module fake_ibex_1772_n_3203 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_688, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_673, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_679, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_672, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3203);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_688;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_673;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_672;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3203;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_850;
wire n_3175;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2333;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2646;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_3117;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3091;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3055;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_907;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2303;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1683;
wire n_1185;
wire n_1122;
wire n_2765;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_1349;
wire n_961;
wire n_1331;
wire n_1223;
wire n_991;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_2862;
wire n_3100;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_768;
wire n_839;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_2818;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_975;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3011;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_786;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3109;
wire n_1961;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3104;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3114;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_866;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_417),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_421),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_594),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_336),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_527),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_222),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_504),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_640),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_272),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_615),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_607),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_199),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_153),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_394),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_80),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_301),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_76),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_599),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_116),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_674),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_667),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_327),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_267),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_348),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_676),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_473),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_31),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_413),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_533),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_192),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_417),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_594),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_690),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_689),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_371),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_401),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_211),
.Y(n_730)
);

CKINVDCx16_ASAP7_75t_R g731 ( 
.A(n_1),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_485),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_502),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_23),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_658),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_181),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_223),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_11),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_393),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_27),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_678),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_626),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_10),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_582),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_62),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_145),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_141),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_305),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_664),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_494),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_683),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_158),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_244),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_370),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_368),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_119),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_639),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_39),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_595),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_215),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_109),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_439),
.Y(n_763)
);

BUFx5_ASAP7_75t_L g764 ( 
.A(n_308),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_226),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_206),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_311),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_397),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_322),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_211),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_18),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_215),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_32),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_408),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_688),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_303),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_474),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_321),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_184),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_388),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_588),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_282),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_574),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_145),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_628),
.Y(n_785)
);

CKINVDCx14_ASAP7_75t_R g786 ( 
.A(n_565),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_80),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_261),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_312),
.Y(n_789)
);

CKINVDCx16_ASAP7_75t_R g790 ( 
.A(n_666),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_4),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_61),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_243),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_216),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_393),
.Y(n_795)
);

BUFx10_ASAP7_75t_L g796 ( 
.A(n_2),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_83),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_299),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_60),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_86),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_291),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_99),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_562),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_252),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_662),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_465),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_488),
.Y(n_807)
);

CKINVDCx11_ASAP7_75t_R g808 ( 
.A(n_112),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_277),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_346),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_3),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_527),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_572),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_563),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_561),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_97),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_474),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_230),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_237),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_521),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_362),
.Y(n_821)
);

CKINVDCx14_ASAP7_75t_R g822 ( 
.A(n_435),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_562),
.Y(n_823)
);

CKINVDCx16_ASAP7_75t_R g824 ( 
.A(n_86),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_671),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_559),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_51),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_672),
.Y(n_828)
);

BUFx10_ASAP7_75t_L g829 ( 
.A(n_123),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_444),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_670),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_288),
.Y(n_832)
);

BUFx5_ASAP7_75t_L g833 ( 
.A(n_112),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_536),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_389),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_387),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_608),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_365),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_521),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_236),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_191),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_685),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_612),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_262),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_271),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_395),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_339),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_1),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_133),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_640),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_661),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_41),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_116),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_436),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_66),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_626),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_367),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_73),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_665),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_0),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_195),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_308),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_569),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_673),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_682),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_87),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_578),
.Y(n_867)
);

BUFx8_ASAP7_75t_SL g868 ( 
.A(n_318),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_140),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_652),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_513),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_307),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_624),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_399),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_184),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_111),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_201),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_61),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_642),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_234),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_602),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_359),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_341),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_637),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_299),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_412),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_687),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_163),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_96),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_448),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_435),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_194),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_512),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_114),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_641),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_24),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_231),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_537),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_373),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_510),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_174),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_349),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_488),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_187),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_119),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_681),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_131),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_494),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_138),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_599),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_13),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_394),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_21),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_608),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_491),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_605),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_437),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_364),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_246),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_357),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_377),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_574),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_575),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_241),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_52),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_283),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_421),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_545),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_114),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_43),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_433),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_70),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_456),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_39),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_316),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_162),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_445),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_543),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_52),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_258),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_506),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_359),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_332),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_233),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_216),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_376),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_344),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_161),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_535),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_503),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_663),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_679),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_391),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_101),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_339),
.Y(n_955)
);

BUFx10_ASAP7_75t_L g956 ( 
.A(n_544),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_126),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_466),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_547),
.Y(n_959)
);

BUFx2_ASAP7_75t_SL g960 ( 
.A(n_380),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_81),
.Y(n_961)
);

BUFx5_ASAP7_75t_L g962 ( 
.A(n_188),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_675),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_218),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_115),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_546),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_467),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_382),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_76),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_306),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_331),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_311),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_323),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_524),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_298),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_100),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_686),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_519),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_570),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_684),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_95),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_48),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_59),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_141),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_94),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_496),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_229),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_368),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_73),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_317),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_202),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_130),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_405),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_159),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_22),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_19),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_399),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_48),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_62),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_370),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_569),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_181),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_571),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_244),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_508),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_534),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_284),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_11),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_96),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_50),
.Y(n_1010)
);

CKINVDCx16_ASAP7_75t_R g1011 ( 
.A(n_526),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_291),
.Y(n_1012)
);

BUFx10_ASAP7_75t_L g1013 ( 
.A(n_360),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_254),
.Y(n_1014)
);

BUFx5_ASAP7_75t_L g1015 ( 
.A(n_356),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_257),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_531),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_170),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_397),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_155),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_143),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_677),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_590),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_369),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_40),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_50),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_103),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_654),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_63),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_508),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_613),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_526),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_578),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_157),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_532),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_25),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_495),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_275),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_8),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_134),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_314),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_78),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_637),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_522),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_47),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_614),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_229),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_269),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_414),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_286),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_161),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_615),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_497),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_122),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_193),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_501),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_152),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_419),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_3),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_0),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_217),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_15),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_790),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_698),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_868),
.Y(n_1065)
);

INVxp67_ASAP7_75t_L g1066 ( 
.A(n_694),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_698),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_711),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_711),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_808),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_733),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_733),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_865),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_831),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_786),
.Y(n_1075)
);

INVxp33_ASAP7_75t_SL g1076 ( 
.A(n_874),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_808),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_753),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_709),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_731),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_753),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_777),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_764),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_822),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_792),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_709),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_721),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_827),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_792),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_848),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_848),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_721),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_824),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_922),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_722),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_720),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_718),
.B(n_4),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_720),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_844),
.B(n_5),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_862),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_846),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_774),
.B(n_6),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_751),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_722),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_935),
.B(n_971),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_723),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_764),
.Y(n_1107)
);

INVxp33_ASAP7_75t_SL g1108 ( 
.A(n_723),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_751),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_984),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1005),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_788),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_794),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_707),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_724),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_794),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_718),
.B(n_6),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_7),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_821),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_726),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_821),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_872),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_953),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_882),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_882),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_724),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_936),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_936),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_986),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_725),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_986),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_725),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_995),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_732),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_732),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_998),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_749),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_865),
.Y(n_1138)
);

INVx4_ASAP7_75t_R g1139 ( 
.A(n_727),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1041),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_761),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_761),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_823),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_834),
.B(n_7),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_823),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_952),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_796),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1041),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_1011),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_691),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_764),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_835),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1042),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1042),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_841),
.B(n_8),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_796),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1043),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_860),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_860),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_903),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_903),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_691),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_712),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_918),
.B(n_9),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1043),
.Y(n_1165)
);

INVxp33_ASAP7_75t_SL g1166 ( 
.A(n_1044),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_693),
.B(n_10),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_919),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1064),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1146),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1079),
.B(n_750),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1067),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1087),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1092),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1073),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1140),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1114),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1068),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1073),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1069),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1083),
.B(n_742),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1150),
.A2(n_739),
.B1(n_759),
.B2(n_712),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1138),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1146),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1114),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1150),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1071),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1130),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1072),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1114),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1081),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1085),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1095),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1107),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1114),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1089),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1090),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1091),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1151),
.A2(n_775),
.B(n_752),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1094),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1137),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1086),
.B(n_1096),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1098),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1100),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1141),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1103),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1109),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1104),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1108),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1120),
.B(n_805),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1112),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1113),
.B(n_825),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1116),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1119),
.B(n_887),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1121),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1122),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1124),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1125),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1127),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1142),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1128),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1129),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1131),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1133),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1110),
.B(n_829),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1070),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1152),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1143),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1076),
.A2(n_759),
.B1(n_771),
.B2(n_739),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1167),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1161),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1145),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1106),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1147),
.B(n_828),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1158),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1166),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1159),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1160),
.Y(n_1239)
);

NAND2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1118),
.B(n_707),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1115),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1066),
.B(n_829),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1168),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1117),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1117),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1156),
.Y(n_1246)
);

NAND2xp33_ASAP7_75t_SL g1247 ( 
.A(n_1063),
.B(n_1075),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1164),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1102),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1105),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1144),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1155),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1126),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1132),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1111),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1134),
.A2(n_1046),
.B1(n_1049),
.B2(n_1045),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1135),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1139),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1093),
.B(n_838),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1065),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1148),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1153),
.B(n_919),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1154),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1123),
.A2(n_793),
.B1(n_795),
.B2(n_771),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1157),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1165),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1149),
.B(n_1084),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1074),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1080),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1080),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1082),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1070),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1077),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1077),
.Y(n_1274)
);

XOR2xp5_ASAP7_75t_L g1275 ( 
.A(n_1082),
.B(n_1062),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1101),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1136),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1162),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1163),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1064),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1073),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1088),
.B(n_838),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1073),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1130),
.Y(n_1285)
);

AND2x2_ASAP7_75t_SL g1286 ( 
.A(n_1097),
.B(n_931),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1064),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1114),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1088),
.B(n_884),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1073),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1120),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1064),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1146),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1064),
.Y(n_1294)
);

INVx5_ASAP7_75t_L g1295 ( 
.A(n_1114),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1130),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1099),
.B(n_707),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1099),
.A2(n_1049),
.B1(n_1061),
.B2(n_1060),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1130),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1087),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1130),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1064),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1073),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1064),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1146),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1064),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1064),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1083),
.B(n_963),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1064),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1065),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1146),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1083),
.A2(n_932),
.B(n_931),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1079),
.B(n_764),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1064),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1064),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1064),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1146),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1064),
.B(n_955),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1130),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1064),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1064),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1079),
.B(n_764),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1064),
.B(n_963),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1099),
.A2(n_1055),
.B1(n_1058),
.B2(n_1053),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1250),
.A2(n_1059),
.B1(n_695),
.B2(n_696),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1291),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1189),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1291),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1201),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1313),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1183),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1176),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1176),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1200),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1291),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1325),
.B(n_697),
.C(n_692),
.Y(n_1338)
);

BUFx10_ASAP7_75t_L g1339 ( 
.A(n_1205),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1205),
.B(n_956),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1170),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1170),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1210),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1184),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1244),
.B(n_713),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1202),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1261),
.B(n_701),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1184),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1266),
.B(n_705),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1230),
.B(n_710),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1245),
.B(n_714),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1230),
.B(n_728),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1293),
.B(n_842),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1298),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1298),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1188),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1237),
.B(n_1231),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1237),
.B(n_996),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1306),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1246),
.B(n_906),
.Y(n_1360)
);

CKINVDCx8_ASAP7_75t_R g1361 ( 
.A(n_1311),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1173),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1206),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1312),
.B(n_1318),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1318),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1228),
.B(n_859),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1169),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1172),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1188),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1264),
.B(n_740),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1232),
.B(n_864),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_L g1372 ( 
.A(n_1254),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1258),
.B(n_706),
.Y(n_1373)
);

XNOR2xp5_ASAP7_75t_L g1374 ( 
.A(n_1275),
.B(n_793),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1174),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1264),
.B(n_765),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1254),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1285),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1206),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1194),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1286),
.B(n_951),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1325),
.B(n_700),
.C(n_699),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1286),
.B(n_977),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1178),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1255),
.B(n_980),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1221),
.Y(n_1386)
);

AND2x6_ASAP7_75t_L g1387 ( 
.A(n_1257),
.B(n_955),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1180),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1260),
.B(n_960),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1221),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1285),
.B(n_803),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1187),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1209),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1277),
.B(n_795),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1241),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1203),
.B(n_1171),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1236),
.Y(n_1397)
);

INVx2_ASAP7_75t_SL g1398 ( 
.A(n_1302),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_SL g1399 ( 
.A(n_1257),
.B(n_1057),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1190),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1211),
.B(n_1022),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1192),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1193),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1301),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1265),
.B(n_1262),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1302),
.B(n_811),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1320),
.B(n_1013),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1257),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1186),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1262),
.B(n_708),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_L g1411 ( 
.A(n_1263),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1296),
.A2(n_1039),
.B1(n_1040),
.B2(n_1037),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_R g1413 ( 
.A(n_1311),
.B(n_1038),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1296),
.A2(n_703),
.B1(n_704),
.B2(n_702),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1238),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1300),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1320),
.B(n_1013),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1197),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1175),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1234),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1179),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1198),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1249),
.B(n_719),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1242),
.B(n_830),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1281),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1235),
.B(n_830),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1199),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1256),
.B(n_853),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1229),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1282),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1324),
.B(n_830),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1263),
.Y(n_1432)
);

INVx4_ASAP7_75t_SL g1433 ( 
.A(n_1263),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1284),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1253),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1287),
.A2(n_730),
.B1(n_734),
.B2(n_729),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1227),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1251),
.B(n_735),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1290),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1292),
.Y(n_1440)
);

AND2x6_ASAP7_75t_L g1441 ( 
.A(n_1259),
.B(n_979),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1294),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_SL g1443 ( 
.A(n_1253),
.B(n_798),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1256),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1299),
.A2(n_716),
.B1(n_717),
.B2(n_715),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1303),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_SL g1447 ( 
.A(n_1272),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1226),
.B(n_836),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1319),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1283),
.B(n_836),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1299),
.A2(n_745),
.B1(n_747),
.B2(n_738),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1305),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1289),
.B(n_836),
.Y(n_1453)
);

AND2x6_ASAP7_75t_L g1454 ( 
.A(n_1267),
.B(n_979),
.Y(n_1454)
);

AO22x2_ASAP7_75t_L g1455 ( 
.A1(n_1182),
.A2(n_826),
.B1(n_845),
.B2(n_798),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1227),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1314),
.A2(n_737),
.B(n_736),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1304),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1307),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1308),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1270),
.B(n_911),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1280),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1310),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1240),
.B(n_855),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1297),
.B(n_855),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1315),
.B(n_1316),
.Y(n_1466)
);

NOR2x1p5_ASAP7_75t_L g1467 ( 
.A(n_1269),
.B(n_754),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1252),
.B(n_1248),
.Y(n_1468)
);

INVx8_ASAP7_75t_L g1469 ( 
.A(n_1269),
.Y(n_1469)
);

CKINVDCx8_ASAP7_75t_R g1470 ( 
.A(n_1186),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1317),
.B(n_755),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1233),
.Y(n_1472)
);

INVx4_ASAP7_75t_SL g1473 ( 
.A(n_1268),
.Y(n_1473)
);

AND2x6_ASAP7_75t_L g1474 ( 
.A(n_1323),
.B(n_1002),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1309),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1321),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1322),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1271),
.A2(n_845),
.B1(n_849),
.B2(n_826),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1239),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1243),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1297),
.B(n_1309),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1214),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1204),
.B(n_757),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1247),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1222),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1207),
.B(n_758),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1223),
.Y(n_1487)
);

AND2x6_ASAP7_75t_L g1488 ( 
.A(n_1208),
.B(n_1002),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1225),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1212),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1216),
.B(n_760),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1217),
.A2(n_1036),
.B1(n_1035),
.B2(n_762),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1218),
.Y(n_1493)
);

BUFx10_ASAP7_75t_L g1494 ( 
.A(n_1276),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1219),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1277),
.B(n_1213),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1220),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1247),
.Y(n_1498)
);

AND2x6_ASAP7_75t_L g1499 ( 
.A(n_1224),
.B(n_1008),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1273),
.Y(n_1500)
);

OR2x6_ASAP7_75t_L g1501 ( 
.A(n_1274),
.B(n_849),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1215),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1278),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1181),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1181),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1195),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1279),
.B(n_741),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1295),
.B(n_743),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1295),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1177),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1185),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1185),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1191),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1191),
.B(n_744),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1191),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1196),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1196),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1288),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1288),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1356),
.A2(n_975),
.B1(n_958),
.B2(n_767),
.C(n_769),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1367),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1368),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1396),
.B(n_763),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1334),
.B(n_746),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1502),
.B(n_766),
.Y(n_1525)
);

BUFx8_ASAP7_75t_L g1526 ( 
.A(n_1447),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1335),
.B(n_748),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1416),
.A2(n_1398),
.B1(n_1378),
.B2(n_1369),
.Y(n_1528)
);

AO22x2_ASAP7_75t_L g1529 ( 
.A1(n_1350),
.A2(n_876),
.B1(n_886),
.B2(n_856),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1339),
.B(n_770),
.Y(n_1530)
);

AO22x2_ASAP7_75t_L g1531 ( 
.A1(n_1352),
.A2(n_886),
.B1(n_899),
.B2(n_876),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1409),
.A2(n_902),
.B1(n_907),
.B2(n_899),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1339),
.B(n_772),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1429),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1429),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1496),
.A2(n_780),
.B1(n_781),
.B2(n_779),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1384),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1473),
.B(n_1328),
.Y(n_1538)
);

AO22x2_ASAP7_75t_L g1539 ( 
.A1(n_1370),
.A2(n_1376),
.B1(n_1420),
.B2(n_1404),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1388),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1437),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1392),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1413),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1400),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1402),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1403),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1343),
.Y(n_1547)
);

AO22x2_ASAP7_75t_L g1548 ( 
.A1(n_1428),
.A2(n_907),
.B1(n_924),
.B2(n_902),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1418),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1375),
.B(n_924),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1422),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1380),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1425),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1473),
.B(n_756),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1393),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1395),
.B(n_940),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1444),
.A2(n_791),
.B1(n_797),
.B2(n_789),
.C(n_787),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1330),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1357),
.B(n_940),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1440),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1391),
.B(n_799),
.Y(n_1561)
);

NAND2x1p5_ASAP7_75t_L g1562 ( 
.A(n_1427),
.B(n_768),
.Y(n_1562)
);

AO22x2_ASAP7_75t_L g1563 ( 
.A1(n_1455),
.A2(n_970),
.B1(n_972),
.B2(n_943),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1442),
.Y(n_1564)
);

AO22x2_ASAP7_75t_L g1565 ( 
.A1(n_1455),
.A2(n_970),
.B1(n_972),
.B2(n_943),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1446),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1452),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1459),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1460),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1463),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1476),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_SL g1572 ( 
.A(n_1389),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1427),
.B(n_800),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1435),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1443),
.Y(n_1575)
);

AO22x2_ASAP7_75t_L g1576 ( 
.A1(n_1406),
.A2(n_1018),
.B1(n_1026),
.B2(n_994),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1477),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1479),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1490),
.Y(n_1579)
);

AO22x2_ASAP7_75t_L g1580 ( 
.A1(n_1478),
.A2(n_1362),
.B1(n_1382),
.B2(n_1338),
.Y(n_1580)
);

CKINVDCx16_ASAP7_75t_R g1581 ( 
.A(n_1394),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1493),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1372),
.B(n_773),
.Y(n_1583)
);

AO22x2_ASAP7_75t_L g1584 ( 
.A1(n_1433),
.A2(n_1026),
.B1(n_1027),
.B2(n_1018),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1326),
.B(n_1329),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1374),
.A2(n_1051),
.B1(n_1052),
.B2(n_1027),
.Y(n_1586)
);

BUFx8_ASAP7_75t_L g1587 ( 
.A(n_1447),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1469),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1361),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_L g1590 ( 
.A(n_1488),
.B(n_833),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1469),
.B(n_1008),
.Y(n_1591)
);

NAND2x1p5_ASAP7_75t_L g1592 ( 
.A(n_1372),
.B(n_776),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1467),
.B(n_1052),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_SL g1594 ( 
.A(n_1500),
.B(n_1062),
.C(n_1057),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1326),
.B(n_802),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1466),
.Y(n_1596)
);

NAND2xp33_ASAP7_75t_L g1597 ( 
.A(n_1488),
.B(n_833),
.Y(n_1597)
);

AO22x2_ASAP7_75t_L g1598 ( 
.A1(n_1410),
.A2(n_1451),
.B1(n_1445),
.B2(n_1347),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1495),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1456),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1497),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1472),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1407),
.B(n_806),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1514),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1411),
.B(n_778),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1411),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1480),
.Y(n_1607)
);

AO22x2_ASAP7_75t_L g1608 ( 
.A1(n_1347),
.A2(n_783),
.B1(n_784),
.B2(n_782),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1389),
.B(n_785),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1514),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1485),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1470),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1489),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1417),
.B(n_810),
.Y(n_1614)
);

AO22x2_ASAP7_75t_L g1615 ( 
.A1(n_1349),
.A2(n_804),
.B1(n_807),
.B2(n_801),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1337),
.B(n_809),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1349),
.A2(n_813),
.B1(n_814),
.B2(n_812),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1501),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1340),
.B(n_1358),
.Y(n_1619)
);

AO22x2_ASAP7_75t_L g1620 ( 
.A1(n_1507),
.A2(n_820),
.B1(n_832),
.B2(n_816),
.Y(n_1620)
);

AO22x2_ASAP7_75t_L g1621 ( 
.A1(n_1507),
.A2(n_839),
.B1(n_843),
.B2(n_837),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1494),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1462),
.A2(n_818),
.B1(n_819),
.B2(n_817),
.C(n_815),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1461),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1364),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1331),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1487),
.B(n_1329),
.Y(n_1627)
);

BUFx8_ASAP7_75t_L g1628 ( 
.A(n_1503),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1449),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1449),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1405),
.B(n_854),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1449),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1341),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1342),
.Y(n_1634)
);

BUFx8_ASAP7_75t_L g1635 ( 
.A(n_1454),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1344),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1348),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1381),
.A2(n_873),
.B1(n_875),
.B2(n_871),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1482),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_L g1640 ( 
.A(n_1412),
.B(n_12),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1354),
.Y(n_1641)
);

BUFx8_ASAP7_75t_L g1642 ( 
.A(n_1454),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1359),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1365),
.Y(n_1644)
);

AO22x2_ASAP7_75t_L g1645 ( 
.A1(n_1399),
.A2(n_889),
.B1(n_896),
.B2(n_881),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1408),
.B(n_898),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1432),
.B(n_900),
.Y(n_1647)
);

AO22x2_ASAP7_75t_L g1648 ( 
.A1(n_1336),
.A2(n_904),
.B1(n_905),
.B2(n_901),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1498),
.B(n_1024),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1432),
.B(n_912),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1383),
.A2(n_916),
.B1(n_926),
.B2(n_913),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1494),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1484),
.Y(n_1653)
);

BUFx8_ASAP7_75t_L g1654 ( 
.A(n_1454),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1474),
.A2(n_927),
.B1(n_930),
.B2(n_929),
.Y(n_1655)
);

AND2x6_ASAP7_75t_L g1656 ( 
.A(n_1508),
.B(n_1024),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1414),
.B(n_840),
.Y(n_1657)
);

AO22x2_ASAP7_75t_L g1658 ( 
.A1(n_1336),
.A2(n_938),
.B1(n_941),
.B2(n_937),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1468),
.Y(n_1659)
);

NAND2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1355),
.B(n_944),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1468),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1355),
.B(n_945),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1419),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1499),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1454),
.A2(n_850),
.B1(n_851),
.B2(n_847),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1421),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1327),
.B(n_852),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1430),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1436),
.A2(n_858),
.B1(n_863),
.B2(n_861),
.C(n_857),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1441),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1441),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1434),
.Y(n_1672)
);

AO22x2_ASAP7_75t_L g1673 ( 
.A1(n_1481),
.A2(n_966),
.B1(n_969),
.B2(n_961),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1508),
.B(n_973),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1373),
.B(n_976),
.Y(n_1675)
);

AO22x2_ASAP7_75t_L g1676 ( 
.A1(n_1423),
.A2(n_990),
.B1(n_997),
.B2(n_987),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1439),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1377),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1415),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1492),
.A2(n_867),
.B1(n_870),
.B2(n_869),
.C(n_866),
.Y(n_1680)
);

AO22x2_ASAP7_75t_L g1681 ( 
.A1(n_1423),
.A2(n_1003),
.B1(n_1006),
.B2(n_1001),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1415),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1385),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1415),
.Y(n_1684)
);

AO22x2_ASAP7_75t_L g1685 ( 
.A1(n_1438),
.A2(n_1016),
.B1(n_1032),
.B2(n_1009),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1475),
.A2(n_1047),
.B1(n_1048),
.B2(n_1034),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1387),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1483),
.A2(n_1491),
.B1(n_1486),
.B2(n_1471),
.C(n_1345),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1506),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1448),
.B(n_1050),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1458),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1387),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1360),
.A2(n_877),
.B1(n_879),
.B2(n_878),
.Y(n_1693)
);

AO22x2_ASAP7_75t_L g1694 ( 
.A1(n_1450),
.A2(n_1054),
.B1(n_1056),
.B2(n_1050),
.Y(n_1694)
);

AO22x2_ASAP7_75t_L g1695 ( 
.A1(n_1453),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1351),
.B(n_880),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1426),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1424),
.B(n_883),
.Y(n_1698)
);

AO22x2_ASAP7_75t_L g1699 ( 
.A1(n_1332),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1366),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1371),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1387),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1457),
.A2(n_888),
.B1(n_891),
.B2(n_890),
.C(n_885),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1353),
.B(n_892),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1401),
.B(n_893),
.Y(n_1705)
);

CKINVDCx14_ASAP7_75t_R g1706 ( 
.A(n_1509),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1333),
.B(n_894),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1363),
.B(n_1379),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1709)
);

AO22x2_ASAP7_75t_L g1710 ( 
.A1(n_1464),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1431),
.B(n_895),
.Y(n_1711)
);

AO22x2_ASAP7_75t_L g1712 ( 
.A1(n_1465),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1390),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1397),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1346),
.B(n_897),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_SL g1716 ( 
.A(n_1510),
.Y(n_1716)
);

NAND2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1510),
.B(n_928),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1386),
.A2(n_962),
.B1(n_1015),
.B2(n_833),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1596),
.B(n_1700),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1524),
.B(n_908),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1574),
.B(n_909),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1528),
.B(n_910),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1547),
.B(n_914),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1575),
.B(n_915),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1622),
.B(n_917),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1701),
.B(n_1511),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1664),
.B(n_1513),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1523),
.B(n_920),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1652),
.B(n_921),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1552),
.B(n_923),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1665),
.B(n_1555),
.Y(n_1731)
);

NAND2xp33_ASAP7_75t_SL g1732 ( 
.A(n_1670),
.B(n_928),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1606),
.B(n_925),
.Y(n_1733)
);

NAND2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1692),
.B(n_928),
.Y(n_1734)
);

NAND2xp33_ASAP7_75t_SL g1735 ( 
.A(n_1692),
.B(n_1687),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1619),
.B(n_933),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1702),
.B(n_934),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1606),
.B(n_939),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1521),
.B(n_942),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1550),
.B(n_946),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_SL g1742 ( 
.A(n_1572),
.B(n_947),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1616),
.B(n_948),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1527),
.B(n_949),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1527),
.B(n_950),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1537),
.B(n_1516),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1635),
.B(n_954),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1642),
.B(n_957),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1654),
.B(n_959),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1540),
.B(n_964),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1660),
.B(n_965),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1662),
.B(n_1031),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1671),
.B(n_1033),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1543),
.B(n_967),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_SL g1755 ( 
.A(n_1716),
.B(n_968),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1542),
.B(n_974),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1675),
.B(n_978),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1583),
.B(n_981),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1592),
.B(n_982),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1544),
.B(n_1518),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1545),
.B(n_983),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1589),
.B(n_985),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1605),
.B(n_1581),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1546),
.B(n_1512),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1588),
.B(n_988),
.Y(n_1765)
);

NAND2xp33_ASAP7_75t_SL g1766 ( 
.A(n_1618),
.B(n_989),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1624),
.B(n_1025),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1628),
.B(n_1536),
.Y(n_1768)
);

AND2x2_ASAP7_75t_SL g1769 ( 
.A(n_1590),
.B(n_934),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_SL g1770 ( 
.A(n_1538),
.B(n_991),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1549),
.B(n_992),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1556),
.B(n_993),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1646),
.B(n_999),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1647),
.B(n_1000),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1538),
.B(n_1004),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1650),
.B(n_1007),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1561),
.B(n_1010),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1674),
.B(n_1012),
.Y(n_1778)
);

NAND2xp33_ASAP7_75t_SL g1779 ( 
.A(n_1627),
.B(n_1014),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1603),
.B(n_1017),
.Y(n_1780)
);

NAND2xp33_ASAP7_75t_SL g1781 ( 
.A(n_1525),
.B(n_1019),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1614),
.B(n_1028),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1559),
.B(n_1029),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1539),
.B(n_1021),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_SL g1785 ( 
.A(n_1532),
.B(n_1023),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1683),
.B(n_1030),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1551),
.B(n_962),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1788)
);

NAND2xp33_ASAP7_75t_SL g1789 ( 
.A(n_1530),
.B(n_1517),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1533),
.B(n_1519),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1560),
.B(n_26),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1564),
.B(n_26),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1566),
.B(n_28),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1567),
.B(n_28),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_SL g1795 ( 
.A(n_1578),
.B(n_29),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1625),
.B(n_29),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1562),
.B(n_30),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1678),
.B(n_32),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1640),
.B(n_1593),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1554),
.B(n_33),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1631),
.B(n_34),
.Y(n_1801)
);

NAND2xp33_ASAP7_75t_SL g1802 ( 
.A(n_1653),
.B(n_35),
.Y(n_1802)
);

NAND2xp33_ASAP7_75t_SL g1803 ( 
.A(n_1599),
.B(n_35),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1631),
.B(n_36),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1655),
.B(n_36),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1693),
.B(n_37),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1609),
.B(n_37),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1657),
.B(n_38),
.Y(n_1808)
);

NAND2xp33_ASAP7_75t_SL g1809 ( 
.A(n_1601),
.B(n_40),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1568),
.B(n_1569),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1570),
.B(n_42),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1602),
.B(n_42),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1571),
.B(n_44),
.Y(n_1813)
);

NAND2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1607),
.B(n_44),
.Y(n_1814)
);

NAND2xp33_ASAP7_75t_SL g1815 ( 
.A(n_1577),
.B(n_45),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_SL g1816 ( 
.A(n_1579),
.B(n_46),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1667),
.B(n_49),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1698),
.B(n_53),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1612),
.B(n_54),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1582),
.B(n_55),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1580),
.B(n_55),
.Y(n_1821)
);

NAND2xp33_ASAP7_75t_SL g1822 ( 
.A(n_1611),
.B(n_56),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1613),
.B(n_56),
.Y(n_1823)
);

AND2x2_ASAP7_75t_SL g1824 ( 
.A(n_1597),
.B(n_57),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1691),
.B(n_58),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1558),
.B(n_63),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1608),
.B(n_1615),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1715),
.B(n_64),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1586),
.B(n_1594),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1615),
.B(n_1617),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1711),
.B(n_65),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1604),
.B(n_67),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1617),
.B(n_68),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1620),
.B(n_69),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1638),
.B(n_70),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1659),
.B(n_71),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_SL g1837 ( 
.A(n_1661),
.B(n_71),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1610),
.B(n_72),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1651),
.B(n_74),
.Y(n_1839)
);

NAND2xp33_ASAP7_75t_SL g1840 ( 
.A(n_1534),
.B(n_75),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1705),
.B(n_75),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1621),
.B(n_77),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1535),
.B(n_79),
.Y(n_1843)
);

NAND2xp33_ASAP7_75t_SL g1844 ( 
.A(n_1663),
.B(n_82),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1666),
.B(n_84),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1668),
.B(n_85),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1686),
.B(n_87),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_SL g1848 ( 
.A(n_1672),
.B(n_88),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1686),
.B(n_88),
.Y(n_1849)
);

NAND2xp33_ASAP7_75t_SL g1850 ( 
.A(n_1677),
.B(n_89),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1689),
.B(n_90),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1629),
.B(n_90),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_SL g1853 ( 
.A(n_1696),
.B(n_91),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1630),
.B(n_91),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1632),
.B(n_92),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1717),
.B(n_93),
.Y(n_1856)
);

NAND2xp33_ASAP7_75t_SL g1857 ( 
.A(n_1595),
.B(n_93),
.Y(n_1857)
);

NAND2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1704),
.B(n_1541),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1600),
.B(n_95),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1688),
.B(n_1557),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1714),
.B(n_98),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1598),
.B(n_99),
.Y(n_1862)
);

NAND2xp33_ASAP7_75t_SL g1863 ( 
.A(n_1656),
.B(n_100),
.Y(n_1863)
);

NAND2xp33_ASAP7_75t_SL g1864 ( 
.A(n_1656),
.B(n_101),
.Y(n_1864)
);

NAND2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1585),
.B(n_102),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1648),
.B(n_104),
.Y(n_1866)
);

NAND2xp33_ASAP7_75t_SL g1867 ( 
.A(n_1639),
.B(n_105),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1713),
.B(n_105),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1626),
.B(n_106),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1526),
.B(n_107),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1648),
.B(n_108),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1658),
.B(n_108),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1587),
.B(n_110),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1633),
.B(n_1634),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1636),
.B(n_110),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1637),
.B(n_113),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1529),
.B(n_113),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1658),
.B(n_115),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1641),
.B(n_117),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1643),
.B(n_118),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_SL g1881 ( 
.A(n_1709),
.B(n_120),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1644),
.B(n_121),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1676),
.B(n_122),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1573),
.B(n_124),
.Y(n_1884)
);

NAND2xp33_ASAP7_75t_SL g1885 ( 
.A(n_1679),
.B(n_124),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1591),
.B(n_125),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1676),
.B(n_127),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1681),
.B(n_1685),
.Y(n_1888)
);

NAND2xp33_ASAP7_75t_SL g1889 ( 
.A(n_1682),
.B(n_127),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1681),
.B(n_128),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_SL g1891 ( 
.A(n_1684),
.B(n_129),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1697),
.B(n_130),
.Y(n_1892)
);

NAND2xp33_ASAP7_75t_SL g1893 ( 
.A(n_1707),
.B(n_132),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1708),
.B(n_133),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1718),
.B(n_135),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1529),
.B(n_136),
.Y(n_1896)
);

NAND2xp33_ASAP7_75t_SL g1897 ( 
.A(n_1584),
.B(n_137),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1706),
.B(n_139),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1680),
.B(n_140),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1591),
.B(n_142),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1649),
.B(n_143),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1531),
.B(n_144),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1520),
.B(n_146),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1649),
.B(n_147),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1690),
.B(n_148),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1531),
.B(n_148),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1623),
.B(n_149),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1673),
.B(n_150),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_SL g1909 ( 
.A(n_1645),
.B(n_1699),
.Y(n_1909)
);

NAND2xp33_ASAP7_75t_SL g1910 ( 
.A(n_1645),
.B(n_151),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1673),
.B(n_152),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1690),
.B(n_153),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1694),
.B(n_154),
.Y(n_1913)
);

NAND2xp33_ASAP7_75t_SL g1914 ( 
.A(n_1699),
.B(n_155),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1576),
.B(n_1703),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1695),
.B(n_156),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1576),
.B(n_157),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1669),
.B(n_159),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1548),
.B(n_160),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1548),
.B(n_160),
.Y(n_1920)
);

NAND2xp33_ASAP7_75t_SL g1921 ( 
.A(n_1710),
.B(n_1712),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1710),
.B(n_164),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1712),
.B(n_165),
.Y(n_1923)
);

NAND2xp33_ASAP7_75t_SL g1924 ( 
.A(n_1563),
.B(n_165),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1563),
.B(n_166),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1565),
.B(n_166),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1565),
.B(n_167),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1524),
.B(n_167),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1596),
.B(n_168),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1524),
.B(n_168),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1596),
.B(n_169),
.Y(n_1931)
);

NAND2xp33_ASAP7_75t_SL g1932 ( 
.A(n_1664),
.B(n_171),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1664),
.B(n_171),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1596),
.B(n_172),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1524),
.B(n_173),
.Y(n_1935)
);

NAND2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1664),
.B(n_174),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1524),
.B(n_175),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_SL g1938 ( 
.A(n_1524),
.B(n_176),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1596),
.B(n_177),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1524),
.B(n_177),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1596),
.B(n_178),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1524),
.B(n_178),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1524),
.B(n_179),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1524),
.B(n_180),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1524),
.B(n_182),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1524),
.B(n_182),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1524),
.B(n_183),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1524),
.B(n_183),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1524),
.B(n_185),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1524),
.B(n_186),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1524),
.B(n_187),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1524),
.B(n_188),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1574),
.B(n_189),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_SL g1954 ( 
.A(n_1664),
.B(n_189),
.Y(n_1954)
);

XNOR2x2_ASAP7_75t_L g1955 ( 
.A(n_1576),
.B(n_190),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1524),
.B(n_191),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1524),
.B(n_192),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1596),
.B(n_193),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1596),
.B(n_196),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1524),
.B(n_197),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1596),
.B(n_198),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_SL g1962 ( 
.A(n_1664),
.B(n_200),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1524),
.B(n_200),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1524),
.B(n_201),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1524),
.B(n_202),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1524),
.B(n_203),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1596),
.B(n_204),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1574),
.B(n_205),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1524),
.B(n_206),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1524),
.B(n_207),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1664),
.B(n_208),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1524),
.B(n_208),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1524),
.B(n_209),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1574),
.B(n_210),
.Y(n_1974)
);

NAND2xp33_ASAP7_75t_SL g1975 ( 
.A(n_1664),
.B(n_212),
.Y(n_1975)
);

NAND2xp33_ASAP7_75t_SL g1976 ( 
.A(n_1664),
.B(n_213),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1596),
.B(n_214),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1574),
.B(n_214),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1524),
.B(n_217),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1524),
.B(n_219),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1524),
.B(n_219),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1524),
.B(n_220),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_SL g1983 ( 
.A(n_1524),
.B(n_221),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1574),
.B(n_221),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1664),
.B(n_222),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1664),
.B(n_223),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1524),
.B(n_224),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1524),
.B(n_224),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1664),
.B(n_225),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1596),
.B(n_226),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1524),
.B(n_227),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1596),
.B(n_227),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1524),
.B(n_228),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1524),
.B(n_228),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1524),
.B(n_230),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1596),
.B(n_231),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1664),
.B(n_232),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1524),
.B(n_232),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1596),
.B(n_235),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1524),
.B(n_238),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1524),
.B(n_238),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1524),
.B(n_239),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1524),
.B(n_239),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1596),
.B(n_240),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1524),
.B(n_240),
.Y(n_2005)
);

NAND2xp33_ASAP7_75t_SL g2006 ( 
.A(n_1664),
.B(n_242),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1574),
.B(n_242),
.Y(n_2007)
);

NAND2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1664),
.B(n_245),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1524),
.B(n_246),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1524),
.B(n_247),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1524),
.B(n_247),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1524),
.B(n_248),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1596),
.B(n_249),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1524),
.B(n_249),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1574),
.B(n_250),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1524),
.B(n_250),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1664),
.B(n_251),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1664),
.B(n_251),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1596),
.B(n_252),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1719),
.Y(n_2020)
);

AO31x2_ASAP7_75t_L g2021 ( 
.A1(n_1821),
.A2(n_255),
.A3(n_253),
.B(n_254),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1931),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1719),
.B(n_253),
.Y(n_2023)
);

BUFx4f_ASAP7_75t_L g2024 ( 
.A(n_1886),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1719),
.B(n_255),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1860),
.B(n_256),
.Y(n_2026)
);

OAI22x1_ASAP7_75t_L g2027 ( 
.A1(n_1925),
.A2(n_1886),
.B1(n_1927),
.B2(n_1926),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1793),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1834),
.B(n_1925),
.Y(n_2029)
);

NAND2x1p5_ASAP7_75t_L g2030 ( 
.A(n_1886),
.B(n_259),
.Y(n_2030)
);

NAND3x1_ASAP7_75t_L g2031 ( 
.A(n_1877),
.B(n_259),
.C(n_260),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1925),
.B(n_260),
.Y(n_2032)
);

O2A1O1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1915),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_SL g2034 ( 
.A1(n_1931),
.A2(n_669),
.B(n_668),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_SL g2035 ( 
.A1(n_1827),
.A2(n_263),
.B(n_264),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1726),
.B(n_264),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1918),
.A2(n_265),
.B(n_266),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1810),
.B(n_266),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1909),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2039)
);

NOR2xp67_ASAP7_75t_L g2040 ( 
.A(n_1731),
.B(n_268),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1931),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1830),
.B(n_273),
.Y(n_2042)
);

AO32x2_ASAP7_75t_L g2043 ( 
.A1(n_1921),
.A2(n_276),
.A3(n_273),
.B1(n_274),
.B2(n_277),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1799),
.B(n_274),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1785),
.B(n_278),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1793),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1888),
.B(n_278),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1958),
.Y(n_2048)
);

NOR2xp67_ASAP7_75t_L g2049 ( 
.A(n_1829),
.B(n_279),
.Y(n_2049)
);

NAND3xp33_ASAP7_75t_L g2050 ( 
.A(n_1914),
.B(n_279),
.C(n_280),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1726),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1770),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1726),
.B(n_281),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1787),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1772),
.B(n_282),
.Y(n_2055)
);

NOR2x1_ASAP7_75t_SL g2056 ( 
.A(n_1913),
.B(n_680),
.Y(n_2056)
);

INVx4_ASAP7_75t_L g2057 ( 
.A(n_1901),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1741),
.B(n_1744),
.Y(n_2058)
);

INVxp67_ASAP7_75t_L g2059 ( 
.A(n_1901),
.Y(n_2059)
);

NOR4xp25_ASAP7_75t_L g2060 ( 
.A(n_1917),
.B(n_287),
.C(n_285),
.D(n_286),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1813),
.Y(n_2061)
);

NOR2xp67_ASAP7_75t_L g2062 ( 
.A(n_1763),
.B(n_285),
.Y(n_2062)
);

OAI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1929),
.A2(n_287),
.B(n_288),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_2019),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_SL g2065 ( 
.A1(n_1958),
.A2(n_289),
.B(n_290),
.Y(n_2065)
);

O2A1O1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_1919),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1899),
.B(n_294),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1745),
.B(n_295),
.Y(n_2068)
);

BUFx8_ASAP7_75t_L g2069 ( 
.A(n_1901),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1904),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1959),
.A2(n_1967),
.B1(n_1992),
.B2(n_1990),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1896),
.B(n_296),
.Y(n_2072)
);

OAI21x1_ASAP7_75t_SL g2073 ( 
.A1(n_1847),
.A2(n_1849),
.B(n_1866),
.Y(n_2073)
);

O2A1O1Ixp5_ASAP7_75t_L g2074 ( 
.A1(n_1734),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_SL g2075 ( 
.A1(n_1959),
.A2(n_297),
.B(n_300),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1959),
.B(n_300),
.Y(n_2076)
);

BUFx12f_ASAP7_75t_L g2077 ( 
.A(n_1904),
.Y(n_2077)
);

CKINVDCx11_ASAP7_75t_R g2078 ( 
.A(n_1904),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1934),
.A2(n_302),
.B(n_304),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1721),
.B(n_309),
.Y(n_2080)
);

INVxp67_ASAP7_75t_SL g2081 ( 
.A(n_1967),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1967),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_1905),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1808),
.B(n_310),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1869),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1817),
.B(n_313),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1990),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_1775),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1990),
.A2(n_318),
.B1(n_315),
.B2(n_317),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1905),
.Y(n_2090)
);

NAND2x1p5_ASAP7_75t_L g2091 ( 
.A(n_1905),
.B(n_319),
.Y(n_2091)
);

AO31x2_ASAP7_75t_L g2092 ( 
.A1(n_1862),
.A2(n_324),
.A3(n_320),
.B(n_322),
.Y(n_2092)
);

OAI21xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1824),
.A2(n_325),
.B(n_326),
.Y(n_2093)
);

CKINVDCx11_ASAP7_75t_R g2094 ( 
.A(n_1912),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_SL g2095 ( 
.A1(n_1871),
.A2(n_325),
.B(n_326),
.Y(n_2095)
);

CKINVDCx20_ASAP7_75t_R g2096 ( 
.A(n_1742),
.Y(n_2096)
);

NOR2x1_ASAP7_75t_L g2097 ( 
.A(n_1768),
.B(n_328),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1902),
.B(n_329),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1874),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2019),
.Y(n_2100)
);

OA22x2_ASAP7_75t_L g2101 ( 
.A1(n_1920),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2101)
);

AO31x2_ASAP7_75t_L g2102 ( 
.A1(n_1916),
.A2(n_334),
.A3(n_330),
.B(n_333),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_2019),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1736),
.B(n_333),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_SL g2105 ( 
.A1(n_1872),
.A2(n_334),
.B(n_335),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1992),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1906),
.B(n_335),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1939),
.B(n_337),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1941),
.B(n_338),
.Y(n_2109)
);

OAI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1961),
.A2(n_340),
.B(n_341),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1992),
.A2(n_343),
.B1(n_340),
.B2(n_342),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1936),
.A2(n_342),
.B(n_343),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1977),
.B(n_344),
.Y(n_2113)
);

NAND2x1_ASAP7_75t_L g2114 ( 
.A(n_2004),
.B(n_345),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1912),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_1953),
.B(n_345),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_2004),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2004),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1762),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1908),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_SL g2121 ( 
.A1(n_1936),
.A2(n_347),
.B(n_349),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1968),
.B(n_350),
.Y(n_2122)
);

OAI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1996),
.A2(n_351),
.B(n_352),
.Y(n_2123)
);

OAI21xp33_ASAP7_75t_L g2124 ( 
.A1(n_1922),
.A2(n_352),
.B(n_353),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_SL g2125 ( 
.A1(n_1912),
.A2(n_353),
.B(n_354),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1999),
.A2(n_354),
.B(n_355),
.Y(n_2126)
);

A2O1A1Ixp33_ASAP7_75t_L g2127 ( 
.A1(n_1822),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1769),
.A2(n_358),
.B(n_360),
.Y(n_2128)
);

AO32x2_ASAP7_75t_L g2129 ( 
.A1(n_1955),
.A2(n_362),
.A3(n_358),
.B1(n_361),
.B2(n_363),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_SL g2130 ( 
.A1(n_1878),
.A2(n_361),
.B(n_363),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1911),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1974),
.B(n_365),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1978),
.B(n_366),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1984),
.B(n_369),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1755),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_1740),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2013),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1722),
.B(n_372),
.Y(n_2138)
);

AO32x2_ASAP7_75t_L g2139 ( 
.A1(n_1923),
.A2(n_376),
.A3(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_2139)
);

AOI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_1907),
.A2(n_375),
.B(n_378),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1740),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1728),
.B(n_379),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1835),
.B(n_381),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1740),
.Y(n_2144)
);

AOI21xp33_ASAP7_75t_L g2145 ( 
.A1(n_1784),
.A2(n_383),
.B(n_384),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_1720),
.B(n_385),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1824),
.B(n_386),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1739),
.B(n_387),
.Y(n_2148)
);

AO31x2_ASAP7_75t_L g2149 ( 
.A1(n_1791),
.A2(n_392),
.A3(n_390),
.B(n_391),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1746),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1750),
.B(n_392),
.Y(n_2151)
);

AOI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1895),
.A2(n_396),
.B(n_398),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1756),
.B(n_396),
.Y(n_2153)
);

BUFx24_ASAP7_75t_L g2154 ( 
.A(n_1897),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2007),
.B(n_400),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_1924),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1792),
.A2(n_402),
.B(n_403),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_1766),
.Y(n_2158)
);

BUFx10_ASAP7_75t_L g2159 ( 
.A(n_1746),
.Y(n_2159)
);

AOI221x1_ASAP7_75t_L g2160 ( 
.A1(n_1910),
.A2(n_407),
.B1(n_404),
.B2(n_406),
.C(n_409),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1761),
.B(n_407),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1794),
.Y(n_2162)
);

AOI221x1_ASAP7_75t_L g2163 ( 
.A1(n_1823),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.C(n_413),
.Y(n_2163)
);

INVx3_ASAP7_75t_SL g2164 ( 
.A(n_1747),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1811),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1751),
.B(n_415),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1771),
.B(n_416),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1858),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1831),
.B(n_418),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1833),
.Y(n_2170)
);

NAND2x1p5_ASAP7_75t_L g2171 ( 
.A(n_1748),
.B(n_419),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1818),
.B(n_420),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_1881),
.B(n_422),
.C(n_423),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1783),
.B(n_424),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_1752),
.B(n_425),
.Y(n_2175)
);

AO32x2_ASAP7_75t_L g2176 ( 
.A1(n_1795),
.A2(n_425),
.A3(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_1796),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1732),
.B(n_429),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1932),
.A2(n_429),
.B(n_430),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_1933),
.A2(n_430),
.B(n_431),
.Y(n_2180)
);

AO22x2_ASAP7_75t_L g2181 ( 
.A1(n_1842),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_2181)
);

BUFx2_ASAP7_75t_L g2182 ( 
.A(n_1863),
.Y(n_2182)
);

NOR2xp67_ASAP7_75t_SL g2183 ( 
.A(n_1749),
.B(n_436),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_1743),
.B(n_437),
.Y(n_2184)
);

AO22x2_ASAP7_75t_L g2185 ( 
.A1(n_1883),
.A2(n_441),
.B1(n_438),
.B2(n_440),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2015),
.B(n_441),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_1887),
.B(n_442),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1890),
.B(n_442),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1806),
.A2(n_443),
.B(n_445),
.Y(n_2189)
);

AO32x2_ASAP7_75t_L g2190 ( 
.A1(n_1795),
.A2(n_446),
.A3(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1764),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1764),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1746),
.Y(n_2193)
);

AOI221x1_ASAP7_75t_L g2194 ( 
.A1(n_1986),
.A2(n_446),
.B1(n_447),
.B2(n_449),
.C(n_450),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1732),
.B(n_451),
.Y(n_2195)
);

A2O1A1Ixp33_ASAP7_75t_L g2196 ( 
.A1(n_1881),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_1777),
.B(n_1757),
.Y(n_2197)
);

A2O1A1Ixp33_ASAP7_75t_L g2198 ( 
.A1(n_1989),
.A2(n_454),
.B(n_452),
.C(n_453),
.Y(n_2198)
);

AO31x2_ASAP7_75t_L g2199 ( 
.A1(n_1989),
.A2(n_458),
.A3(n_455),
.B(n_457),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_1903),
.A2(n_457),
.B(n_458),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1788),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1788),
.Y(n_2202)
);

A2O1A1Ixp33_ASAP7_75t_L g2203 ( 
.A1(n_1997),
.A2(n_461),
.B(n_459),
.C(n_460),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1737),
.B(n_459),
.Y(n_2204)
);

INVxp67_ASAP7_75t_SL g2205 ( 
.A(n_1760),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_1773),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_1778),
.B(n_462),
.Y(n_2207)
);

OAI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_1828),
.A2(n_462),
.B(n_463),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_1760),
.Y(n_2209)
);

AOI21xp5_ASAP7_75t_SL g2210 ( 
.A1(n_1737),
.A2(n_464),
.B(n_466),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1780),
.B(n_468),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1782),
.B(n_468),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_1997),
.B(n_469),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_2006),
.B(n_470),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2006),
.B(n_471),
.Y(n_2215)
);

AOI21xp5_ASAP7_75t_SL g2216 ( 
.A1(n_2008),
.A2(n_472),
.B(n_473),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1760),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_1954),
.A2(n_475),
.B(n_476),
.Y(n_2218)
);

A2O1A1Ixp33_ASAP7_75t_L g2219 ( 
.A1(n_2008),
.A2(n_2018),
.B(n_2017),
.C(n_1816),
.Y(n_2219)
);

OAI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1805),
.A2(n_1841),
.B(n_1839),
.Y(n_2220)
);

INVx1_ASAP7_75t_SL g2221 ( 
.A(n_1774),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1856),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_1928),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_2223)
);

AO31x2_ASAP7_75t_L g2224 ( 
.A1(n_2017),
.A2(n_477),
.A3(n_478),
.B(n_480),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_2018),
.B(n_480),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_1898),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_1753),
.B(n_481),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1801),
.B(n_482),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1804),
.B(n_483),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1776),
.B(n_484),
.Y(n_2230)
);

AO31x2_ASAP7_75t_L g2231 ( 
.A1(n_1840),
.A2(n_486),
.A3(n_487),
.B(n_489),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1832),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1786),
.B(n_489),
.Y(n_2233)
);

AOI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_1864),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_1800),
.Y(n_2235)
);

NAND2x1p5_ASAP7_75t_L g2236 ( 
.A(n_1900),
.B(n_493),
.Y(n_2236)
);

CKINVDCx16_ASAP7_75t_R g2237 ( 
.A(n_1802),
.Y(n_2237)
);

NOR2xp67_ASAP7_75t_SL g2238 ( 
.A(n_1870),
.B(n_1873),
.Y(n_2238)
);

INVx5_ASAP7_75t_L g2239 ( 
.A(n_1727),
.Y(n_2239)
);

INVx4_ASAP7_75t_L g2240 ( 
.A(n_1832),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_1754),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1838),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1724),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_1767),
.Y(n_2244)
);

AOI221x1_ASAP7_75t_L g2245 ( 
.A1(n_1840),
.A2(n_1867),
.B1(n_1843),
.B2(n_1889),
.C(n_1885),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_1930),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_2246)
);

BUFx2_ASAP7_75t_L g2247 ( 
.A(n_1861),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1826),
.Y(n_2248)
);

OR2x6_ASAP7_75t_L g2249 ( 
.A(n_1758),
.B(n_502),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1820),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1875),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_1962),
.A2(n_505),
.B(n_507),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1807),
.B(n_509),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_1971),
.A2(n_511),
.B(n_512),
.Y(n_2254)
);

AO32x2_ASAP7_75t_L g2255 ( 
.A1(n_1838),
.A2(n_514),
.A3(n_515),
.B1(n_516),
.B2(n_517),
.Y(n_2255)
);

AO31x2_ASAP7_75t_L g2256 ( 
.A1(n_1843),
.A2(n_514),
.A3(n_515),
.B(n_516),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1759),
.B(n_518),
.Y(n_2257)
);

BUFx2_ASAP7_75t_L g2258 ( 
.A(n_1779),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1876),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_SL g2260 ( 
.A(n_1859),
.B(n_520),
.C(n_523),
.Y(n_2260)
);

AO31x2_ASAP7_75t_L g2261 ( 
.A1(n_1867),
.A2(n_523),
.A3(n_524),
.B(n_525),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1894),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_1723),
.B(n_525),
.Y(n_2263)
);

NOR2xp67_ASAP7_75t_L g2264 ( 
.A(n_1730),
.B(n_528),
.Y(n_2264)
);

AO32x2_ASAP7_75t_L g2265 ( 
.A1(n_1885),
.A2(n_528),
.A3(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_2265)
);

AO21x2_ASAP7_75t_L g2266 ( 
.A1(n_1892),
.A2(n_529),
.B(n_532),
.Y(n_2266)
);

INVx3_ASAP7_75t_L g2267 ( 
.A(n_1735),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1781),
.B(n_533),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1879),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1975),
.B(n_1976),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_1733),
.B(n_537),
.Y(n_2271)
);

AO31x2_ASAP7_75t_L g2272 ( 
.A1(n_1889),
.A2(n_538),
.A3(n_539),
.B(n_540),
.Y(n_2272)
);

NOR2xp67_ASAP7_75t_L g2273 ( 
.A(n_1725),
.B(n_540),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_1985),
.A2(n_541),
.B(n_542),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1880),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_1819),
.B(n_543),
.Y(n_2276)
);

BUFx6f_ASAP7_75t_L g2277 ( 
.A(n_1797),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_1935),
.B(n_547),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2120),
.B(n_1882),
.Y(n_2279)
);

INVx1_ASAP7_75t_SL g2280 ( 
.A(n_2090),
.Y(n_2280)
);

INVx8_ASAP7_75t_L g2281 ( 
.A(n_2077),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2029),
.B(n_1729),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2042),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2047),
.Y(n_2284)
);

OR3x4_ASAP7_75t_SL g2285 ( 
.A(n_2078),
.B(n_548),
.C(n_549),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2030),
.B(n_1937),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2181),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2069),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_2239),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2094),
.A2(n_1815),
.B1(n_1809),
.B2(n_1812),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2181),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2096),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2091),
.B(n_1938),
.Y(n_2293)
);

BUFx2_ASAP7_75t_L g2294 ( 
.A(n_2069),
.Y(n_2294)
);

O2A1O1Ixp33_ASAP7_75t_SL g2295 ( 
.A1(n_2219),
.A2(n_1940),
.B(n_1943),
.C(n_1942),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2045),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2185),
.Y(n_2297)
);

O2A1O1Ixp33_ASAP7_75t_L g2298 ( 
.A1(n_2026),
.A2(n_2016),
.B(n_1944),
.C(n_1946),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2146),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_2239),
.Y(n_2300)
);

AOI22xp33_ASAP7_75t_L g2301 ( 
.A1(n_2147),
.A2(n_1814),
.B1(n_1803),
.B2(n_1844),
.Y(n_2301)
);

CKINVDCx11_ASAP7_75t_R g2302 ( 
.A(n_2164),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2071),
.A2(n_1947),
.B1(n_1948),
.B2(n_1945),
.Y(n_2303)
);

INVx1_ASAP7_75t_SL g2304 ( 
.A(n_2115),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2239),
.Y(n_2305)
);

NAND2x1p5_ASAP7_75t_L g2306 ( 
.A(n_2024),
.B(n_1949),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2036),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2036),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2053),
.Y(n_2309)
);

OA21x2_ASAP7_75t_L g2310 ( 
.A1(n_2245),
.A2(n_1854),
.B(n_1852),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2099),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2131),
.B(n_1836),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2170),
.B(n_1837),
.Y(n_2313)
);

AO21x2_ASAP7_75t_L g2314 ( 
.A1(n_2073),
.A2(n_1855),
.B(n_1825),
.Y(n_2314)
);

CKINVDCx8_ASAP7_75t_R g2315 ( 
.A(n_2135),
.Y(n_2315)
);

INVx3_ASAP7_75t_SL g2316 ( 
.A(n_2119),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2053),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2024),
.B(n_1950),
.Y(n_2318)
);

CKINVDCx16_ASAP7_75t_R g2319 ( 
.A(n_2237),
.Y(n_2319)
);

NAND2x1p5_ASAP7_75t_L g2320 ( 
.A(n_2057),
.B(n_1951),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2022),
.A2(n_2014),
.B1(n_2012),
.B2(n_2011),
.Y(n_2321)
);

BUFx2_ASAP7_75t_SL g2322 ( 
.A(n_2057),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2076),
.A2(n_1845),
.B1(n_1846),
.B2(n_1848),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_2064),
.Y(n_2324)
);

OAI22xp33_ASAP7_75t_L g2325 ( 
.A1(n_2048),
.A2(n_1966),
.B1(n_2009),
.B2(n_2005),
.Y(n_2325)
);

NOR2xp67_ASAP7_75t_SL g2326 ( 
.A(n_2210),
.B(n_1952),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_2241),
.Y(n_2327)
);

OAI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_2140),
.A2(n_1957),
.B(n_1956),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_2081),
.B(n_1868),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2076),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_SL g2331 ( 
.A(n_2240),
.B(n_1891),
.Y(n_2331)
);

INVx3_ASAP7_75t_SL g2332 ( 
.A(n_2168),
.Y(n_2332)
);

OAI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2117),
.A2(n_1969),
.B1(n_2003),
.B2(n_2002),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_2243),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2070),
.Y(n_2335)
);

INVxp67_ASAP7_75t_SL g2336 ( 
.A(n_2064),
.Y(n_2336)
);

NAND2xp33_ASAP7_75t_SL g2337 ( 
.A(n_2082),
.B(n_1960),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2020),
.Y(n_2338)
);

INVx2_ASAP7_75t_SL g2339 ( 
.A(n_2159),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2072),
.B(n_1963),
.Y(n_2340)
);

AOI21xp33_ASAP7_75t_L g2341 ( 
.A1(n_2027),
.A2(n_1965),
.B(n_1964),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2240),
.A2(n_2010),
.B1(n_2001),
.B2(n_2000),
.Y(n_2342)
);

AO21x1_ASAP7_75t_L g2343 ( 
.A1(n_2213),
.A2(n_1891),
.B(n_1850),
.Y(n_2343)
);

BUFx12f_ASAP7_75t_L g2344 ( 
.A(n_2158),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2159),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2112),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2098),
.B(n_1970),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2087),
.B(n_1972),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2107),
.B(n_1973),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2154),
.Y(n_2350)
);

BUFx3_ASAP7_75t_L g2351 ( 
.A(n_2051),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2051),
.Y(n_2352)
);

OR2x6_ASAP7_75t_L g2353 ( 
.A(n_2082),
.B(n_1979),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2116),
.B(n_1980),
.Y(n_2354)
);

OA21x2_ASAP7_75t_L g2355 ( 
.A1(n_2232),
.A2(n_1982),
.B(n_1981),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2051),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2059),
.B(n_1765),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_2136),
.Y(n_2358)
);

OAI21x1_ASAP7_75t_L g2359 ( 
.A1(n_2232),
.A2(n_1987),
.B(n_1983),
.Y(n_2359)
);

OR2x6_ASAP7_75t_L g2360 ( 
.A(n_2082),
.B(n_1988),
.Y(n_2360)
);

INVx2_ASAP7_75t_SL g2361 ( 
.A(n_2136),
.Y(n_2361)
);

BUFx8_ASAP7_75t_SL g2362 ( 
.A(n_2249),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2100),
.B(n_1991),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2149),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2160),
.B(n_1851),
.C(n_1865),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2226),
.B(n_1738),
.Y(n_2366)
);

OAI21x1_ASAP7_75t_L g2367 ( 
.A1(n_2242),
.A2(n_1994),
.B(n_1993),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2122),
.B(n_1995),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2149),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2193),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2103),
.Y(n_2371)
);

INVx1_ASAP7_75t_SL g2372 ( 
.A(n_2103),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_2193),
.Y(n_2373)
);

AOI21x1_ASAP7_75t_L g2374 ( 
.A1(n_2270),
.A2(n_1998),
.B(n_1798),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2132),
.B(n_548),
.Y(n_2375)
);

BUFx2_ASAP7_75t_L g2376 ( 
.A(n_2052),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2193),
.B(n_1735),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2221),
.B(n_1853),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2093),
.A2(n_1857),
.B(n_1893),
.C(n_1884),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2106),
.B(n_1790),
.Y(n_2380)
);

BUFx8_ASAP7_75t_SL g2381 ( 
.A(n_2249),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2133),
.B(n_549),
.Y(n_2382)
);

OA21x2_ASAP7_75t_L g2383 ( 
.A1(n_2194),
.A2(n_1789),
.B(n_551),
.Y(n_2383)
);

O2A1O1Ixp33_ASAP7_75t_SL g2384 ( 
.A1(n_2198),
.A2(n_550),
.B(n_552),
.C(n_553),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2114),
.A2(n_550),
.B1(n_552),
.B2(n_553),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2118),
.B(n_554),
.Y(n_2386)
);

OAI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2088),
.A2(n_555),
.B1(n_556),
.B2(n_557),
.Y(n_2387)
);

AOI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2182),
.A2(n_556),
.B(n_557),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2028),
.B(n_558),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_SL g2390 ( 
.A1(n_2056),
.A2(n_560),
.B(n_563),
.Y(n_2390)
);

NAND3xp33_ASAP7_75t_L g2391 ( 
.A(n_2163),
.B(n_564),
.C(n_566),
.Y(n_2391)
);

O2A1O1Ixp33_ASAP7_75t_L g2392 ( 
.A1(n_2067),
.A2(n_567),
.B(n_568),
.C(n_570),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2083),
.B(n_2134),
.Y(n_2393)
);

NAND2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2258),
.B(n_573),
.Y(n_2394)
);

OR2x6_ASAP7_75t_SL g2395 ( 
.A(n_2041),
.B(n_576),
.Y(n_2395)
);

NAND2x1p5_ASAP7_75t_L g2396 ( 
.A(n_2183),
.B(n_577),
.Y(n_2396)
);

OR2x2_ASAP7_75t_SL g2397 ( 
.A(n_2260),
.B(n_577),
.Y(n_2397)
);

NOR2xp67_ASAP7_75t_L g2398 ( 
.A(n_2267),
.B(n_579),
.Y(n_2398)
);

INVxp33_ASAP7_75t_L g2399 ( 
.A(n_2238),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2217),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2149),
.Y(n_2401)
);

NAND2x1p5_ASAP7_75t_L g2402 ( 
.A(n_2141),
.B(n_581),
.Y(n_2402)
);

OAI211xp5_ASAP7_75t_L g2403 ( 
.A1(n_2125),
.A2(n_2040),
.B(n_2145),
.C(n_2097),
.Y(n_2403)
);

AOI21xp33_ASAP7_75t_L g2404 ( 
.A1(n_2033),
.A2(n_582),
.B(n_583),
.Y(n_2404)
);

NOR2x1_ASAP7_75t_L g2405 ( 
.A(n_2050),
.B(n_583),
.Y(n_2405)
);

OAI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2037),
.A2(n_584),
.B(n_585),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2046),
.B(n_584),
.Y(n_2407)
);

NOR2xp67_ASAP7_75t_L g2408 ( 
.A(n_2173),
.B(n_585),
.Y(n_2408)
);

OR2x6_ASAP7_75t_L g2409 ( 
.A(n_2065),
.B(n_586),
.Y(n_2409)
);

A2O1A1Ixp33_ASAP7_75t_L g2410 ( 
.A1(n_2128),
.A2(n_587),
.B(n_588),
.C(n_589),
.Y(n_2410)
);

OAI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2200),
.A2(n_587),
.B(n_589),
.Y(n_2411)
);

INVx4_ASAP7_75t_SL g2412 ( 
.A(n_2199),
.Y(n_2412)
);

BUFx3_ASAP7_75t_L g2413 ( 
.A(n_2141),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2191),
.B(n_2192),
.Y(n_2414)
);

OAI221xp5_ASAP7_75t_L g2415 ( 
.A1(n_2111),
.A2(n_660),
.B1(n_591),
.B2(n_592),
.C(n_593),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_2205),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2191),
.B(n_590),
.Y(n_2417)
);

AO21x2_ASAP7_75t_L g2418 ( 
.A1(n_2095),
.A2(n_596),
.B(n_597),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_2144),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2244),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2061),
.A2(n_598),
.B1(n_600),
.B2(n_601),
.Y(n_2421)
);

BUFx12f_ASAP7_75t_L g2422 ( 
.A(n_2206),
.Y(n_2422)
);

BUFx12f_ASAP7_75t_L g2423 ( 
.A(n_2171),
.Y(n_2423)
);

INVx5_ASAP7_75t_L g2424 ( 
.A(n_2144),
.Y(n_2424)
);

NAND2x1p5_ASAP7_75t_L g2425 ( 
.A(n_2150),
.B(n_602),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2102),
.Y(n_2426)
);

CKINVDCx11_ASAP7_75t_R g2427 ( 
.A(n_2166),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2102),
.Y(n_2428)
);

AND2x4_ASAP7_75t_L g2429 ( 
.A(n_2192),
.B(n_603),
.Y(n_2429)
);

BUFx3_ASAP7_75t_L g2430 ( 
.A(n_2209),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2263),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_2247),
.B(n_604),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2058),
.Y(n_2433)
);

AO21x2_ASAP7_75t_L g2434 ( 
.A1(n_2105),
.A2(n_605),
.B(n_606),
.Y(n_2434)
);

OR2x2_ASAP7_75t_L g2435 ( 
.A(n_2155),
.B(n_606),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2207),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2143),
.A2(n_609),
.B(n_610),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2197),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2186),
.B(n_611),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2184),
.Y(n_2440)
);

AO21x2_ASAP7_75t_L g2441 ( 
.A1(n_2130),
.A2(n_616),
.B(n_617),
.Y(n_2441)
);

CKINVDCx6p67_ASAP7_75t_R g2442 ( 
.A(n_2175),
.Y(n_2442)
);

AOI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2235),
.A2(n_616),
.B1(n_618),
.B2(n_619),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2139),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2201),
.B(n_620),
.Y(n_2445)
);

OAI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2220),
.A2(n_621),
.B(n_622),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2214),
.A2(n_623),
.B(n_624),
.Y(n_2447)
);

AOI22xp33_ASAP7_75t_L g2448 ( 
.A1(n_2032),
.A2(n_623),
.B1(n_625),
.B2(n_627),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2138),
.A2(n_629),
.B1(n_630),
.B2(n_631),
.Y(n_2449)
);

AND2x4_ASAP7_75t_L g2450 ( 
.A(n_2201),
.B(n_632),
.Y(n_2450)
);

AO21x2_ASAP7_75t_L g2451 ( 
.A1(n_2035),
.A2(n_633),
.B(n_634),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2202),
.B(n_633),
.Y(n_2452)
);

OAI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_2189),
.A2(n_635),
.B(n_636),
.Y(n_2453)
);

AO22x2_ASAP7_75t_L g2454 ( 
.A1(n_2089),
.A2(n_2215),
.B1(n_2225),
.B2(n_2085),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2023),
.Y(n_2455)
);

AND2x6_ASAP7_75t_L g2456 ( 
.A(n_2202),
.B(n_638),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2187),
.B(n_642),
.Y(n_2457)
);

O2A1O1Ixp33_ASAP7_75t_SL g2458 ( 
.A1(n_2203),
.A2(n_643),
.B(n_644),
.C(n_645),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2137),
.Y(n_2459)
);

AOI22xp33_ASAP7_75t_L g2460 ( 
.A1(n_2162),
.A2(n_643),
.B1(n_645),
.B2(n_646),
.Y(n_2460)
);

OR2x6_ASAP7_75t_L g2461 ( 
.A(n_2075),
.B(n_647),
.Y(n_2461)
);

INVx2_ASAP7_75t_SL g2462 ( 
.A(n_2271),
.Y(n_2462)
);

OA21x2_ASAP7_75t_L g2463 ( 
.A1(n_2074),
.A2(n_647),
.B(n_648),
.Y(n_2463)
);

OAI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2152),
.A2(n_648),
.B(n_649),
.Y(n_2464)
);

OAI21x1_ASAP7_75t_SL g2465 ( 
.A1(n_2056),
.A2(n_650),
.B(n_651),
.Y(n_2465)
);

INVx2_ASAP7_75t_SL g2466 ( 
.A(n_2271),
.Y(n_2466)
);

BUFx8_ASAP7_75t_L g2467 ( 
.A(n_2129),
.Y(n_2467)
);

OAI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2177),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_2468)
);

OAI221xp5_ASAP7_75t_L g2469 ( 
.A1(n_2165),
.A2(n_2104),
.B1(n_2124),
.B2(n_2039),
.C(n_2157),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2188),
.B(n_656),
.Y(n_2470)
);

AOI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2068),
.A2(n_657),
.B1(n_658),
.B2(n_659),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2092),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2025),
.B(n_2080),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2257),
.B(n_2253),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2062),
.B(n_2262),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_2209),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2054),
.B(n_2250),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_2063),
.A2(n_2110),
.B(n_2079),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_2227),
.Y(n_2479)
);

AOI22xp33_ASAP7_75t_L g2480 ( 
.A1(n_2251),
.A2(n_2275),
.B1(n_2269),
.B2(n_2259),
.Y(n_2480)
);

AOI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2034),
.A2(n_2195),
.B(n_2178),
.Y(n_2481)
);

AO31x2_ASAP7_75t_L g2482 ( 
.A1(n_2127),
.A2(n_2196),
.A3(n_2054),
.B(n_2274),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2231),
.Y(n_2483)
);

OA21x2_ASAP7_75t_L g2484 ( 
.A1(n_2123),
.A2(n_2126),
.B(n_2180),
.Y(n_2484)
);

OA21x2_ASAP7_75t_L g2485 ( 
.A1(n_2179),
.A2(n_2252),
.B(n_2254),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2276),
.B(n_2264),
.Y(n_2486)
);

O2A1O1Ixp33_ASAP7_75t_L g2487 ( 
.A1(n_2142),
.A2(n_2148),
.B(n_2151),
.C(n_2167),
.Y(n_2487)
);

AOI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2204),
.A2(n_2049),
.B(n_2218),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2256),
.Y(n_2489)
);

O2A1O1Ixp33_ASAP7_75t_L g2490 ( 
.A1(n_2153),
.A2(n_2161),
.B(n_2230),
.C(n_2233),
.Y(n_2490)
);

CKINVDCx20_ASAP7_75t_R g2491 ( 
.A(n_2211),
.Y(n_2491)
);

NAND2x1p5_ASAP7_75t_L g2492 ( 
.A(n_2273),
.B(n_2262),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2236),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2248),
.B(n_2262),
.Y(n_2494)
);

AOI22xp33_ASAP7_75t_L g2495 ( 
.A1(n_2101),
.A2(n_2055),
.B1(n_2208),
.B2(n_2278),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2212),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2222),
.B(n_2277),
.Y(n_2497)
);

OAI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2156),
.A2(n_2031),
.B1(n_2234),
.B2(n_2216),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2302),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2459),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2416),
.Y(n_2501)
);

BUFx8_ASAP7_75t_SL g2502 ( 
.A(n_2350),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2344),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2289),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_2362),
.Y(n_2505)
);

OAI21xp5_ASAP7_75t_L g2506 ( 
.A1(n_2391),
.A2(n_2066),
.B(n_2060),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2477),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2289),
.B(n_2224),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2431),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2299),
.Y(n_2510)
);

BUFx2_ASAP7_75t_L g2511 ( 
.A(n_2294),
.Y(n_2511)
);

BUFx12f_ASAP7_75t_L g2512 ( 
.A(n_2288),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2435),
.B(n_2021),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2436),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2376),
.B(n_2021),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2338),
.Y(n_2516)
);

INVx2_ASAP7_75t_SL g2517 ( 
.A(n_2281),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2440),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2283),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2311),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2375),
.B(n_2129),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2284),
.Y(n_2522)
);

OR2x6_ASAP7_75t_L g2523 ( 
.A(n_2322),
.B(n_2121),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2382),
.B(n_2129),
.Y(n_2524)
);

INVx5_ASAP7_75t_SL g2525 ( 
.A(n_2442),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2287),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2291),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2300),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2300),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2297),
.Y(n_2530)
);

OR2x6_ASAP7_75t_L g2531 ( 
.A(n_2281),
.B(n_2222),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2345),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2417),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2305),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2439),
.B(n_2043),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2417),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2281),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2483),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2305),
.B(n_2224),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2414),
.B(n_2021),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2489),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2429),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2429),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2445),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2444),
.Y(n_2545)
);

AOI22xp33_ASAP7_75t_L g2546 ( 
.A1(n_2427),
.A2(n_2113),
.B1(n_2108),
.B2(n_2109),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2351),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2474),
.B(n_2043),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2419),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2450),
.Y(n_2550)
);

INVx3_ASAP7_75t_L g2551 ( 
.A(n_2419),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2414),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2452),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2282),
.B(n_2190),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2393),
.B(n_2319),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2457),
.B(n_2190),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2452),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2409),
.A2(n_2084),
.B1(n_2038),
.B2(n_2044),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2327),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2386),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2470),
.B(n_2347),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2412),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_2412),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2386),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_2346),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2349),
.B(n_2190),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2389),
.Y(n_2567)
);

INVxp67_ASAP7_75t_SL g2568 ( 
.A(n_2331),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2389),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2407),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2407),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_SL g2572 ( 
.A1(n_2467),
.A2(n_2223),
.B1(n_2246),
.B2(n_2277),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2316),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2340),
.B(n_2169),
.Y(n_2574)
);

BUFx2_ASAP7_75t_L g2575 ( 
.A(n_2352),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2319),
.B(n_2176),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_2373),
.B(n_2224),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2280),
.B(n_2272),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_2423),
.Y(n_2579)
);

NAND2xp33_ASAP7_75t_R g2580 ( 
.A(n_2383),
.B(n_2268),
.Y(n_2580)
);

OA21x2_ASAP7_75t_L g2581 ( 
.A1(n_2364),
.A2(n_2401),
.B(n_2369),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2356),
.Y(n_2582)
);

AOI22xp33_ASAP7_75t_L g2583 ( 
.A1(n_2409),
.A2(n_2086),
.B1(n_2229),
.B2(n_2228),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2354),
.B(n_2176),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2373),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_2381),
.Y(n_2586)
);

BUFx5_ASAP7_75t_L g2587 ( 
.A(n_2456),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2395),
.B(n_2172),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2330),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2307),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2308),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2358),
.Y(n_2592)
);

CKINVDCx10_ASAP7_75t_R g2593 ( 
.A(n_2409),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2309),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2368),
.B(n_2176),
.Y(n_2595)
);

INVx1_ASAP7_75t_SL g2596 ( 
.A(n_2280),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2426),
.B(n_2428),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2317),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2377),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2462),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2466),
.Y(n_2601)
);

INVx5_ASAP7_75t_L g2602 ( 
.A(n_2456),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2336),
.B(n_2272),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2388),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2456),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2456),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2486),
.B(n_2255),
.Y(n_2607)
);

BUFx12f_ASAP7_75t_SL g2608 ( 
.A(n_2461),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2339),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2473),
.B(n_2174),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2424),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2472),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2324),
.B(n_2256),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2424),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2398),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_2461),
.A2(n_2266),
.B1(n_2277),
.B2(n_2222),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2324),
.B(n_2261),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2421),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2421),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2334),
.Y(n_2620)
);

OR2x6_ASAP7_75t_L g2621 ( 
.A(n_2461),
.B(n_2255),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_2370),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2402),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2400),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2399),
.B(n_2255),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2286),
.B(n_2265),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_2331),
.A2(n_2265),
.B(n_2261),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2425),
.Y(n_2628)
);

AND2x2_ASAP7_75t_L g2629 ( 
.A(n_2455),
.B(n_2265),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2424),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2418),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2434),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2335),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2441),
.Y(n_2634)
);

BUFx3_ASAP7_75t_L g2635 ( 
.A(n_2413),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2430),
.Y(n_2636)
);

HB1xp67_ASAP7_75t_L g2637 ( 
.A(n_2304),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2304),
.B(n_2433),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2292),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2361),
.Y(n_2640)
);

BUFx4f_ASAP7_75t_L g2641 ( 
.A(n_2394),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2441),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2438),
.B(n_2496),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2296),
.B(n_2437),
.Y(n_2644)
);

HB1xp67_ASAP7_75t_L g2645 ( 
.A(n_2371),
.Y(n_2645)
);

CKINVDCx6p67_ASAP7_75t_R g2646 ( 
.A(n_2332),
.Y(n_2646)
);

AOI21x1_ASAP7_75t_L g2647 ( 
.A1(n_2488),
.A2(n_2343),
.B(n_2408),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2279),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2385),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2467),
.A2(n_2498),
.B1(n_2415),
.B2(n_2469),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2372),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2385),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2312),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2312),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2313),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2313),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2446),
.Y(n_2657)
);

BUFx10_ASAP7_75t_L g2658 ( 
.A(n_2517),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2561),
.B(n_2494),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2602),
.B(n_2587),
.Y(n_2660)
);

NAND2xp33_ASAP7_75t_R g2661 ( 
.A(n_2505),
.B(n_2420),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_R g2662 ( 
.A(n_2608),
.B(n_2315),
.Y(n_2662)
);

BUFx10_ASAP7_75t_L g2663 ( 
.A(n_2537),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_2502),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2509),
.B(n_2480),
.Y(n_2665)
);

NAND2xp33_ASAP7_75t_R g2666 ( 
.A(n_2505),
.B(n_2285),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2510),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2514),
.B(n_2495),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_R g2669 ( 
.A(n_2593),
.B(n_2422),
.Y(n_2669)
);

XNOR2xp5_ASAP7_75t_L g2670 ( 
.A(n_2499),
.B(n_2491),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2518),
.B(n_2454),
.Y(n_2671)
);

NOR2xp33_ASAP7_75t_R g2672 ( 
.A(n_2593),
.B(n_2479),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2501),
.B(n_2497),
.Y(n_2673)
);

NAND2xp33_ASAP7_75t_R g2674 ( 
.A(n_2586),
.B(n_2378),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2501),
.B(n_2497),
.Y(n_2675)
);

NAND2xp33_ASAP7_75t_R g2676 ( 
.A(n_2586),
.B(n_2293),
.Y(n_2676)
);

NAND2xp33_ASAP7_75t_R g2677 ( 
.A(n_2511),
.B(n_2478),
.Y(n_2677)
);

NAND2xp33_ASAP7_75t_R g2678 ( 
.A(n_2503),
.B(n_2523),
.Y(n_2678)
);

INVxp67_ASAP7_75t_L g2679 ( 
.A(n_2637),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2519),
.B(n_2454),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2522),
.B(n_2494),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2500),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2602),
.B(n_2493),
.Y(n_2683)
);

CKINVDCx16_ASAP7_75t_R g2684 ( 
.A(n_2499),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2502),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2596),
.B(n_2476),
.Y(n_2686)
);

NAND2xp33_ASAP7_75t_R g2687 ( 
.A(n_2523),
.B(n_2318),
.Y(n_2687)
);

AND2x2_ASAP7_75t_L g2688 ( 
.A(n_2596),
.B(n_2476),
.Y(n_2688)
);

AND2x2_ASAP7_75t_SL g2689 ( 
.A(n_2641),
.B(n_2290),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_R g2690 ( 
.A(n_2646),
.B(n_2337),
.Y(n_2690)
);

CKINVDCx11_ASAP7_75t_R g2691 ( 
.A(n_2512),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2637),
.Y(n_2692)
);

INVxp67_ASAP7_75t_L g2693 ( 
.A(n_2633),
.Y(n_2693)
);

AND2x4_ASAP7_75t_L g2694 ( 
.A(n_2602),
.B(n_2329),
.Y(n_2694)
);

NAND2xp33_ASAP7_75t_R g2695 ( 
.A(n_2523),
.B(n_2549),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2633),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2589),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2576),
.B(n_2451),
.Y(n_2698)
);

NAND2xp33_ASAP7_75t_R g2699 ( 
.A(n_2549),
.B(n_2366),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2590),
.Y(n_2700)
);

NAND2xp33_ASAP7_75t_SL g2701 ( 
.A(n_2650),
.B(n_2323),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2591),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_2579),
.Y(n_2703)
);

NAND2xp33_ASAP7_75t_R g2704 ( 
.A(n_2551),
.B(n_2446),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2585),
.Y(n_2705)
);

INVxp67_ASAP7_75t_L g2706 ( 
.A(n_2532),
.Y(n_2706)
);

CKINVDCx16_ASAP7_75t_R g2707 ( 
.A(n_2532),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2638),
.B(n_2451),
.Y(n_2708)
);

OR2x6_ASAP7_75t_L g2709 ( 
.A(n_2531),
.B(n_2492),
.Y(n_2709)
);

NAND2xp33_ASAP7_75t_SL g2710 ( 
.A(n_2650),
.B(n_2551),
.Y(n_2710)
);

NAND2xp33_ASAP7_75t_R g2711 ( 
.A(n_2643),
.B(n_2484),
.Y(n_2711)
);

NAND2xp33_ASAP7_75t_R g2712 ( 
.A(n_2531),
.B(n_2484),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2548),
.B(n_2355),
.Y(n_2713)
);

NAND2xp33_ASAP7_75t_R g2714 ( 
.A(n_2531),
.B(n_2453),
.Y(n_2714)
);

NAND2xp33_ASAP7_75t_R g2715 ( 
.A(n_2621),
.B(n_2453),
.Y(n_2715)
);

NAND2xp33_ASAP7_75t_R g2716 ( 
.A(n_2621),
.B(n_2463),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_R g2717 ( 
.A(n_2621),
.B(n_2588),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_R g2718 ( 
.A(n_2641),
.B(n_2357),
.Y(n_2718)
);

BUFx10_ASAP7_75t_L g2719 ( 
.A(n_2573),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2525),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2516),
.Y(n_2721)
);

NAND2xp33_ASAP7_75t_R g2722 ( 
.A(n_2588),
.B(n_2463),
.Y(n_2722)
);

INVxp33_ASAP7_75t_L g2723 ( 
.A(n_2636),
.Y(n_2723)
);

NAND2xp33_ASAP7_75t_R g2724 ( 
.A(n_2611),
.B(n_2406),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2599),
.B(n_2475),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2594),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2599),
.B(n_2526),
.Y(n_2727)
);

NAND2xp33_ASAP7_75t_R g2728 ( 
.A(n_2611),
.B(n_2406),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2644),
.B(n_2355),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2527),
.B(n_2408),
.Y(n_2730)
);

INVx5_ASAP7_75t_L g2731 ( 
.A(n_2525),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2598),
.Y(n_2732)
);

XNOR2xp5_ASAP7_75t_L g2733 ( 
.A(n_2639),
.B(n_2498),
.Y(n_2733)
);

INVxp67_ASAP7_75t_L g2734 ( 
.A(n_2609),
.Y(n_2734)
);

XNOR2xp5_ASAP7_75t_L g2735 ( 
.A(n_2559),
.B(n_2620),
.Y(n_2735)
);

OR2x4_ASAP7_75t_L g2736 ( 
.A(n_2555),
.B(n_2625),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2530),
.Y(n_2737)
);

NAND2xp33_ASAP7_75t_SL g2738 ( 
.A(n_2513),
.B(n_2326),
.Y(n_2738)
);

NAND2xp33_ASAP7_75t_R g2739 ( 
.A(n_2614),
.B(n_2411),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_SL g2740 ( 
.A(n_2587),
.B(n_2403),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2507),
.Y(n_2741)
);

INVx2_ASAP7_75t_SL g2742 ( 
.A(n_2609),
.Y(n_2742)
);

CKINVDCx20_ASAP7_75t_R g2743 ( 
.A(n_2525),
.Y(n_2743)
);

BUFx3_ASAP7_75t_L g2744 ( 
.A(n_2635),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2520),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_R g2746 ( 
.A(n_2587),
.B(n_2374),
.Y(n_2746)
);

XNOR2xp5_ASAP7_75t_L g2747 ( 
.A(n_2546),
.B(n_2397),
.Y(n_2747)
);

NAND2xp33_ASAP7_75t_R g2748 ( 
.A(n_2614),
.B(n_2411),
.Y(n_2748)
);

INVxp67_ASAP7_75t_L g2749 ( 
.A(n_2547),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2552),
.B(n_2405),
.Y(n_2750)
);

NAND2xp33_ASAP7_75t_R g2751 ( 
.A(n_2630),
.B(n_2310),
.Y(n_2751)
);

NAND2xp33_ASAP7_75t_R g2752 ( 
.A(n_2630),
.B(n_2310),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2508),
.B(n_2353),
.Y(n_2753)
);

AND2x4_ASAP7_75t_L g2754 ( 
.A(n_2508),
.B(n_2353),
.Y(n_2754)
);

NAND2xp33_ASAP7_75t_R g2755 ( 
.A(n_2575),
.B(n_2485),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2600),
.B(n_2405),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2648),
.B(n_2363),
.Y(n_2757)
);

INVxp67_ASAP7_75t_L g2758 ( 
.A(n_2582),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2601),
.B(n_2380),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_2635),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_2636),
.Y(n_2761)
);

XNOR2xp5_ASAP7_75t_L g2762 ( 
.A(n_2546),
.B(n_2396),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2539),
.B(n_2360),
.Y(n_2763)
);

INVxp67_ASAP7_75t_L g2764 ( 
.A(n_2592),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2607),
.B(n_2554),
.Y(n_2765)
);

XOR2x2_ASAP7_75t_SL g2766 ( 
.A(n_2572),
.B(n_2468),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2539),
.B(n_2360),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2622),
.Y(n_2768)
);

NAND2xp33_ASAP7_75t_SL g2769 ( 
.A(n_2515),
.B(n_2301),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2566),
.B(n_2482),
.Y(n_2770)
);

BUFx3_ASAP7_75t_L g2771 ( 
.A(n_2622),
.Y(n_2771)
);

XNOR2xp5_ASAP7_75t_L g2772 ( 
.A(n_2572),
.B(n_2468),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2538),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2584),
.B(n_2482),
.Y(n_2774)
);

NAND2xp33_ASAP7_75t_R g2775 ( 
.A(n_2504),
.B(n_2360),
.Y(n_2775)
);

AND2x4_ASAP7_75t_L g2776 ( 
.A(n_2613),
.B(n_2314),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2595),
.B(n_2482),
.Y(n_2777)
);

INVxp67_ASAP7_75t_L g2778 ( 
.A(n_2624),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_R g2779 ( 
.A(n_2624),
.B(n_2448),
.Y(n_2779)
);

INVxp67_ASAP7_75t_L g2780 ( 
.A(n_2645),
.Y(n_2780)
);

NAND2xp33_ASAP7_75t_R g2781 ( 
.A(n_2528),
.B(n_2464),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2521),
.B(n_2314),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2613),
.B(n_2359),
.Y(n_2783)
);

XNOR2xp5_ASAP7_75t_L g2784 ( 
.A(n_2524),
.B(n_2387),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2556),
.B(n_2367),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_R g2786 ( 
.A(n_2623),
.B(n_2471),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_2645),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2653),
.B(n_2363),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_R g2789 ( 
.A(n_2628),
.B(n_2443),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2617),
.B(n_2577),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_R g2791 ( 
.A(n_2528),
.B(n_2449),
.Y(n_2791)
);

INVxp67_ASAP7_75t_L g2792 ( 
.A(n_2651),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2654),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_R g2794 ( 
.A(n_2529),
.B(n_2348),
.Y(n_2794)
);

XNOR2xp5_ASAP7_75t_L g2795 ( 
.A(n_2535),
.B(n_2306),
.Y(n_2795)
);

NAND2xp33_ASAP7_75t_R g2796 ( 
.A(n_2534),
.B(n_2629),
.Y(n_2796)
);

OR2x2_ASAP7_75t_L g2797 ( 
.A(n_2655),
.B(n_2432),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2640),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2656),
.Y(n_2799)
);

CKINVDCx16_ASAP7_75t_R g2800 ( 
.A(n_2640),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2533),
.B(n_2341),
.Y(n_2801)
);

HB1xp67_ASAP7_75t_L g2802 ( 
.A(n_2651),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2597),
.Y(n_2803)
);

NAND2xp33_ASAP7_75t_R g2804 ( 
.A(n_2534),
.B(n_2464),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2610),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2560),
.B(n_2487),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_R g2807 ( 
.A(n_2580),
.B(n_2460),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2564),
.B(n_2490),
.Y(n_2808)
);

XNOR2xp5_ASAP7_75t_L g2809 ( 
.A(n_2558),
.B(n_2415),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2577),
.B(n_2465),
.Y(n_2810)
);

INVxp67_ASAP7_75t_L g2811 ( 
.A(n_2610),
.Y(n_2811)
);

XNOR2xp5_ASAP7_75t_L g2812 ( 
.A(n_2558),
.B(n_2342),
.Y(n_2812)
);

NAND2xp33_ASAP7_75t_R g2813 ( 
.A(n_2625),
.B(n_2447),
.Y(n_2813)
);

INVxp67_ASAP7_75t_L g2814 ( 
.A(n_2574),
.Y(n_2814)
);

INVxp67_ASAP7_75t_L g2815 ( 
.A(n_2574),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2790),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2765),
.B(n_2541),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2729),
.B(n_2545),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2696),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2667),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2773),
.Y(n_2821)
);

AOI22xp33_ASAP7_75t_L g2822 ( 
.A1(n_2701),
.A2(n_2652),
.B1(n_2649),
.B2(n_2619),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2682),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2737),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2697),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2713),
.B(n_2545),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2705),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2770),
.B(n_2581),
.Y(n_2828)
);

AOI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2772),
.A2(n_2618),
.B1(n_2626),
.B2(n_2657),
.Y(n_2829)
);

BUFx6f_ASAP7_75t_L g2830 ( 
.A(n_2761),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2700),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2774),
.B(n_2777),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2790),
.B(n_2562),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2702),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2726),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2776),
.B(n_2562),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2785),
.B(n_2581),
.Y(n_2837)
);

INVx1_ASAP7_75t_SL g2838 ( 
.A(n_2707),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2721),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2812),
.A2(n_2626),
.B1(n_2615),
.B2(n_2469),
.Y(n_2840)
);

AND2x4_ASAP7_75t_L g2841 ( 
.A(n_2776),
.B(n_2563),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2745),
.Y(n_2842)
);

AND2x4_ASAP7_75t_L g2843 ( 
.A(n_2783),
.B(n_2563),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2747),
.B(n_2536),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2806),
.B(n_2542),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2668),
.B(n_2567),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2732),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_L g2848 ( 
.A1(n_2809),
.A2(n_2605),
.B1(n_2606),
.B2(n_2583),
.Y(n_2848)
);

INVx4_ASAP7_75t_L g2849 ( 
.A(n_2731),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2741),
.B(n_2569),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2782),
.B(n_2603),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2698),
.B(n_2603),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2708),
.B(n_2565),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2693),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2803),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2793),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2801),
.B(n_2565),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2799),
.B(n_2570),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_2731),
.Y(n_2859)
);

INVxp67_ASAP7_75t_SL g2860 ( 
.A(n_2787),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2762),
.A2(n_2800),
.B1(n_2733),
.B2(n_2731),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2679),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2759),
.B(n_2612),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2727),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2744),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2727),
.Y(n_2866)
);

INVxp67_ASAP7_75t_SL g2867 ( 
.A(n_2802),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2771),
.Y(n_2868)
);

HB1xp67_ASAP7_75t_L g2869 ( 
.A(n_2692),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2681),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2730),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2753),
.B(n_2568),
.Y(n_2872)
);

OAI221xp5_ASAP7_75t_SL g2873 ( 
.A1(n_2766),
.A2(n_2583),
.B1(n_2616),
.B2(n_2627),
.C(n_2379),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2730),
.Y(n_2874)
);

AOI22xp33_ASAP7_75t_SL g2875 ( 
.A1(n_2794),
.A2(n_2568),
.B1(n_2543),
.B2(n_2544),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2750),
.Y(n_2876)
);

NOR3xp33_ASAP7_75t_L g2877 ( 
.A(n_2808),
.B(n_2506),
.C(n_2342),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2699),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2753),
.B(n_2631),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2754),
.B(n_2632),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2780),
.Y(n_2881)
);

NAND2x1p5_ASAP7_75t_L g2882 ( 
.A(n_2798),
.B(n_2660),
.Y(n_2882)
);

OAI21xp33_ASAP7_75t_L g2883 ( 
.A1(n_2807),
.A2(n_2627),
.B(n_2616),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2671),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2757),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2768),
.Y(n_2886)
);

INVx4_ASAP7_75t_L g2887 ( 
.A(n_2768),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2788),
.Y(n_2888)
);

OAI221xp5_ASAP7_75t_SL g2889 ( 
.A1(n_2784),
.A2(n_2392),
.B1(n_2557),
.B2(n_2553),
.C(n_2550),
.Y(n_2889)
);

INVxp67_ASAP7_75t_SL g2890 ( 
.A(n_2792),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2805),
.B(n_2571),
.Y(n_2891)
);

HB1xp67_ASAP7_75t_L g2892 ( 
.A(n_2778),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2680),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2659),
.Y(n_2894)
);

OAI21x1_ASAP7_75t_L g2895 ( 
.A1(n_2882),
.A2(n_2647),
.B(n_2740),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2885),
.B(n_2634),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2885),
.B(n_2642),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2827),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2865),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2820),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2824),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2817),
.B(n_2673),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2833),
.B(n_2763),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2821),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2817),
.B(n_2578),
.Y(n_2905)
);

NAND4xp25_ASAP7_75t_L g2906 ( 
.A(n_2873),
.B(n_2666),
.C(n_2678),
.D(n_2717),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2825),
.Y(n_2907)
);

INVx1_ASAP7_75t_SL g2908 ( 
.A(n_2868),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2851),
.B(n_2673),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2849),
.B(n_2720),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2888),
.B(n_2828),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2831),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2833),
.Y(n_2913)
);

BUFx4f_ASAP7_75t_SL g2914 ( 
.A(n_2865),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2851),
.B(n_2675),
.Y(n_2915)
);

NAND3xp33_ASAP7_75t_L g2916 ( 
.A(n_2883),
.B(n_2711),
.C(n_2677),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2832),
.B(n_2749),
.Y(n_2917)
);

OAI31xp33_ASAP7_75t_L g2918 ( 
.A1(n_2889),
.A2(n_2710),
.A3(n_2769),
.B(n_2738),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2832),
.B(n_2852),
.Y(n_2919)
);

OR2x2_ASAP7_75t_L g2920 ( 
.A(n_2888),
.B(n_2758),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2852),
.B(n_2675),
.Y(n_2921)
);

OAI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2877),
.A2(n_2689),
.B(n_2706),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2822),
.A2(n_2715),
.B1(n_2804),
.B2(n_2781),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2834),
.Y(n_2924)
);

AOI22xp5_ASAP7_75t_L g2925 ( 
.A1(n_2848),
.A2(n_2813),
.B1(n_2704),
.B2(n_2714),
.Y(n_2925)
);

OR2x6_ASAP7_75t_L g2926 ( 
.A(n_2849),
.B(n_2694),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2835),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2860),
.Y(n_2928)
);

BUFx3_ASAP7_75t_L g2929 ( 
.A(n_2886),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2886),
.Y(n_2930)
);

AO21x2_ASAP7_75t_L g2931 ( 
.A1(n_2891),
.A2(n_2746),
.B(n_2604),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2816),
.B(n_2686),
.Y(n_2932)
);

AND2x4_ASAP7_75t_L g2933 ( 
.A(n_2833),
.B(n_2763),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2839),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2847),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2823),
.Y(n_2936)
);

BUFx3_ASAP7_75t_L g2937 ( 
.A(n_2887),
.Y(n_2937)
);

HB1xp67_ASAP7_75t_L g2938 ( 
.A(n_2867),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2838),
.A2(n_2743),
.B1(n_2684),
.B2(n_2664),
.Y(n_2939)
);

AND2x4_ASAP7_75t_SL g2940 ( 
.A(n_2887),
.B(n_2761),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2842),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2856),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2887),
.Y(n_2943)
);

OR2x2_ASAP7_75t_L g2944 ( 
.A(n_2876),
.B(n_2764),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2816),
.B(n_2688),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2816),
.B(n_2864),
.Y(n_2946)
);

AOI221xp5_ASAP7_75t_L g2947 ( 
.A1(n_2829),
.A2(n_2815),
.B1(n_2814),
.B2(n_2811),
.C(n_2669),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2842),
.Y(n_2948)
);

OR2x2_ASAP7_75t_L g2949 ( 
.A(n_2876),
.B(n_2540),
.Y(n_2949)
);

INVx3_ASAP7_75t_L g2950 ( 
.A(n_2849),
.Y(n_2950)
);

AND2x4_ASAP7_75t_L g2951 ( 
.A(n_2843),
.B(n_2767),
.Y(n_2951)
);

CKINVDCx20_ASAP7_75t_R g2952 ( 
.A(n_2861),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2826),
.B(n_2540),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2855),
.Y(n_2954)
);

OAI33xp33_ASAP7_75t_L g2955 ( 
.A1(n_2878),
.A2(n_2734),
.A3(n_2760),
.B1(n_2665),
.B2(n_2703),
.B3(n_2797),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2855),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2819),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2928),
.B(n_2828),
.Y(n_2958)
);

AND2x2_ASAP7_75t_SL g2959 ( 
.A(n_2951),
.B(n_2843),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2904),
.Y(n_2960)
);

HB1xp67_ASAP7_75t_L g2961 ( 
.A(n_2928),
.Y(n_2961)
);

AND2x2_ASAP7_75t_L g2962 ( 
.A(n_2919),
.B(n_2837),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2938),
.Y(n_2963)
);

AND2x4_ASAP7_75t_L g2964 ( 
.A(n_2916),
.B(n_2843),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2909),
.B(n_2837),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2938),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2915),
.B(n_2871),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2914),
.B(n_2875),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2911),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2911),
.B(n_2826),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2898),
.B(n_2818),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2900),
.Y(n_2972)
);

HB1xp67_ASAP7_75t_L g2973 ( 
.A(n_2908),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2923),
.B(n_2884),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2902),
.B(n_2818),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2901),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2907),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2912),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2924),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2927),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2905),
.B(n_2869),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2935),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2936),
.Y(n_2983)
);

OR2x2_ASAP7_75t_L g2984 ( 
.A(n_2953),
.B(n_2949),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2942),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2952),
.B(n_2892),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2946),
.B(n_2853),
.Y(n_2987)
);

NAND2x1_ASAP7_75t_L g2988 ( 
.A(n_2926),
.B(n_2859),
.Y(n_2988)
);

BUFx2_ASAP7_75t_L g2989 ( 
.A(n_2914),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2957),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2921),
.B(n_2871),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2899),
.B(n_2882),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2954),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2899),
.Y(n_2994)
);

AOI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2918),
.A2(n_2859),
.B(n_2736),
.Y(n_2995)
);

OR2x2_ASAP7_75t_L g2996 ( 
.A(n_2917),
.B(n_2881),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2956),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2908),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2925),
.B(n_2893),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2904),
.Y(n_3000)
);

NAND2x1p5_ASAP7_75t_L g3001 ( 
.A(n_2937),
.B(n_2859),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2920),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2932),
.B(n_2853),
.Y(n_3003)
);

AND2x4_ASAP7_75t_L g3004 ( 
.A(n_2931),
.B(n_2836),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2934),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2896),
.Y(n_3006)
);

AND2x2_ASAP7_75t_SL g3007 ( 
.A(n_2951),
.B(n_2836),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2945),
.B(n_2857),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2896),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2897),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2913),
.B(n_2874),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2897),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2941),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2948),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2963),
.B(n_2840),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2966),
.B(n_2890),
.Y(n_3016)
);

NOR2x1_ASAP7_75t_L g3017 ( 
.A(n_2989),
.B(n_2906),
.Y(n_3017)
);

OAI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2995),
.A2(n_2906),
.B1(n_2926),
.B2(n_2952),
.Y(n_3018)
);

NOR4xp25_ASAP7_75t_SL g3019 ( 
.A(n_2968),
.B(n_2695),
.C(n_2676),
.D(n_2722),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_3006),
.B(n_2947),
.Y(n_3020)
);

AO221x2_ASAP7_75t_L g3021 ( 
.A1(n_3007),
.A2(n_2939),
.B1(n_2922),
.B2(n_2672),
.C(n_2662),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_3007),
.B(n_2913),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_R g3023 ( 
.A(n_2994),
.B(n_2691),
.Y(n_3023)
);

INVxp33_ASAP7_75t_SL g3024 ( 
.A(n_2986),
.Y(n_3024)
);

AO221x2_ASAP7_75t_L g3025 ( 
.A1(n_2959),
.A2(n_2922),
.B1(n_2955),
.B2(n_2894),
.C(n_2661),
.Y(n_3025)
);

AO221x2_ASAP7_75t_L g3026 ( 
.A1(n_2959),
.A2(n_2955),
.B1(n_2685),
.B2(n_2670),
.C(n_2926),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2958),
.B(n_2944),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_3009),
.B(n_2947),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2968),
.A2(n_2844),
.B1(n_2845),
.B2(n_2724),
.Y(n_3029)
);

INVx2_ASAP7_75t_SL g3030 ( 
.A(n_2994),
.Y(n_3030)
);

BUFx2_ASAP7_75t_L g3031 ( 
.A(n_2973),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_3010),
.B(n_2845),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_2998),
.Y(n_3033)
);

INVxp67_ASAP7_75t_L g3034 ( 
.A(n_2973),
.Y(n_3034)
);

AOI21xp33_ASAP7_75t_L g3035 ( 
.A1(n_2974),
.A2(n_2918),
.B(n_2674),
.Y(n_3035)
);

AO221x2_ASAP7_75t_L g3036 ( 
.A1(n_2988),
.A2(n_2735),
.B1(n_2719),
.B2(n_2866),
.C(n_2718),
.Y(n_3036)
);

NAND2xp33_ASAP7_75t_R g3037 ( 
.A(n_3004),
.B(n_2690),
.Y(n_3037)
);

INVxp67_ASAP7_75t_SL g3038 ( 
.A(n_2961),
.Y(n_3038)
);

NOR4xp25_ASAP7_75t_SL g3039 ( 
.A(n_2992),
.B(n_2687),
.C(n_2739),
.D(n_2728),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_3012),
.B(n_2862),
.Y(n_3040)
);

NAND2xp33_ASAP7_75t_SL g3041 ( 
.A(n_3004),
.B(n_2930),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2969),
.B(n_2854),
.Y(n_3042)
);

NOR4xp25_ASAP7_75t_SL g3043 ( 
.A(n_2992),
.B(n_2748),
.C(n_2716),
.D(n_2751),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2986),
.A2(n_2844),
.B1(n_2874),
.B2(n_2863),
.Y(n_3044)
);

NOR2x1_ASAP7_75t_L g3045 ( 
.A(n_3004),
.B(n_2937),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2999),
.B(n_2863),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2970),
.B(n_2870),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2996),
.B(n_2929),
.Y(n_3048)
);

INVx3_ASAP7_75t_L g3049 ( 
.A(n_3001),
.Y(n_3049)
);

NAND2xp33_ASAP7_75t_SL g3050 ( 
.A(n_2961),
.B(n_2950),
.Y(n_3050)
);

AO221x2_ASAP7_75t_L g3051 ( 
.A1(n_3001),
.A2(n_2943),
.B1(n_2933),
.B2(n_2903),
.C(n_2929),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_3038),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_3051),
.B(n_2964),
.Y(n_3053)
);

OR2x2_ASAP7_75t_L g3054 ( 
.A(n_3051),
.B(n_2984),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_3017),
.B(n_2964),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_3031),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_3020),
.B(n_2972),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_3040),
.Y(n_3058)
);

INVx1_ASAP7_75t_SL g3059 ( 
.A(n_3033),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3042),
.Y(n_3060)
);

INVx2_ASAP7_75t_SL g3061 ( 
.A(n_3023),
.Y(n_3061)
);

BUFx3_ASAP7_75t_L g3062 ( 
.A(n_3030),
.Y(n_3062)
);

NOR2xp33_ASAP7_75t_R g3063 ( 
.A(n_3037),
.B(n_2658),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3034),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_3024),
.B(n_2976),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_3016),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_3036),
.A2(n_2931),
.B(n_2964),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_3041),
.B(n_2943),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_3018),
.B(n_2977),
.Y(n_3069)
);

NAND3xp33_ASAP7_75t_L g3070 ( 
.A(n_3035),
.B(n_2755),
.C(n_2978),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3047),
.Y(n_3071)
);

INVx1_ASAP7_75t_SL g3072 ( 
.A(n_3050),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_3028),
.B(n_2979),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_3021),
.B(n_2965),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_3032),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_3021),
.B(n_2970),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_3027),
.Y(n_3077)
);

AO21x2_ASAP7_75t_L g3078 ( 
.A1(n_3029),
.A2(n_2390),
.B(n_2895),
.Y(n_3078)
);

AND2x4_ASAP7_75t_L g3079 ( 
.A(n_3045),
.B(n_2903),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_3015),
.B(n_2981),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_3036),
.B(n_3022),
.Y(n_3081)
);

BUFx2_ASAP7_75t_L g3082 ( 
.A(n_3049),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_3026),
.B(n_3019),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_3026),
.B(n_2962),
.Y(n_3084)
);

OAI21xp33_ASAP7_75t_L g3085 ( 
.A1(n_3044),
.A2(n_3002),
.B(n_2982),
.Y(n_3085)
);

INVx1_ASAP7_75t_SL g3086 ( 
.A(n_3048),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_3046),
.B(n_2933),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_3039),
.B(n_3008),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3025),
.Y(n_3089)
);

AOI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_3069),
.A2(n_3025),
.B1(n_2983),
.B2(n_2985),
.Y(n_3090)
);

INVxp67_ASAP7_75t_SL g3091 ( 
.A(n_3062),
.Y(n_3091)
);

OA21x2_ASAP7_75t_L g3092 ( 
.A1(n_3089),
.A2(n_3000),
.B(n_2960),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3052),
.Y(n_3093)
);

AND2x4_ASAP7_75t_SL g3094 ( 
.A(n_3061),
.B(n_2663),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_3059),
.B(n_2980),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_SL g3096 ( 
.A1(n_3072),
.A2(n_2742),
.B1(n_2910),
.B2(n_2950),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_3076),
.A2(n_2880),
.B1(n_2872),
.B2(n_2879),
.Y(n_3097)
);

OAI221xp5_ASAP7_75t_L g3098 ( 
.A1(n_3067),
.A2(n_2910),
.B1(n_2990),
.B2(n_2846),
.C(n_2712),
.Y(n_3098)
);

INVxp67_ASAP7_75t_L g3099 ( 
.A(n_3059),
.Y(n_3099)
);

NAND2xp33_ASAP7_75t_R g3100 ( 
.A(n_3063),
.B(n_3043),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3077),
.Y(n_3101)
);

AOI322xp5_ASAP7_75t_L g3102 ( 
.A1(n_3081),
.A2(n_3008),
.A3(n_3003),
.B1(n_2987),
.B2(n_2971),
.C1(n_2975),
.C2(n_3011),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3064),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_3086),
.B(n_2971),
.Y(n_3104)
);

AOI32xp33_ASAP7_75t_L g3105 ( 
.A1(n_3083),
.A2(n_2940),
.A3(n_3003),
.B1(n_2975),
.B2(n_2756),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_3079),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_3056),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_3082),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3075),
.B(n_2987),
.Y(n_3109)
);

AOI221xp5_ASAP7_75t_L g3110 ( 
.A1(n_3069),
.A2(n_2993),
.B1(n_2997),
.B2(n_3014),
.C(n_2858),
.Y(n_3110)
);

AOI21xp33_ASAP7_75t_SL g3111 ( 
.A1(n_3070),
.A2(n_2683),
.B(n_2709),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_3066),
.Y(n_3112)
);

OR2x2_ASAP7_75t_L g3113 ( 
.A(n_3057),
.B(n_3013),
.Y(n_3113)
);

AOI222xp33_ASAP7_75t_L g3114 ( 
.A1(n_3072),
.A2(n_2850),
.B1(n_3000),
.B2(n_2960),
.C1(n_3013),
.C2(n_3005),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_3080),
.B(n_2967),
.Y(n_3115)
);

INVxp67_ASAP7_75t_L g3116 ( 
.A(n_3065),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3091),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_3099),
.B(n_3058),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_3116),
.B(n_3060),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_3108),
.B(n_3057),
.Y(n_3120)
);

INVx1_ASAP7_75t_SL g3121 ( 
.A(n_3094),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3106),
.B(n_3053),
.Y(n_3122)
);

INVx1_ASAP7_75t_SL g3123 ( 
.A(n_3107),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_3106),
.B(n_3074),
.Y(n_3124)
);

INVx1_ASAP7_75t_SL g3125 ( 
.A(n_3103),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3104),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3110),
.B(n_3073),
.Y(n_3127)
);

INVx1_ASAP7_75t_SL g3128 ( 
.A(n_3093),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_3095),
.B(n_3086),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3109),
.Y(n_3130)
);

INVxp67_ASAP7_75t_L g3131 ( 
.A(n_3112),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_3092),
.Y(n_3132)
);

INVxp67_ASAP7_75t_L g3133 ( 
.A(n_3101),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_3102),
.B(n_3073),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3115),
.B(n_3071),
.Y(n_3135)
);

NAND2x1_ASAP7_75t_L g3136 ( 
.A(n_3092),
.B(n_3055),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_3114),
.B(n_3065),
.Y(n_3137)
);

CKINVDCx5p33_ASAP7_75t_R g3138 ( 
.A(n_3117),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_3121),
.B(n_3137),
.Y(n_3139)
);

HB1xp67_ASAP7_75t_L g3140 ( 
.A(n_3118),
.Y(n_3140)
);

CKINVDCx20_ASAP7_75t_R g3141 ( 
.A(n_3129),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3132),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_3132),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_3123),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3120),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3126),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3119),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3122),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3124),
.Y(n_3149)
);

INVx1_ASAP7_75t_SL g3150 ( 
.A(n_3125),
.Y(n_3150)
);

INVxp33_ASAP7_75t_L g3151 ( 
.A(n_3136),
.Y(n_3151)
);

INVx8_ASAP7_75t_L g3152 ( 
.A(n_3128),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3135),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3133),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3133),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3130),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_3142),
.B(n_3055),
.Y(n_3157)
);

NAND5xp2_ASAP7_75t_L g3158 ( 
.A(n_3139),
.B(n_3134),
.C(n_3105),
.D(n_3090),
.E(n_3067),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_3151),
.A2(n_3131),
.B(n_3127),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_3141),
.B(n_3096),
.Y(n_3160)
);

NOR4xp25_ASAP7_75t_L g3161 ( 
.A(n_3150),
.B(n_3131),
.C(n_3098),
.D(n_3088),
.Y(n_3161)
);

NAND3xp33_ASAP7_75t_L g3162 ( 
.A(n_3138),
.B(n_3100),
.C(n_3111),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3150),
.B(n_3085),
.Y(n_3163)
);

NOR2xp33_ASAP7_75t_SL g3164 ( 
.A(n_3144),
.B(n_3054),
.Y(n_3164)
);

NOR2x1_ASAP7_75t_L g3165 ( 
.A(n_3143),
.B(n_3084),
.Y(n_3165)
);

NAND3xp33_ASAP7_75t_SL g3166 ( 
.A(n_3154),
.B(n_3097),
.C(n_3068),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_3148),
.B(n_3079),
.Y(n_3167)
);

NAND4xp25_ASAP7_75t_L g3168 ( 
.A(n_3149),
.B(n_3113),
.C(n_2447),
.D(n_2410),
.Y(n_3168)
);

NAND3xp33_ASAP7_75t_SL g3169 ( 
.A(n_3155),
.B(n_2789),
.C(n_2786),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_3164),
.B(n_3152),
.Y(n_3170)
);

OAI211xp5_ASAP7_75t_L g3171 ( 
.A1(n_3162),
.A2(n_3159),
.B(n_3152),
.C(n_3160),
.Y(n_3171)
);

AOI222xp33_ASAP7_75t_L g3172 ( 
.A1(n_3163),
.A2(n_3145),
.B1(n_3152),
.B2(n_3153),
.C1(n_3147),
.C2(n_3146),
.Y(n_3172)
);

NOR4xp25_ASAP7_75t_L g3173 ( 
.A(n_3166),
.B(n_3156),
.C(n_3140),
.D(n_2298),
.Y(n_3173)
);

NAND3xp33_ASAP7_75t_SL g3174 ( 
.A(n_3161),
.B(n_3167),
.C(n_3158),
.Y(n_3174)
);

NOR3xp33_ASAP7_75t_L g3175 ( 
.A(n_3169),
.B(n_2333),
.C(n_2404),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_L g3176 ( 
.A1(n_3165),
.A2(n_3078),
.B1(n_3087),
.B2(n_2725),
.Y(n_3176)
);

AND3x1_ASAP7_75t_L g3177 ( 
.A(n_3157),
.B(n_3078),
.C(n_2506),
.Y(n_3177)
);

O2A1O1Ixp33_ASAP7_75t_L g3178 ( 
.A1(n_3168),
.A2(n_2458),
.B(n_2384),
.C(n_3087),
.Y(n_3178)
);

OAI211xp5_ASAP7_75t_SL g3179 ( 
.A1(n_3160),
.A2(n_2404),
.B(n_2328),
.C(n_2295),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_3170),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_3171),
.B(n_2723),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_3177),
.Y(n_3182)
);

NAND4xp75_ASAP7_75t_L g3183 ( 
.A(n_3172),
.B(n_2328),
.C(n_2810),
.D(n_2481),
.Y(n_3183)
);

AO22x1_ASAP7_75t_L g3184 ( 
.A1(n_3175),
.A2(n_2725),
.B1(n_2321),
.B2(n_2303),
.Y(n_3184)
);

XNOR2xp5_ASAP7_75t_L g3185 ( 
.A(n_3183),
.B(n_3174),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3184),
.B(n_3173),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_SL g3187 ( 
.A(n_3180),
.B(n_3176),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_R g3188 ( 
.A(n_3181),
.B(n_3179),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3182),
.B(n_3178),
.Y(n_3189)
);

AOI21xp33_ASAP7_75t_L g3190 ( 
.A1(n_3185),
.A2(n_2709),
.B(n_2321),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3187),
.B(n_3188),
.Y(n_3191)
);

OAI22x1_ASAP7_75t_L g3192 ( 
.A1(n_3186),
.A2(n_2320),
.B1(n_2365),
.B2(n_2694),
.Y(n_3192)
);

INVxp67_ASAP7_75t_L g3193 ( 
.A(n_3189),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3191),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3193),
.B(n_2940),
.Y(n_3195)
);

NAND2x1p5_ASAP7_75t_L g3196 ( 
.A(n_3194),
.B(n_3190),
.Y(n_3196)
);

AOI31xp33_ASAP7_75t_L g3197 ( 
.A1(n_3196),
.A2(n_3195),
.A3(n_3192),
.B(n_2365),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3196),
.A2(n_2830),
.B1(n_2779),
.B2(n_2991),
.Y(n_3198)
);

XOR2xp5_ASAP7_75t_L g3199 ( 
.A(n_3198),
.B(n_2830),
.Y(n_3199)
);

AOI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_3199),
.A2(n_3197),
.B1(n_2841),
.B2(n_2836),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3200),
.Y(n_3201)
);

OAI221xp5_ASAP7_75t_R g3202 ( 
.A1(n_3201),
.A2(n_2795),
.B1(n_2775),
.B2(n_2752),
.C(n_2796),
.Y(n_3202)
);

AOI211xp5_ASAP7_75t_L g3203 ( 
.A1(n_3202),
.A2(n_2325),
.B(n_2830),
.C(n_2791),
.Y(n_3203)
);


endmodule