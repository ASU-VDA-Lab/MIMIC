module fake_netlist_5_1628_n_1255 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1255);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1255;

wire n_924;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1182;
wire n_579;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_533;
wire n_1251;
wire n_278;

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_40),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_90),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_88),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_72),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_32),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_145),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_56),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_117),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_15),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_64),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_47),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_144),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_71),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_67),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_66),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_24),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_23),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_135),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_65),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_167),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_2),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_32),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_55),
.Y(n_229)
);

CKINVDCx6p67_ASAP7_75t_R g230 ( 
.A(n_60),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_83),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_0),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_82),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_152),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_81),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_181),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_189),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_191),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_192),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_202),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

CKINVDCx11_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_255),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_182),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_263),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_263),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_244),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_247),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_241),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_251),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_237),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_255),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_264),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_237),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_267),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_293),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_271),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_277),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_315),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_289),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_290),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_290),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_289),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_291),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_291),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_292),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_292),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_299),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_299),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_284),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_300),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_300),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_300),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_356),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_302),
.Y(n_375)
);

BUFx8_ASAP7_75t_SL g376 ( 
.A(n_318),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_300),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_307),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_298),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_203),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_203),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_302),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_223),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_343),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_223),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_335),
.B(n_199),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

BUFx8_ASAP7_75t_SL g396 ( 
.A(n_321),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_304),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_304),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_344),
.B(n_204),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

BUFx12f_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_312),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_312),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_390),
.A2(n_321),
.B1(n_362),
.B2(n_348),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_339),
.Y(n_417)
);

NAND2x1p5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_208),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_395),
.A2(n_377),
.B(n_381),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_390),
.A2(n_362),
.B1(n_352),
.B2(n_348),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_371),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_379),
.A2(n_386),
.B(n_385),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_380),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_400),
.A2(n_316),
.B1(n_340),
.B2(n_353),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_368),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_349),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_316),
.B1(n_226),
.B2(n_221),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_209),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_215),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_357),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_389),
.B(n_359),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_376),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_373),
.B(n_195),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_394),
.B(n_387),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_387),
.A2(n_399),
.B1(n_406),
.B2(n_405),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_392),
.A2(n_220),
.B(n_180),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_409),
.A2(n_352),
.B1(n_355),
.B2(n_350),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_373),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_396),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_231),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_399),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_373),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_196),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_403),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_408),
.B(n_323),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_405),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_182),
.Y(n_469)
);

AOI22x1_ASAP7_75t_SL g470 ( 
.A1(n_409),
.A2(n_226),
.B1(n_232),
.B2(n_198),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_406),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_406),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_393),
.B(n_210),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_382),
.B(n_285),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_411),
.B(n_232),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

AND3x2_ASAP7_75t_L g485 ( 
.A(n_407),
.B(n_184),
.C(n_206),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_222),
.Y(n_487)
);

OAI22x1_ASAP7_75t_SL g488 ( 
.A1(n_410),
.A2(n_224),
.B1(n_213),
.B2(n_186),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_401),
.A2(n_303),
.B(n_301),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_233),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_378),
.B(n_185),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

CKINVDCx6p67_ASAP7_75t_R g497 ( 
.A(n_410),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_398),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_388),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_443),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_443),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_456),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_456),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_464),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_464),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_414),
.A2(n_410),
.B1(n_216),
.B2(n_214),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_466),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_427),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_481),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_422),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_497),
.B(n_410),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_452),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_416),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_R g524 ( 
.A(n_497),
.B(n_438),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_466),
.B(n_378),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_428),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_487),
.B(n_372),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_440),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_487),
.B(n_463),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_440),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_436),
.B(n_388),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_436),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_413),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_438),
.B(n_391),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_465),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_465),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_431),
.B(n_391),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_R g548 ( 
.A(n_417),
.B(n_391),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_470),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_413),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_488),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_467),
.B(n_378),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_417),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_431),
.B(n_391),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_483),
.B(n_230),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_432),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_471),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_479),
.B(n_404),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_482),
.B(n_404),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_444),
.B(n_190),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_490),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_444),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_521),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_521),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_528),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_528),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_500),
.B(n_476),
.C(n_485),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_537),
.B(n_444),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_502),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_538),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_554),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_494),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_524),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_517),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

INVx8_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_540),
.B(n_478),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_560),
.B(n_453),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_545),
.B(n_538),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_550),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

AOI21x1_ASAP7_75t_L g591 ( 
.A1(n_531),
.A2(n_469),
.B(n_458),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_555),
.B(n_482),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_503),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_551),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_501),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_529),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_557),
.B(n_489),
.C(n_484),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_448),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_460),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_541),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_530),
.B(n_535),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_558),
.B(n_478),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_526),
.B(n_418),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_568),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_597),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_565),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_580),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_597),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_600),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_573),
.B(n_524),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_576),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_584),
.B(n_455),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_600),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_575),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_577),
.B(n_518),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_596),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_596),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_575),
.Y(n_627)
);

CKINVDCx6p67_ASAP7_75t_R g628 ( 
.A(n_576),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_572),
.B(n_579),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_572),
.B(n_512),
.C(n_559),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_586),
.B(n_592),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_601),
.B(n_561),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_601),
.B(n_592),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_570),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_590),
.B(n_544),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_598),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_581),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_578),
.Y(n_642)
);

INVxp67_ASAP7_75t_R g643 ( 
.A(n_580),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_602),
.B(n_544),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_598),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_596),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_582),
.B(n_506),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_578),
.B(n_566),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_599),
.B(n_520),
.C(n_606),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_606),
.B(n_532),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_596),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_571),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_603),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_578),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_587),
.B(n_532),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g658 ( 
.A(n_582),
.B(n_450),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_599),
.A2(n_519),
.B1(n_548),
.B2(n_184),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_585),
.B(n_548),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_574),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_605),
.B(n_493),
.C(n_492),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_581),
.B(n_516),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_584),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_583),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_505),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_584),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_593),
.A2(n_491),
.B1(n_523),
.B2(n_522),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_595),
.B(n_477),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_594),
.B(n_496),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_595),
.B(n_571),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_583),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_584),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_569),
.B(n_498),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_583),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_591),
.B(n_499),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_591),
.B(n_478),
.C(n_553),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_584),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_455),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_577),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_584),
.B(n_518),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_573),
.B(n_467),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_596),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_573),
.B(n_467),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

AND3x2_ASAP7_75t_L g689 ( 
.A(n_586),
.B(n_459),
.C(n_457),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_667),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_650),
.B(n_478),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_639),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_631),
.B(n_644),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_608),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_613),
.B(n_513),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_611),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_629),
.A2(n_680),
.B(n_659),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_418),
.Y(n_698)
);

XOR2xp5_ASAP7_75t_L g699 ( 
.A(n_648),
.B(n_507),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_612),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_636),
.B(n_491),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_613),
.B(n_513),
.Y(n_702)
);

XOR2xp5_ASAP7_75t_L g703 ( 
.A(n_610),
.B(n_508),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_617),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_632),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_634),
.Y(n_707)
);

BUFx6f_ASAP7_75t_SL g708 ( 
.A(n_618),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_509),
.Y(n_709)
);

XNOR2xp5_ASAP7_75t_L g710 ( 
.A(n_614),
.B(n_510),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_638),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_688),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_618),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g714 ( 
.A(n_614),
.B(n_511),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_629),
.B(n_491),
.Y(n_715)
);

AND2x2_ASAP7_75t_SL g716 ( 
.A(n_684),
.B(n_501),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_651),
.B(n_190),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_616),
.B(n_457),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_684),
.A2(n_556),
.B(n_527),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_677),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_659),
.A2(n_437),
.B(n_434),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_677),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_609),
.B(n_639),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_673),
.Y(n_724)
);

CKINVDCx16_ASAP7_75t_R g725 ( 
.A(n_620),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_657),
.B(n_515),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_657),
.B(n_549),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_640),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_652),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_645),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_620),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_653),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_621),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_655),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_661),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_666),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_678),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_683),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_672),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_619),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_619),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_615),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_633),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_627),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_627),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_635),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_635),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_658),
.B(n_230),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_652),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_607),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_642),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_642),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_623),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_656),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_656),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_685),
.A2(n_556),
.B(n_527),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_641),
.Y(n_758)
);

INVxp33_ASAP7_75t_L g759 ( 
.A(n_660),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_658),
.B(n_183),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_665),
.B(n_491),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_665),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_624),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_674),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_674),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_630),
.B(n_183),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_637),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_654),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_685),
.B(n_491),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_687),
.B(n_442),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_660),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_670),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_687),
.B(n_442),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_679),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_774),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_694),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_740),
.B(n_720),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_693),
.B(n_643),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_690),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_696),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_723),
.B(n_630),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_692),
.B(n_186),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_758),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_772),
.B(n_671),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_671),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_744),
.B(n_649),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_725),
.B(n_681),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_732),
.B(n_649),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_726),
.B(n_212),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_700),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_749),
.A2(n_682),
.B1(n_616),
.B2(n_668),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_704),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_709),
.B(n_212),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_705),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_766),
.A2(n_682),
.B1(n_616),
.B2(n_668),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_713),
.B(n_662),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_710),
.B(n_662),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_729),
.B(n_649),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_706),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_760),
.A2(n_504),
.B1(n_682),
.B2(n_207),
.Y(n_800)
);

NAND2x1p5_ASAP7_75t_L g801 ( 
.A(n_716),
.B(n_626),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_707),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_698),
.B(n_622),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_714),
.B(n_504),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_711),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_771),
.A2(n_504),
.B1(n_207),
.B2(n_664),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_712),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_731),
.B(n_649),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_733),
.B(n_649),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_735),
.B(n_689),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_736),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_737),
.B(n_689),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_759),
.B(n_622),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_741),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_767),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_697),
.B(n_664),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_717),
.B(n_675),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_739),
.B(n_214),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_743),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_745),
.B(n_646),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_697),
.A2(n_669),
.B(n_233),
.C(n_234),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_691),
.A2(n_727),
.B1(n_708),
.B2(n_728),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_715),
.B(n_652),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_708),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_701),
.A2(n_504),
.B1(n_207),
.B2(n_179),
.Y(n_829)
);

NOR2x1p5_ASAP7_75t_L g830 ( 
.A(n_701),
.B(n_675),
.Y(n_830)
);

AOI221xp5_ASAP7_75t_L g831 ( 
.A1(n_715),
.A2(n_234),
.B1(n_216),
.B2(n_185),
.C(n_187),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_768),
.B(n_646),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_721),
.A2(n_504),
.B1(n_185),
.B2(n_187),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_751),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_746),
.B(n_647),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_699),
.B(n_703),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_718),
.B(n_652),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_695),
.B(n_229),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_754),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_695),
.B(n_702),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_235),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_763),
.B(n_676),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_730),
.B(n_750),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_769),
.B(n_773),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_730),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_730),
.B(n_236),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_747),
.B(n_647),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_750),
.Y(n_848)
);

NAND2x1_ASAP7_75t_L g849 ( 
.A(n_718),
.B(n_686),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_775),
.B(n_718),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_820),
.B(n_750),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_826),
.A2(n_669),
.B1(n_719),
.B2(n_769),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_825),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_SL g854 ( 
.A(n_795),
.B(n_801),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_791),
.B(n_719),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_779),
.B(n_770),
.Y(n_856)
);

OAI22xp33_ASAP7_75t_L g857 ( 
.A1(n_800),
.A2(n_773),
.B1(n_770),
.B2(n_757),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_793),
.B(n_761),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_789),
.B(n_761),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_777),
.B(n_748),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_801),
.B(n_757),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_780),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_776),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_794),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_781),
.B(n_686),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_802),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_797),
.A2(n_721),
.B(n_764),
.C(n_762),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_783),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_837),
.B(n_752),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_778),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_828),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_790),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_796),
.B(n_187),
.C(n_753),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_804),
.A2(n_786),
.B1(n_788),
.B2(n_782),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_792),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_822),
.B(n_0),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_819),
.A2(n_756),
.B(n_755),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_844),
.B(n_686),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_777),
.B(n_765),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_830),
.A2(n_187),
.B1(n_563),
.B2(n_562),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_799),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_840),
.B(n_1),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_805),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_836),
.B(n_3),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_807),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_817),
.B(n_686),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_784),
.B(n_626),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_808),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_809),
.B(n_3),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_816),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_838),
.B(n_841),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_785),
.B(n_626),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_821),
.B(n_4),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_834),
.B(n_4),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_848),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_839),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_846),
.B(n_803),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_787),
.A2(n_833),
.B1(n_806),
.B2(n_831),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_824),
.A2(n_495),
.B(n_513),
.C(n_547),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_812),
.B(n_626),
.Y(n_903)
);

AO22x1_ASAP7_75t_L g904 ( 
.A1(n_812),
.A2(n_424),
.B1(n_6),
.B2(n_7),
.Y(n_904)
);

OAI221xp5_ASAP7_75t_L g905 ( 
.A1(n_814),
.A2(n_462),
.B1(n_472),
.B2(n_468),
.C(n_461),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_814),
.B(n_501),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_823),
.B(n_835),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_847),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_823),
.B(n_5),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_847),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_845),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_837),
.B(n_451),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_810),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_832),
.B(n_5),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_798),
.B(n_7),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_848),
.B(n_501),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_849),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_811),
.B(n_8),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_829),
.A2(n_425),
.B(n_419),
.Y(n_919)
);

BUFx12f_ASAP7_75t_L g920 ( 
.A(n_837),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_810),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_842),
.B(n_525),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_827),
.B(n_8),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_827),
.B(n_9),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_843),
.B(n_9),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_827),
.B(n_10),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_827),
.A2(n_563),
.B1(n_562),
.B2(n_424),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_828),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_826),
.A2(n_547),
.B1(n_474),
.B2(n_473),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_825),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_861),
.B(n_855),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_853),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_854),
.B(n_525),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_871),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_873),
.A2(n_547),
.B1(n_525),
.B2(n_425),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_854),
.B(n_525),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_920),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_853),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_908),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_917),
.B(n_419),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_917),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_861),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_SL g944 ( 
.A(n_851),
.B(n_475),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_928),
.B(n_10),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_921),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_910),
.B(n_11),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_928),
.Y(n_948)
);

AND2x4_ASAP7_75t_SL g949 ( 
.A(n_868),
.B(n_445),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_872),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_881),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_L g952 ( 
.A(n_873),
.B(n_475),
.Y(n_952)
);

OR2x2_ASAP7_75t_SL g953 ( 
.A(n_909),
.B(n_425),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_913),
.B(n_11),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_892),
.B(n_12),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_885),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_850),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_911),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_870),
.B(n_12),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_930),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_850),
.B(n_13),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_916),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_907),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_862),
.B(n_14),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_889),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_SL g966 ( 
.A(n_896),
.B(n_14),
.C(n_15),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_895),
.B(n_16),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_894),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_916),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_900),
.B(n_884),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_875),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_883),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_888),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_891),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_898),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_864),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_899),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_869),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_860),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_867),
.B(n_475),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_879),
.B(n_16),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_869),
.B(n_17),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_874),
.B(n_858),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_856),
.B(n_17),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_886),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_948),
.B(n_943),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_956),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_934),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_948),
.B(n_915),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_932),
.Y(n_991)
);

AND3x1_ASAP7_75t_L g992 ( 
.A(n_966),
.B(n_876),
.C(n_925),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_938),
.B(n_918),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_978),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_942),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_986),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_934),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_958),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_934),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_963),
.B(n_865),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_956),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_979),
.B(n_857),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_939),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_958),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_933),
.B(n_924),
.C(n_923),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_962),
.B(n_861),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_985),
.B(n_903),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_931),
.B(n_906),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_972),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_958),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_983),
.B(n_882),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_982),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_937),
.B(n_914),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_953),
.B(n_893),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_931),
.B(n_887),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_R g1016 ( 
.A(n_960),
.B(n_926),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_941),
.B(n_877),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_950),
.B(n_922),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_SL g1019 ( 
.A(n_966),
.B(n_878),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_972),
.Y(n_1020)
);

BUFx4f_ASAP7_75t_L g1021 ( 
.A(n_982),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_936),
.A2(n_901),
.B1(n_880),
.B2(n_905),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_943),
.B(n_859),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_931),
.B(n_890),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_980),
.B(n_904),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_973),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_973),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_967),
.A2(n_929),
.B1(n_852),
.B2(n_927),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_951),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_965),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_943),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_968),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_955),
.A2(n_970),
.B1(n_945),
.B2(n_957),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_954),
.B(n_946),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_976),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_977),
.Y(n_1036)
);

AND2x4_ASAP7_75t_SL g1037 ( 
.A(n_961),
.B(n_912),
.Y(n_1037)
);

NOR2x1_ASAP7_75t_L g1038 ( 
.A(n_947),
.B(n_897),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_971),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_947),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_954),
.B(n_919),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_974),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_964),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_975),
.B(n_943),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_964),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_981),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_961),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_944),
.B(n_916),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_952),
.A2(n_912),
.B1(n_916),
.B2(n_447),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_981),
.B(n_902),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1040),
.B(n_1045),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1019),
.B(n_959),
.C(n_984),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_1012),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1011),
.A2(n_935),
.B1(n_940),
.B2(n_984),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_935),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1012),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1025),
.A2(n_940),
.B(n_949),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1029),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1025),
.A2(n_969),
.B(n_962),
.Y(n_1060)
);

AO32x1_ASAP7_75t_L g1061 ( 
.A1(n_1022),
.A2(n_969),
.A3(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1025),
.A2(n_992),
.B(n_1041),
.Y(n_1062)
);

BUFx4f_ASAP7_75t_L g1063 ( 
.A(n_989),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_1023),
.A2(n_495),
.B(n_454),
.C(n_445),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_991),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_997),
.B(n_424),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_994),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1030),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1043),
.B(n_18),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1036),
.B(n_18),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1065),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1062),
.B(n_1038),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1070),
.A2(n_1069),
.B(n_1060),
.Y(n_1073)
);

AND3x4_ASAP7_75t_L g1074 ( 
.A(n_1057),
.B(n_1004),
.C(n_1005),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_1070),
.A2(n_987),
.B(n_998),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1053),
.A2(n_996),
.B(n_994),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_1063),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_1052),
.A2(n_1051),
.B(n_1056),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1054),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_1053),
.B(n_989),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_1063),
.A2(n_1021),
.B(n_1033),
.C(n_1050),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1067),
.B(n_1044),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_1058),
.A2(n_996),
.B(n_988),
.Y(n_1083)
);

BUFx8_ASAP7_75t_L g1084 ( 
.A(n_1054),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1055),
.B(n_1002),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1054),
.B(n_991),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1059),
.Y(n_1087)
);

NAND2x1_ASAP7_75t_L g1088 ( 
.A(n_1068),
.B(n_1015),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_L g1089 ( 
.A(n_1061),
.B(n_1015),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1061),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1061),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1064),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_1066),
.B(n_997),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1059),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_1071),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1086),
.B(n_997),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1090),
.A2(n_1024),
.B1(n_1014),
.B2(n_1028),
.Y(n_1098)
);

OAI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1081),
.A2(n_992),
.B1(n_993),
.B2(n_1013),
.C(n_1021),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1090),
.A2(n_1006),
.B1(n_1024),
.B2(n_1008),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1084),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1084),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_1081),
.B(n_1078),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_SL g1104 ( 
.A(n_1102),
.B(n_999),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1104),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1103),
.A2(n_1099),
.B1(n_1078),
.B2(n_1072),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1105),
.Y(n_1107)
);

OAI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1106),
.A2(n_1089),
.B1(n_1072),
.B2(n_1091),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_1096),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_1101),
.B(n_1098),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1107),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1110),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1110),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1112),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1112),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1116),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1115),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1118),
.A2(n_1112),
.B1(n_1114),
.B2(n_1109),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1117),
.B(n_1097),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_1114),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_1113),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_1100),
.B1(n_1080),
.B2(n_1077),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1124),
.B(n_1080),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1126),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1125),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_1079),
.B1(n_1080),
.B2(n_1074),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1128),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1127),
.B(n_1079),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1129),
.B(n_1079),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1130),
.A2(n_1087),
.B1(n_1092),
.B2(n_1095),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1131),
.B(n_1073),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1134),
.B(n_1132),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1133),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1135),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1136),
.Y(n_1138)
);

OAI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_1137),
.A2(n_1085),
.B1(n_1010),
.B2(n_1075),
.C(n_1088),
.Y(n_1139)
);

AO221x2_ASAP7_75t_L g1140 ( 
.A1(n_1138),
.A2(n_1094),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1140),
.B(n_1082),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1141),
.B(n_1142),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1141),
.B(n_19),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1144),
.Y(n_1145)
);

OR2x2_ASAP7_75t_L g1146 ( 
.A(n_1143),
.B(n_22),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_23),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1147),
.Y(n_1148)
);

AOI222xp33_ASAP7_75t_L g1149 ( 
.A1(n_1145),
.A2(n_1094),
.B1(n_1093),
.B2(n_990),
.C1(n_27),
.C2(n_28),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1146),
.B(n_24),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1148),
.B(n_1076),
.Y(n_1151)
);

AOI221xp5_ASAP7_75t_L g1152 ( 
.A1(n_1150),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_1149),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1152),
.A2(n_280),
.B(n_301),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_25),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1154),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1155),
.A2(n_1156),
.B1(n_29),
.B2(n_30),
.Y(n_1157)
);

OAI221xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1155),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.C(n_33),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_1157),
.B(n_31),
.C(n_33),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1159),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1160),
.Y(n_1162)
);

OAI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1161),
.A2(n_1093),
.B1(n_1047),
.B2(n_1031),
.Y(n_1163)
);

AOI211x1_ASAP7_75t_SL g1164 ( 
.A1(n_1162),
.A2(n_280),
.B(n_1034),
.C(n_305),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1161),
.A2(n_995),
.B1(n_1031),
.B2(n_404),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1164),
.A2(n_305),
.B1(n_995),
.B2(n_36),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_SL g1167 ( 
.A(n_1165),
.B(n_280),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_1163),
.B(n_280),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_L g1169 ( 
.A1(n_1167),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1168),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1170),
.B(n_1166),
.Y(n_1171)
);

AOI211xp5_ASAP7_75t_L g1172 ( 
.A1(n_1169),
.A2(n_280),
.B(n_276),
.C(n_41),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1171),
.A2(n_276),
.B(n_39),
.C(n_42),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1172),
.B(n_38),
.Y(n_1174)
);

OAI211xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1174),
.A2(n_276),
.B(n_44),
.C(n_45),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1173),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1176),
.B(n_1083),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_1175),
.B(n_276),
.C(n_43),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1178),
.B(n_276),
.C(n_404),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1177),
.B(n_276),
.C(n_404),
.Y(n_1180)
);

XNOR2x1_ASAP7_75t_L g1181 ( 
.A(n_1179),
.B(n_46),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1180),
.B(n_276),
.C(n_48),
.Y(n_1182)
);

NAND5xp2_ASAP7_75t_L g1183 ( 
.A(n_1179),
.B(n_49),
.C(n_51),
.D(n_52),
.E(n_53),
.Y(n_1183)
);

NOR3x1_ASAP7_75t_L g1184 ( 
.A(n_1181),
.B(n_54),
.C(n_57),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1182),
.B(n_58),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1183),
.B(n_1031),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1186),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_1185),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1187),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1188),
.A2(n_1184),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_1190)
);

AND2x2_ASAP7_75t_SL g1191 ( 
.A(n_1189),
.B(n_59),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1190),
.B(n_68),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1192),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1191),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1193),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1194),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1195),
.Y(n_1197)
);

OAI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1196),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.C(n_77),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1197),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1198),
.A2(n_404),
.B1(n_79),
.B2(n_84),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_L g1201 ( 
.A(n_1197),
.B(n_78),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1199),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1200),
.A2(n_85),
.B(n_86),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1201),
.A2(n_87),
.B(n_89),
.Y(n_1204)
);

AOI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1202),
.A2(n_1203),
.B1(n_1204),
.B2(n_95),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1202),
.A2(n_1048),
.B1(n_446),
.B2(n_441),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1205),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1206),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1208),
.B(n_420),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1207),
.B(n_91),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1209),
.B(n_93),
.Y(n_1211)
);

OAI21xp33_ASAP7_75t_L g1212 ( 
.A1(n_1210),
.A2(n_1016),
.B(n_97),
.Y(n_1212)
);

AOI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1209),
.A2(n_96),
.B(n_98),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1211),
.Y(n_1214)
);

AOI21xp33_ASAP7_75t_L g1215 ( 
.A1(n_1213),
.A2(n_99),
.B(n_100),
.Y(n_1215)
);

AO22x1_ASAP7_75t_L g1216 ( 
.A1(n_1212),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1214),
.A2(n_1006),
.B1(n_446),
.B2(n_441),
.Y(n_1217)
);

AO22x1_ASAP7_75t_L g1218 ( 
.A1(n_1216),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1215),
.A2(n_446),
.B1(n_441),
.B2(n_420),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1219),
.B(n_107),
.Y(n_1220)
);

XNOR2xp5_ASAP7_75t_L g1221 ( 
.A(n_1218),
.B(n_109),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1217),
.A2(n_110),
.B(n_111),
.Y(n_1222)
);

OAI222xp33_ASAP7_75t_SL g1223 ( 
.A1(n_1219),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.C1(n_116),
.C2(n_118),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1219),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_1224)
);

OA21x2_ASAP7_75t_L g1225 ( 
.A1(n_1219),
.A2(n_123),
.B(n_124),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1219),
.A2(n_125),
.B(n_126),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1219),
.A2(n_420),
.B1(n_441),
.B2(n_446),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1219),
.A2(n_127),
.B(n_130),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1219),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1219),
.B(n_132),
.Y(n_1230)
);

OAI321xp33_ASAP7_75t_L g1231 ( 
.A1(n_1219),
.A2(n_136),
.A3(n_137),
.B1(n_139),
.B2(n_140),
.C(n_141),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_SL g1232 ( 
.A1(n_1219),
.A2(n_142),
.B(n_147),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1229),
.A2(n_149),
.B(n_151),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1221),
.A2(n_153),
.B(n_154),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_156),
.B(n_157),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1230),
.A2(n_158),
.B(n_159),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1220),
.B(n_160),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1222),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1225),
.B(n_162),
.Y(n_1239)
);

NAND2x1_ASAP7_75t_L g1240 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1231),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1241),
.A2(n_1228),
.B1(n_1226),
.B2(n_1223),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1238),
.A2(n_1224),
.B1(n_164),
.B2(n_165),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1240),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1239),
.A2(n_1037),
.B1(n_420),
.B2(n_168),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1235),
.A2(n_163),
.B1(n_166),
.B2(n_170),
.Y(n_1246)
);

AOI322xp5_ASAP7_75t_L g1247 ( 
.A1(n_1237),
.A2(n_171),
.A3(n_172),
.B1(n_173),
.B2(n_176),
.C1(n_1008),
.C2(n_1049),
.Y(n_1247)
);

OA22x2_ASAP7_75t_L g1248 ( 
.A1(n_1244),
.A2(n_1237),
.B1(n_1234),
.B2(n_1236),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1242),
.A2(n_1233),
.B1(n_1001),
.B2(n_1027),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1243),
.B(n_1246),
.Y(n_1250)
);

AOI221xp5_ASAP7_75t_L g1251 ( 
.A1(n_1248),
.A2(n_1245),
.B1(n_1247),
.B2(n_1020),
.C(n_1009),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1251),
.A2(n_1250),
.B1(n_1249),
.B2(n_1026),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1252),
.A2(n_1035),
.B1(n_1032),
.B2(n_1042),
.Y(n_1253)
);

AOI211xp5_ASAP7_75t_L g1254 ( 
.A1(n_1253),
.A2(n_1007),
.B(n_1000),
.C(n_1018),
.Y(n_1254)
);

AOI211xp5_ASAP7_75t_L g1255 ( 
.A1(n_1254),
.A2(n_1017),
.B(n_1039),
.C(n_1003),
.Y(n_1255)
);


endmodule