module real_jpeg_28579_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_287, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_287;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_167;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_18),
.B1(n_19),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_23),
.B(n_26),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_44),
.B1(n_72),
.B2(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_0),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_22),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_0),
.A2(n_50),
.B(n_55),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_0),
.A2(n_8),
.B(n_73),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_0),
.B(n_49),
.Y(n_173)
);

INVx11_ASAP7_75t_SL g74 ( 
.A(n_1),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_5),
.A2(n_33),
.B1(n_72),
.B2(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_5),
.A2(n_33),
.B1(n_50),
.B2(n_52),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_61),
.Y(n_119)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_17),
.B1(n_50),
.B2(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_17),
.B1(n_72),
.B2(n_73),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_36),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_29),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_18),
.A2(n_25),
.B(n_44),
.C(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_21),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_27),
.B1(n_43),
.B2(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_23),
.A2(n_24),
.B1(n_51),
.B2(n_55),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_23),
.A2(n_44),
.B(n_56),
.C(n_148),
.Y(n_147)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_30),
.B(n_38),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_76),
.B(n_285),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_39),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_39),
.B(n_283),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.CI(n_57),
.CON(n_39),
.SN(n_39)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_41),
.A2(n_42),
.B(n_60),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_43),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_44),
.A2(n_50),
.B(n_70),
.C(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_44),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_44),
.B(n_71),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_49),
.B1(n_53),
.B2(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_48),
.B(n_88),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_49),
.A2(n_63),
.B(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_89),
.Y(n_108)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_58),
.B(n_92),
.C(n_93),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_58),
.A2(n_91),
.B1(n_107),
.B2(n_132),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_58),
.B(n_132),
.C(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_58),
.A2(n_91),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_62),
.A2(n_64),
.B1(n_264),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_62),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_64),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_64),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_67),
.A2(n_71),
.B1(n_112),
.B2(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_67),
.A2(n_71),
.B1(n_75),
.B2(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_71),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_72),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_100),
.Y(n_99)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_282),
.B(n_284),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_256),
.A3(n_275),
.B1(n_280),
.B2(n_281),
.C(n_287),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_239),
.B(n_255),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_220),
.B(n_238),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_141),
.B(n_203),
.C(n_219),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_129),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_82),
.B(n_129),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_104),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_83),
.B(n_105),
.C(n_115),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_138),
.C(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_85),
.A2(n_92),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_85),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_85),
.B(n_245),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_90),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_90),
.B(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_136),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_97),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_97),
.B(n_187),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_162),
.C(n_174),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_103),
.B(n_126),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_99),
.B(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_99),
.A2(n_103),
.B1(n_124),
.B2(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.C(n_113),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_107),
.A2(n_116),
.B1(n_117),
.B2(n_132),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_108),
.Y(n_263)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_113),
.A2(n_133),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_113),
.A2(n_133),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_113),
.A2(n_133),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_113),
.B(n_262),
.C(n_264),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_113),
.B(n_269),
.C(n_274),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_117),
.B1(n_169),
.B2(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_123),
.Y(n_213)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_132),
.C(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B(n_121),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_121),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.C(n_137),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_133),
.B(n_213),
.C(n_215),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_137),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_138),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_202),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_197),
.B(n_201),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_165),
.B(n_196),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_153),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_162),
.C(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_156),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_164),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_209),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_191),
.B(n_195),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_176),
.B(n_190),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_171),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B(n_189),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_188),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_204),
.B(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_217),
.B2(n_218),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_212),
.C(n_218),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_217),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_222),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_229),
.C(n_237),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_234),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_234),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_248),
.B(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_240),
.B(n_241),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_253),
.B2(n_254),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_247),
.C(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_258),
.C(n_265),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_258),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_267),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_266),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);


endmodule