module real_aes_15548_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_0), .Y(n_572) );
AND2x4_ASAP7_75t_L g121 ( .A(n_1), .B(n_122), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_2), .A2(n_4), .B1(n_275), .B2(n_276), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_3), .A2(n_22), .B1(n_175), .B2(n_256), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_5), .A2(n_54), .B1(n_183), .B2(n_212), .Y(n_211) );
BUFx3_ASAP7_75t_L g606 ( .A(n_6), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_7), .A2(n_14), .B1(n_146), .B2(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g122 ( .A(n_8), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_9), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_10), .B(n_181), .Y(n_620) );
BUFx2_ASAP7_75t_L g110 ( .A(n_11), .Y(n_110) );
OR2x2_ASAP7_75t_L g856 ( .A(n_11), .B(n_33), .Y(n_856) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_13), .Y(n_886) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_15), .B(n_217), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_16), .B(n_190), .Y(n_588) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_16), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_17), .A2(n_87), .B1(n_217), .B2(n_256), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_18), .A2(n_60), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_18), .Y(n_130) );
INVx1_ASAP7_75t_L g874 ( .A(n_19), .Y(n_874) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_20), .A2(n_50), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_21), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_23), .B(n_175), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_24), .B(n_151), .Y(n_231) );
INVx4_ASAP7_75t_R g199 ( .A(n_25), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_26), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_27), .A2(n_885), .B(n_890), .Y(n_889) );
AO32x2_ASAP7_75t_L g531 ( .A1(n_28), .A2(n_169), .A3(n_170), .B1(n_532), .B2(n_535), .Y(n_531) );
AO32x1_ASAP7_75t_L g636 ( .A1(n_28), .A2(n_169), .A3(n_170), .B1(n_532), .B2(n_535), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_29), .B(n_175), .Y(n_238) );
INVx1_ASAP7_75t_L g280 ( .A(n_30), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_SL g253 ( .A1(n_31), .A2(n_146), .B(n_150), .C(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_32), .A2(n_47), .B1(n_146), .B2(n_153), .Y(n_262) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_34), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_35), .A2(n_53), .B1(n_175), .B2(n_200), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_36), .A2(n_93), .B1(n_153), .B2(n_256), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_37), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g898 ( .A(n_38), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_39), .B(n_544), .Y(n_548) );
INVx1_ASAP7_75t_L g235 ( .A(n_40), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_41), .B(n_146), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_42), .A2(n_70), .B1(n_153), .B2(n_557), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_43), .Y(n_173) );
INVx2_ASAP7_75t_L g851 ( .A(n_44), .Y(n_851) );
INVx1_ASAP7_75t_L g116 ( .A(n_45), .Y(n_116) );
BUFx3_ASAP7_75t_L g854 ( .A(n_45), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_46), .B(n_550), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_48), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_49), .A2(n_86), .B1(n_146), .B2(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_51), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_52), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_55), .A2(n_80), .B1(n_219), .B2(n_544), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_56), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_57), .A2(n_84), .B1(n_217), .B2(n_256), .Y(n_602) );
INVx1_ASAP7_75t_L g159 ( .A(n_58), .Y(n_159) );
AND2x4_ASAP7_75t_L g161 ( .A(n_59), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g131 ( .A(n_60), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_61), .A2(n_92), .B1(n_153), .B2(n_273), .Y(n_272) );
AO22x1_ASAP7_75t_L g215 ( .A1(n_62), .A2(n_75), .B1(n_216), .B2(n_218), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_63), .B(n_256), .Y(n_619) );
INVx1_ASAP7_75t_L g162 ( .A(n_64), .Y(n_162) );
AND2x2_ASAP7_75t_L g257 ( .A(n_65), .B(n_169), .Y(n_257) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_66), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_67), .B(n_169), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_68), .A2(n_183), .B(n_210), .C(n_571), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_69), .B(n_256), .C(n_623), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_71), .B(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_72), .Y(n_248) );
AND2x2_ASAP7_75t_L g573 ( .A(n_73), .B(n_204), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_74), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_76), .B(n_175), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_77), .A2(n_98), .B1(n_217), .B2(n_219), .Y(n_595) );
INVx2_ASAP7_75t_L g151 ( .A(n_78), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_79), .B(n_176), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_81), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_82), .B(n_169), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_83), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_85), .B(n_157), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_88), .B(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_89), .A2(n_103), .B1(n_153), .B2(n_200), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_90), .B(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_91), .A2(n_128), .B1(n_129), .B2(n_132), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_91), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_94), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g120 ( .A(n_95), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_95), .B(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_96), .B(n_190), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_97), .A2(n_155), .B(n_183), .C(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g203 ( .A(n_99), .B(n_204), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g180 ( .A(n_100), .B(n_181), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_101), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
CKINVDCx14_ASAP7_75t_R g865 ( .A(n_101), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_102), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_897), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx10_ASAP7_75t_L g899 ( .A(n_108), .Y(n_899) );
AND2x6_ASAP7_75t_SL g108 ( .A(n_109), .B(n_113), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND3x2_ASAP7_75t_L g871 ( .A(n_115), .B(n_119), .C(n_855), .Y(n_871) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g883 ( .A(n_116), .Y(n_883) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g522 ( .A(n_120), .Y(n_522) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_846), .B(n_857), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_133), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
AOI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_520), .B1(n_523), .B2(n_843), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
XNOR2x1_ASAP7_75t_L g872 ( .A(n_135), .B(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_429), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_345), .C(n_376), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_311), .Y(n_137) );
AOI211x1_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_223), .B(n_266), .C(n_297), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_187), .Y(n_140) );
AND2x2_ASAP7_75t_L g452 ( .A(n_141), .B(n_327), .Y(n_452) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_166), .Y(n_141) );
INVx1_ASAP7_75t_L g337 ( .A(n_142), .Y(n_337) );
OR2x2_ASAP7_75t_L g458 ( .A(n_142), .B(n_309), .Y(n_458) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g294 ( .A(n_143), .B(n_167), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_143), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g326 ( .A(n_143), .Y(n_326) );
OR2x2_ASAP7_75t_L g357 ( .A(n_143), .B(n_188), .Y(n_357) );
AND2x2_ASAP7_75t_L g371 ( .A(n_143), .B(n_188), .Y(n_371) );
AND2x2_ASAP7_75t_L g408 ( .A(n_143), .B(n_364), .Y(n_408) );
AO31x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_156), .A3(n_160), .B(n_163), .Y(n_143) );
OAI22x1_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B1(n_152), .B2(n_154), .Y(n_144) );
INVx4_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
INVx1_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_147), .Y(n_217) );
INVx1_ASAP7_75t_L g219 ( .A(n_147), .Y(n_219) );
INVx1_ASAP7_75t_L g250 ( .A(n_147), .Y(n_250) );
INVx2_ASAP7_75t_L g256 ( .A(n_147), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_148), .A2(n_173), .B(n_174), .C(n_176), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_149), .A2(n_209), .B1(n_261), .B2(n_262), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_149), .A2(n_154), .B1(n_272), .B2(n_274), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_149), .A2(n_548), .B(n_549), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_149), .A2(n_209), .B1(n_556), .B2(n_558), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_149), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_149), .A2(n_150), .B1(n_602), .B2(n_603), .Y(n_601) );
INVx6_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_150), .A2(n_180), .B(n_182), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_150), .B(n_215), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_150), .A2(n_208), .B(n_215), .C(n_221), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_150), .A2(n_252), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_150), .A2(n_619), .B(n_620), .Y(n_618) );
BUFx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g155 ( .A(n_151), .Y(n_155) );
INVx2_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx1_ASAP7_75t_L g234 ( .A(n_151), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_153), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g275 ( .A(n_153), .Y(n_275) );
INVx2_ASAP7_75t_L g546 ( .A(n_153), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_154), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g569 ( .A(n_155), .Y(n_569) );
INVx1_ASAP7_75t_SL g594 ( .A(n_155), .Y(n_594) );
INVx2_ASAP7_75t_L g616 ( .A(n_156), .Y(n_616) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
INVx2_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
OAI21xp33_ASAP7_75t_L g221 ( .A1(n_157), .A2(n_213), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_158), .Y(n_170) );
INVx2_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
BUFx10_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx10_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
INVx1_ASAP7_75t_L g278 ( .A(n_161), .Y(n_278) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_161), .A2(n_554), .A3(n_555), .B(n_559), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx2_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
BUFx2_ASAP7_75t_L g244 ( .A(n_165), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_165), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_165), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_165), .B(n_597), .Y(n_596) );
BUFx2_ASAP7_75t_L g288 ( .A(n_166), .Y(n_288) );
AND2x2_ASAP7_75t_L g339 ( .A(n_166), .B(n_205), .Y(n_339) );
AND2x2_ASAP7_75t_L g482 ( .A(n_166), .B(n_188), .Y(n_482) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g306 ( .A(n_167), .Y(n_306) );
AND2x2_ASAP7_75t_L g325 ( .A(n_167), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g362 ( .A(n_167), .Y(n_362) );
AND2x2_ASAP7_75t_L g386 ( .A(n_167), .B(n_188), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_168), .B(n_171), .Y(n_167) );
NOR2x1_ASAP7_75t_L g184 ( .A(n_169), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g263 ( .A(n_169), .Y(n_263) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g239 ( .A(n_170), .B(n_186), .Y(n_239) );
INVx2_ASAP7_75t_SL g540 ( .A(n_170), .Y(n_540) );
BUFx3_ASAP7_75t_L g554 ( .A(n_170), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_170), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_170), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_170), .B(n_605), .Y(n_604) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_179), .B(n_184), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_175), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g557 ( .A(n_175), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_175), .A2(n_200), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx2_ASAP7_75t_SL g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_177), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_584) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx3_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_181), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_198) );
INVx2_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AO31x2_ASAP7_75t_L g259 ( .A1(n_186), .A2(n_260), .A3(n_263), .B(n_264), .Y(n_259) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_186), .A2(n_581), .B(n_584), .Y(n_580) );
AOI31xp67_ASAP7_75t_L g600 ( .A1(n_186), .A2(n_263), .A3(n_601), .B(n_604), .Y(n_600) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_186), .A2(n_618), .B(n_621), .Y(n_617) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_187), .Y(n_286) );
AND2x2_ASAP7_75t_L g347 ( .A(n_187), .B(n_336), .Y(n_347) );
INVx2_ASAP7_75t_L g479 ( .A(n_187), .Y(n_479) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_205), .Y(n_187) );
INVx1_ASAP7_75t_L g284 ( .A(n_188), .Y(n_284) );
AND2x4_ASAP7_75t_L g296 ( .A(n_188), .B(n_206), .Y(n_296) );
INVx2_ASAP7_75t_L g364 ( .A(n_188), .Y(n_364) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_192), .B(n_203), .Y(n_188) );
AOI21x1_ASAP7_75t_L g563 ( .A1(n_189), .A2(n_564), .B(n_573), .Y(n_563) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_197), .B(n_202), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx2_ASAP7_75t_L g212 ( .A(n_195), .Y(n_212) );
INVx1_ASAP7_75t_L g586 ( .A(n_200), .Y(n_586) );
AND2x2_ASAP7_75t_L g363 ( .A(n_205), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g370 ( .A(n_205), .Y(n_370) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g448 ( .A(n_206), .B(n_364), .Y(n_448) );
AOI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_214), .B(n_220), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B(n_213), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_209), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21x1_ASAP7_75t_L g542 ( .A1(n_209), .A2(n_543), .B(n_545), .Y(n_542) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g550 ( .A(n_217), .Y(n_550) );
OAI21xp33_ASAP7_75t_SL g230 ( .A1(n_218), .A2(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_219), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_222), .A2(n_246), .B(n_253), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_222), .A2(n_565), .B(n_570), .Y(n_564) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
OR2x2_ASAP7_75t_L g353 ( .A(n_225), .B(n_241), .Y(n_353) );
AND2x2_ASAP7_75t_L g491 ( .A(n_225), .B(n_435), .Y(n_491) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g268 ( .A(n_226), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g373 ( .A(n_226), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_226), .B(n_315), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_226), .B(n_291), .Y(n_428) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g285 ( .A(n_227), .Y(n_285) );
AND2x2_ASAP7_75t_L g301 ( .A(n_227), .B(n_302), .Y(n_301) );
NAND2x1p5_ASAP7_75t_SL g314 ( .A(n_227), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g322 ( .A(n_227), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_227), .B(n_291), .Y(n_393) );
AND2x2_ASAP7_75t_L g441 ( .A(n_227), .B(n_270), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_227), .B(n_269), .Y(n_484) );
BUFx2_ASAP7_75t_L g503 ( .A(n_227), .Y(n_503) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B(n_239), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
BUFx4f_ASAP7_75t_L g252 ( .A(n_234), .Y(n_252) );
INVx1_ASAP7_75t_L g623 ( .A(n_234), .Y(n_623) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g287 ( .A(n_241), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g400 ( .A(n_241), .Y(n_400) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_258), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_242), .B(n_270), .Y(n_303) );
INVx2_ASAP7_75t_L g315 ( .A(n_242), .Y(n_315) );
AND2x2_ASAP7_75t_L g351 ( .A(n_242), .B(n_259), .Y(n_351) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g291 ( .A(n_243), .Y(n_291) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_257), .Y(n_243) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_271), .A3(n_277), .B(n_279), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_252), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g276 ( .A(n_250), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g581 ( .A1(n_252), .A2(n_276), .B(n_582), .C(n_583), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_SL g544 ( .A(n_256), .Y(n_544) );
INVx1_ASAP7_75t_L g375 ( .A(n_258), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_258), .B(n_270), .Y(n_392) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g302 ( .A(n_259), .Y(n_302) );
OR2x2_ASAP7_75t_L g334 ( .A(n_259), .B(n_270), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_259), .B(n_270), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_287), .B1(n_289), .B2(n_293), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_281), .B1(n_285), .B2(n_286), .Y(n_267) );
INVx2_ASAP7_75t_L g292 ( .A(n_268), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_268), .B(n_351), .Y(n_365) );
AND2x2_ASAP7_75t_L g399 ( .A(n_268), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
INVx1_ASAP7_75t_L g323 ( .A(n_270), .Y(n_323) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_277), .A2(n_554), .A3(n_592), .B(n_596), .Y(n_591) );
INVx2_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_SL g535 ( .A(n_278), .Y(n_535) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g457 ( .A(n_283), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
AND3x1_ASAP7_75t_L g442 ( .A(n_284), .B(n_305), .C(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g398 ( .A(n_285), .Y(n_398) );
AND2x4_ASAP7_75t_L g434 ( .A(n_285), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g472 ( .A(n_288), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_289), .Y(n_476) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
OR2x2_ASAP7_75t_L g449 ( .A(n_290), .B(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_290), .Y(n_497) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g397 ( .A(n_291), .B(n_375), .Y(n_397) );
AND2x2_ASAP7_75t_L g439 ( .A(n_291), .B(n_306), .Y(n_439) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_291), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_295), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_294), .A2(n_295), .B(n_359), .C(n_365), .Y(n_358) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_294), .B(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_294), .B(n_452), .Y(n_498) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_296), .B(n_325), .Y(n_344) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_304), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_303), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_304), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AND2x2_ASAP7_75t_L g354 ( .A(n_305), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_305), .B(n_371), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_305), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_305), .B(n_363), .Y(n_519) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g502 ( .A(n_306), .Y(n_502) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_324), .B(n_329), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_318), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
OAI33xp33_ASAP7_75t_L g378 ( .A1(n_314), .A2(n_319), .A3(n_379), .B1(n_380), .B2(n_382), .B3(n_383), .Y(n_378) );
OR2x2_ASAP7_75t_L g510 ( .A(n_314), .B(n_334), .Y(n_510) );
INVx2_ASAP7_75t_L g512 ( .A(n_314), .Y(n_512) );
INVx1_ASAP7_75t_L g333 ( .A(n_315), .Y(n_333) );
OR2x2_ASAP7_75t_L g374 ( .A(n_315), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g382 ( .A(n_319), .Y(n_382) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_319), .B(n_501), .C(n_503), .Y(n_500) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_320), .B(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_320), .B(n_484), .Y(n_488) );
AND2x4_ASAP7_75t_L g517 ( .A(n_320), .B(n_518), .Y(n_517) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g343 ( .A(n_322), .Y(n_343) );
OR2x2_ASAP7_75t_L g349 ( .A(n_322), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g462 ( .A(n_322), .B(n_397), .Y(n_462) );
INVx1_ASAP7_75t_L g518 ( .A(n_322), .Y(n_518) );
AND2x4_ASAP7_75t_SL g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
INVx1_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
AND2x2_ASAP7_75t_L g425 ( .A(n_326), .B(n_328), .Y(n_425) );
INVx1_ASAP7_75t_L g465 ( .A(n_327), .Y(n_465) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g356 ( .A(n_328), .B(n_357), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_335), .B1(n_342), .B2(n_344), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g421 ( .A(n_334), .Y(n_421) );
INVx2_ASAP7_75t_L g435 ( .A(n_334), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B(n_339), .C(n_340), .Y(n_335) );
INVx1_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_337), .B(n_362), .Y(n_464) );
OR2x2_ASAP7_75t_L g480 ( .A(n_337), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g493 ( .A(n_337), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_339), .B(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_366), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_352), .B2(n_354), .C(n_358), .Y(n_346) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI32xp33_ASAP7_75t_L g515 ( .A1(n_349), .A2(n_446), .A3(n_464), .B1(n_516), .B2(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g485 ( .A(n_351), .Y(n_485) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_354), .A2(n_367), .B(n_372), .Y(n_366) );
NAND2x1_ASAP7_75t_L g514 ( .A(n_355), .B(n_502), .Y(n_514) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
AND2x2_ASAP7_75t_L g508 ( .A(n_361), .B(n_389), .Y(n_508) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g456 ( .A(n_362), .Y(n_456) );
INVx2_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
AND2x2_ASAP7_75t_L g385 ( .A(n_369), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g404 ( .A(n_370), .Y(n_404) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_394), .C(n_405), .D(n_416), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_385), .B1(n_387), .B2(n_390), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_379), .A2(n_507), .B1(n_509), .B2(n_510), .Y(n_506) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g489 ( .A(n_384), .B(n_448), .Y(n_489) );
AND2x2_ASAP7_75t_L g492 ( .A(n_386), .B(n_493), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_387), .A2(n_406), .B1(n_410), .B2(n_413), .Y(n_405) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OR2x2_ASAP7_75t_L g427 ( .A(n_392), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g411 ( .A(n_393), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g422 ( .A(n_393), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_399), .B(n_401), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_395), .A2(n_500), .B(n_504), .C(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g474 ( .A(n_397), .Y(n_474) );
AND2x4_ASAP7_75t_L g467 ( .A(n_400), .B(n_441), .Y(n_467) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_407), .A2(n_433), .B(n_436), .Y(n_432) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g438 ( .A(n_408), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_408), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g414 ( .A(n_412), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_414), .A2(n_445), .B1(n_449), .B2(n_451), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_423), .B2(n_426), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_421), .Y(n_437) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_494), .Y(n_429) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_431), .B(n_453), .C(n_469), .D(n_486), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_444), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g496 ( .A(n_434), .B(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_440), .B2(n_442), .Y(n_436) );
INVxp67_ASAP7_75t_L g460 ( .A(n_440), .Y(n_460) );
BUFx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g450 ( .A(n_441), .Y(n_450) );
AND2x2_ASAP7_75t_L g473 ( .A(n_441), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_459), .B(n_461), .Y(n_453) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x6_ASAP7_75t_L g478 ( .A(n_456), .B(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g475 ( .A(n_457), .Y(n_475) );
OAI32xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .A3(n_465), .B1(n_466), .B2(n_468), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B1(n_475), .B2(n_476), .C(n_477), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B(n_483), .Y(n_477) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g509 ( .A(n_488), .Y(n_509) );
INVx1_ASAP7_75t_L g505 ( .A(n_489), .Y(n_505) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g494 ( .A1(n_495), .A2(n_498), .B(n_499), .C(n_511), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVxp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_515), .Y(n_511) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
BUFx8_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_522), .Y(n_845) );
AND2x2_ASAP7_75t_L g895 ( .A(n_522), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NOR2x1p5_ASAP7_75t_L g524 ( .A(n_525), .B(n_751), .Y(n_524) );
NAND4xp75_ASAP7_75t_L g525 ( .A(n_526), .B(n_648), .C(n_682), .D(n_731), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_574), .B(n_607), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_536), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g727 ( .A(n_530), .Y(n_727) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g612 ( .A(n_531), .B(n_538), .Y(n_612) );
AND2x4_ASAP7_75t_L g643 ( .A(n_531), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g664 ( .A(n_531), .Y(n_664) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_535), .A2(n_542), .B(n_547), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_536), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_552), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_537), .B(n_678), .Y(n_755) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_537), .Y(n_782) );
OR2x2_ASAP7_75t_L g831 ( .A(n_537), .B(n_635), .Y(n_831) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g647 ( .A(n_538), .Y(n_647) );
INVx3_ASAP7_75t_L g655 ( .A(n_538), .Y(n_655) );
OR2x2_ASAP7_75t_L g663 ( .A(n_538), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g691 ( .A(n_538), .B(n_661), .Y(n_691) );
INVx1_ASAP7_75t_L g702 ( .A(n_538), .Y(n_702) );
AND2x2_ASAP7_75t_L g723 ( .A(n_538), .B(n_664), .Y(n_723) );
INVxp67_ASAP7_75t_L g747 ( .A(n_538), .Y(n_747) );
BUFx2_ASAP7_75t_L g791 ( .A(n_538), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_538), .B(n_553), .Y(n_800) );
AND2x2_ASAP7_75t_L g807 ( .A(n_538), .B(n_808), .Y(n_807) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_551), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_546), .A2(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g665 ( .A(n_552), .B(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_552), .A2(n_577), .B1(n_781), .B2(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
OR2x2_ASAP7_75t_L g635 ( .A(n_553), .B(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g644 ( .A(n_553), .Y(n_644) );
AND2x2_ASAP7_75t_L g656 ( .A(n_553), .B(n_636), .Y(n_656) );
AND2x2_ASAP7_75t_L g714 ( .A(n_553), .B(n_562), .Y(n_714) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
INVx1_ASAP7_75t_L g705 ( .A(n_562), .Y(n_705) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_562), .Y(n_808) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g661 ( .A(n_563), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_566), .B(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_589), .Y(n_575) );
AND2x2_ASAP7_75t_L g762 ( .A(n_576), .B(n_708), .Y(n_762) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI32xp33_ASAP7_75t_L g792 ( .A1(n_577), .A2(n_685), .A3(n_759), .B1(n_793), .B2(n_795), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_577), .B(n_822), .Y(n_821) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g614 ( .A(n_578), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g631 ( .A(n_578), .B(n_591), .Y(n_631) );
BUFx2_ASAP7_75t_L g650 ( .A(n_578), .Y(n_650) );
INVx1_ASAP7_75t_L g697 ( .A(n_578), .Y(n_697) );
AND2x2_ASAP7_75t_L g730 ( .A(n_578), .B(n_709), .Y(n_730) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B(n_588), .Y(n_578) );
OA21x2_ASAP7_75t_L g676 ( .A1(n_579), .A2(n_580), .B(n_588), .Y(n_676) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g613 ( .A(n_590), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g818 ( .A(n_590), .B(n_702), .Y(n_818) );
INVx1_ASAP7_75t_L g822 ( .A(n_590), .Y(n_822) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_598), .Y(n_590) );
INVx2_ASAP7_75t_L g646 ( .A(n_591), .Y(n_646) );
AND2x2_ASAP7_75t_L g670 ( .A(n_591), .B(n_629), .Y(n_670) );
AND2x2_ASAP7_75t_L g681 ( .A(n_591), .B(n_676), .Y(n_681) );
INVx1_ASAP7_75t_L g688 ( .A(n_591), .Y(n_688) );
AND2x2_ASAP7_75t_L g696 ( .A(n_591), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
AND2x2_ASAP7_75t_L g775 ( .A(n_591), .B(n_598), .Y(n_775) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g639 ( .A(n_599), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g629 ( .A(n_600), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_613), .B1(n_626), .B2(n_632), .C(n_637), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_609), .A2(n_759), .B(n_762), .Y(n_758) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
AND2x4_ASAP7_75t_L g834 ( .A(n_610), .B(n_634), .Y(n_834) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g678 ( .A(n_611), .B(n_644), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_612), .B(n_713), .Y(n_712) );
BUFx2_ASAP7_75t_L g743 ( .A(n_612), .Y(n_743) );
OR2x2_ASAP7_75t_L g687 ( .A(n_614), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g749 ( .A(n_614), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g820 ( .A(n_614), .Y(n_820) );
AND2x2_ASAP7_75t_L g628 ( .A(n_615), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g777 ( .A(n_615), .B(n_676), .Y(n_777) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_625), .Y(n_615) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_616), .A2(n_617), .B(n_625), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_626), .A2(n_658), .B1(n_659), .B2(n_668), .C(n_677), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_626), .A2(n_741), .B1(n_754), .B2(n_756), .C(n_758), .Y(n_753) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND2x2_ASAP7_75t_L g680 ( .A(n_628), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_629), .B(n_676), .Y(n_693) );
INVx2_ASAP7_75t_L g699 ( .A(n_629), .Y(n_699) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_632), .A2(n_764), .B1(n_769), .B2(n_773), .C(n_778), .Y(n_763) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g815 ( .A(n_635), .B(n_785), .Y(n_815) );
INVx1_ASAP7_75t_L g667 ( .A(n_636), .Y(n_667) );
INVx1_ASAP7_75t_L g704 ( .A(n_636), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g653 ( .A(n_639), .Y(n_653) );
OR2x2_ASAP7_75t_L g716 ( .A(n_639), .B(n_652), .Y(n_716) );
INVx2_ASAP7_75t_L g729 ( .A(n_639), .Y(n_729) );
INVx2_ASAP7_75t_L g674 ( .A(n_640), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g679 ( .A(n_643), .Y(n_679) );
AND2x4_ASAP7_75t_L g685 ( .A(n_643), .B(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_643), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g759 ( .A(n_643), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g836 ( .A(n_643), .B(n_791), .Y(n_836) );
AND2x2_ASAP7_75t_L g660 ( .A(n_644), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g722 ( .A(n_644), .Y(n_722) );
INVx1_ASAP7_75t_L g781 ( .A(n_644), .Y(n_781) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_SL g652 ( .A(n_646), .Y(n_652) );
AND2x2_ASAP7_75t_L g694 ( .A(n_646), .B(n_673), .Y(n_694) );
AND2x2_ASAP7_75t_L g768 ( .A(n_647), .B(n_722), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_654), .B(n_657), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g734 ( .A(n_650), .Y(n_734) );
AND2x2_ASAP7_75t_L g801 ( .A(n_650), .B(n_729), .Y(n_801) );
AND2x2_ASAP7_75t_L g816 ( .A(n_650), .B(n_775), .Y(n_816) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_L g770 ( .A(n_652), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_652), .B(n_777), .Y(n_787) );
OAI33xp33_ASAP7_75t_L g824 ( .A1(n_652), .A2(n_726), .A3(n_794), .B1(n_825), .B2(n_826), .B3(n_827), .Y(n_824) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_655), .B(n_661), .Y(n_785) );
AND2x2_ASAP7_75t_L g813 ( .A(n_656), .B(n_761), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_665), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g686 ( .A(n_661), .Y(n_686) );
INVx1_ASAP7_75t_L g761 ( .A(n_661), .Y(n_761) );
OAI32xp33_ASAP7_75t_L g706 ( .A1(n_662), .A2(n_687), .A3(n_707), .B1(n_710), .B2(n_712), .Y(n_706) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g741 ( .A(n_663), .B(n_686), .Y(n_741) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g719 ( .A(n_667), .Y(n_719) );
INVx2_ASAP7_75t_L g767 ( .A(n_667), .Y(n_767) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g750 ( .A(n_670), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_671), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g810 ( .A(n_671), .B(n_757), .Y(n_810) );
INVx2_ASAP7_75t_L g841 ( .A(n_671), .Y(n_841) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g756 ( .A(n_672), .B(n_757), .Y(n_756) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
AND2x2_ASAP7_75t_L g698 ( .A(n_673), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g740 ( .A(n_674), .Y(n_740) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_680), .Y(n_677) );
INVx2_ASAP7_75t_L g748 ( .A(n_678), .Y(n_748) );
AND2x2_ASAP7_75t_L g732 ( .A(n_679), .B(n_733), .Y(n_732) );
NOR3x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_706), .C(n_715), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_687), .B(n_689), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_686), .B(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_688), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B1(n_695), .B2(n_700), .Y(n_689) );
INVx3_ASAP7_75t_L g724 ( .A(n_691), .Y(n_724) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVxp67_ASAP7_75t_L g737 ( .A(n_693), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_693), .B(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_L g838 ( .A(n_696), .B(n_729), .Y(n_838) );
AND2x2_ASAP7_75t_L g708 ( .A(n_699), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g757 ( .A(n_699), .Y(n_757) );
INVx1_ASAP7_75t_L g794 ( .A(n_699), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_699), .B(n_740), .Y(n_828) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g825 ( .A(n_703), .Y(n_825) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g711 ( .A(n_705), .Y(n_711) );
AND2x2_ASAP7_75t_L g837 ( .A(n_708), .B(n_777), .Y(n_837) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx2_ASAP7_75t_L g745 ( .A(n_714), .Y(n_745) );
AND2x2_ASAP7_75t_L g842 ( .A(n_714), .B(n_723), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_725), .B2(n_728), .Y(n_715) );
AOI211xp5_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_720), .B(n_723), .C(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g799 ( .A(n_719), .B(n_800), .Y(n_799) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp33_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g733 ( .A(n_729), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g811 ( .A(n_730), .B(n_772), .Y(n_811) );
INVx1_ASAP7_75t_L g826 ( .A(n_730), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .C(n_742), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_741), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g772 ( .A(n_740), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B(n_746), .C(n_749), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_743), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_803), .Y(n_751) );
NOR3xp33_ASAP7_75t_SL g752 ( .A(n_753), .B(n_763), .C(n_788), .Y(n_752) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_759), .A2(n_798), .B1(n_801), .B2(n_802), .Y(n_797) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
AND2x2_ASAP7_75t_L g783 ( .A(n_766), .B(n_784), .Y(n_783) );
AND2x4_ASAP7_75t_L g806 ( .A(n_766), .B(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OR2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g802 ( .A(n_771), .Y(n_802) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_777), .B(n_794), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_783), .B(n_786), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_783), .A2(n_838), .B1(n_840), .B2(n_842), .Y(n_839) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI21xp33_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_792), .B(n_797), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_790), .B(n_834), .Y(n_833) );
BUFx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g829 ( .A(n_800), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_802), .A2(n_824), .B1(n_829), .B2(n_830), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_832), .Y(n_803) );
OAI211xp5_ASAP7_75t_SL g804 ( .A1(n_805), .A2(n_809), .B(n_812), .C(n_823), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NOR2x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
O2A1O1Ixp5_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_814), .B(n_816), .C(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_815), .A2(n_818), .B1(n_819), .B2(n_821), .Y(n_817) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_826), .A2(n_833), .B(n_835), .C(n_839), .Y(n_832) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx8_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
BUFx12f_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVxp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_848), .Y(n_847) );
BUFx12f_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
AND2x6_ASAP7_75t_SL g849 ( .A(n_850), .B(n_852), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx3_ASAP7_75t_L g861 ( .A(n_851), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_851), .B(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_854), .B(n_856), .Y(n_896) );
AND2x6_ASAP7_75t_SL g881 ( .A(n_855), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_862), .B(n_889), .Y(n_857) );
INVx1_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
CKINVDCx11_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_868), .B(n_876), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_864), .B(n_878), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_872), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OAI21xp33_ASAP7_75t_L g876 ( .A1(n_872), .A2(n_877), .B(n_884), .Y(n_876) );
XOR2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
INVx4_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx3_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
CKINVDCx8_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
INVx4_ASAP7_75t_L g888 ( .A(n_881), .Y(n_888) );
INVxp67_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
BUFx12f_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx10_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NOR2xp33_ASAP7_75t_R g897 ( .A(n_898), .B(n_899), .Y(n_897) );
endmodule