module fake_jpeg_12141_n_494 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_50),
.B(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_59),
.Y(n_145)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_63),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_10),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_74),
.Y(n_154)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_10),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_21),
.Y(n_83)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_46),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_26),
.B1(n_44),
.B2(n_46),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_118),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_44),
.B1(n_46),
.B2(n_38),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_43),
.B1(n_44),
.B2(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_110),
.B(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_39),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_44),
.B1(n_38),
.B2(n_29),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_39),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_128),
.B(n_143),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_43),
.B1(n_27),
.B2(n_30),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_135),
.B1(n_139),
.B2(n_60),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_35),
.B1(n_21),
.B2(n_30),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_75),
.A2(n_30),
.B1(n_27),
.B2(n_45),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_20),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_66),
.A2(n_30),
.B1(n_27),
.B2(n_35),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_57),
.B1(n_64),
.B2(n_58),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_53),
.B(n_45),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_69),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_157),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_159),
.Y(n_222)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_93),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_161),
.B(n_34),
.C(n_11),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_162),
.B(n_173),
.Y(n_235)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_166),
.A2(n_197),
.B1(n_202),
.B2(n_207),
.Y(n_234)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_103),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_111),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_171),
.A2(n_190),
.B1(n_196),
.B2(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_104),
.B(n_47),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_174),
.B(n_186),
.Y(n_238)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_42),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_184),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_61),
.B1(n_92),
.B2(n_70),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_182),
.A2(n_208),
.B1(n_34),
.B2(n_1),
.Y(n_254)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_40),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_102),
.B(n_42),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_31),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_192),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_100),
.A2(n_68),
.B1(n_67),
.B2(n_89),
.Y(n_190)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_74),
.A3(n_21),
.B1(n_33),
.B2(n_41),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_198),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_31),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_95),
.A2(n_83),
.B(n_21),
.C(n_24),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_34),
.B(n_41),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_135),
.A2(n_88),
.B1(n_87),
.B2(n_79),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_97),
.A2(n_20),
.B1(n_47),
.B2(n_40),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_201),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_0),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_0),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_97),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_126),
.A2(n_84),
.B1(n_94),
.B2(n_91),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_107),
.B(n_56),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_145),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_210),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_126),
.A2(n_35),
.B1(n_32),
.B2(n_82),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_132),
.A2(n_41),
.B1(n_33),
.B2(n_32),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_136),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_209),
.Y(n_257)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_96),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_211),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_122),
.A2(n_41),
.B1(n_33),
.B2(n_24),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_140),
.B1(n_24),
.B2(n_34),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_138),
.B1(n_119),
.B2(n_101),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_217),
.B(n_251),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_98),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_256),
.C(n_188),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_232),
.B1(n_236),
.B2(n_203),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_166),
.A2(n_118),
.B1(n_105),
.B2(n_138),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_226),
.A2(n_244),
.B1(n_254),
.B2(n_261),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_164),
.A2(n_161),
.B1(n_196),
.B2(n_189),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_161),
.A2(n_105),
.B1(n_119),
.B2(n_117),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_185),
.A2(n_117),
.B1(n_146),
.B2(n_24),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_144),
.B(n_130),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_237),
.A2(n_241),
.B(n_193),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_184),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_41),
.B1(n_34),
.B2(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_0),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_169),
.B(n_11),
.C(n_16),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_0),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_170),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_208),
.B1(n_181),
.B2(n_176),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_264),
.A2(n_280),
.B1(n_287),
.B2(n_222),
.Y(n_332)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_257),
.A2(n_167),
.B1(n_178),
.B2(n_194),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_180),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_276),
.C(n_278),
.Y(n_317)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

BUFx24_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_216),
.A2(n_209),
.A3(n_199),
.B1(n_172),
.B2(n_157),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_271),
.A2(n_288),
.B(n_231),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_273),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_165),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_274),
.B(n_279),
.Y(n_335)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_155),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_217),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_221),
.B(n_156),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_210),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_223),
.A2(n_187),
.B1(n_198),
.B2(n_160),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_228),
.B(n_163),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_209),
.C(n_175),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_246),
.C(n_260),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_177),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_291),
.Y(n_320)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_213),
.A2(n_183),
.B1(n_201),
.B2(n_211),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_205),
.B1(n_6),
.B2(n_12),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_290),
.A2(n_292),
.B1(n_299),
.B2(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_0),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_234),
.A2(n_6),
.B1(n_15),
.B2(n_3),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_214),
.B(n_6),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_260),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_297),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_252),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_1),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_304),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_241),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_300),
.A2(n_301),
.B1(n_305),
.B2(n_306),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_257),
.A2(n_13),
.B1(n_15),
.B2(n_3),
.Y(n_301)
);

NOR2xp67_ASAP7_75t_R g302 ( 
.A(n_251),
.B(n_3),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_240),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_248),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_1),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_265),
.A2(n_237),
.B1(n_217),
.B2(n_225),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_309),
.A2(n_321),
.B1(n_327),
.B2(n_334),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_263),
.B(n_256),
.CI(n_249),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_231),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_315),
.A2(n_287),
.B1(n_280),
.B2(n_286),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_265),
.A2(n_249),
.B(n_260),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_324),
.B(n_342),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_273),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_323),
.C(n_330),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_224),
.B(n_246),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_264),
.A2(n_215),
.B1(n_255),
.B2(n_240),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_329),
.B(n_345),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_272),
.A2(n_217),
.B1(n_219),
.B2(n_215),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_337),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_272),
.A2(n_289),
.B1(n_292),
.B2(n_285),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_222),
.B1(n_259),
.B2(n_233),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_336),
.A2(n_227),
.B1(n_2),
.B2(n_14),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_259),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_270),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_340),
.B(n_341),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_275),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_281),
.A2(n_227),
.B(n_247),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_276),
.B(n_233),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_281),
.C(n_291),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_284),
.B1(n_281),
.B2(n_290),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_346),
.A2(n_359),
.B1(n_361),
.B2(n_364),
.Y(n_388)
);

XOR2x2_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_278),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_310),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_351),
.C(n_353),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_283),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_354),
.A2(n_355),
.B1(n_343),
.B2(n_352),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_303),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_362),
.C(n_369),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_325),
.A2(n_299),
.B1(n_304),
.B2(n_298),
.Y(n_359)
);

INVx3_ASAP7_75t_SL g360 ( 
.A(n_333),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_366),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_337),
.A2(n_295),
.B1(n_296),
.B2(n_266),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_302),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_363),
.B(n_326),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_247),
.B1(n_227),
.B2(n_2),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_365),
.A2(n_338),
.B1(n_313),
.B2(n_322),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_320),
.B(n_2),
.Y(n_367)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

OAI32xp33_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_4),
.A3(n_14),
.B1(n_17),
.B2(n_320),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_370),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_4),
.C(n_17),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_307),
.Y(n_371)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_372),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_4),
.C(n_345),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_313),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_318),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_329),
.A2(n_331),
.B(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_375),
.B(n_309),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_316),
.A2(n_311),
.B1(n_315),
.B2(n_331),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_311),
.B1(n_315),
.B2(n_326),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_314),
.B(n_335),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_378),
.Y(n_393)
);

AOI21xp33_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_357),
.B(n_368),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_383),
.B(n_396),
.Y(n_411)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_359),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_374),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_387),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_390),
.A2(n_397),
.B1(n_358),
.B2(n_367),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_355),
.A2(n_352),
.B1(n_354),
.B2(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_395),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_353),
.B(n_322),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_346),
.A2(n_338),
.B1(n_339),
.B2(n_312),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_339),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_401),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_376),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_399),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_348),
.B(n_347),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_347),
.B(n_312),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_404),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_318),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_369),
.C(n_375),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_377),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_410),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_426),
.B1(n_428),
.B2(n_384),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_357),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_392),
.Y(n_436)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_393),
.B1(n_389),
.B2(n_394),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_362),
.C(n_371),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.C(n_423),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_372),
.C(n_364),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_365),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_396),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_360),
.C(n_370),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_360),
.C(n_366),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_392),
.C(n_387),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_308),
.B1(n_349),
.B2(n_390),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_388),
.A2(n_308),
.B1(n_397),
.B2(n_379),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_413),
.A2(n_417),
.B1(n_427),
.B2(n_428),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_432),
.A2(n_446),
.B1(n_445),
.B2(n_430),
.Y(n_455)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_409),
.Y(n_435)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_439),
.C(n_421),
.Y(n_462)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_440),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_391),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_441),
.A2(n_415),
.B1(n_412),
.B2(n_419),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_418),
.A2(n_394),
.B1(n_400),
.B2(n_382),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_443),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_423),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_391),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_421),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_417),
.A2(n_383),
.B1(n_387),
.B2(n_308),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_410),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_414),
.B(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_408),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_461),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_462),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_455),
.A2(n_445),
.B1(n_439),
.B2(n_432),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_458),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_453),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_459),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_468),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_434),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_434),
.C(n_436),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_470),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_424),
.C(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_454),
.C(n_452),
.Y(n_471)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_472),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_440),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_466),
.A2(n_469),
.B(n_464),
.Y(n_474)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_480),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_471),
.A2(n_460),
.B1(n_450),
.B2(n_470),
.Y(n_477)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_477),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_463),
.B(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_479),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_476),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_476),
.Y(n_485)
);

A2O1A1O1Ixp25_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_481),
.B(n_473),
.C(n_475),
.D(n_472),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_483),
.A2(n_478),
.B(n_463),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_487),
.B(n_480),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_457),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_489),
.C(n_455),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_473),
.C(n_453),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_449),
.B(n_431),
.Y(n_492)
);

AOI31xp33_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_453),
.A3(n_449),
.B(n_431),
.Y(n_493)
);

OAI311xp33_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_308),
.A3(n_411),
.B1(n_438),
.C1(n_459),
.Y(n_494)
);


endmodule