module fake_jpeg_21427_n_148 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_76),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_2),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_87),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_66),
.B1(n_49),
.B2(n_59),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_54),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_101),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_59),
.B1(n_49),
.B2(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_97),
.B1(n_100),
.B2(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_103),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_68),
.B1(n_64),
.B2(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_51),
.B1(n_57),
.B2(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_55),
.B1(n_62),
.B2(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_3),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_3),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_113),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_122),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_97),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_120),
.C(n_121),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_55),
.B(n_6),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_5),
.B(n_6),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_23),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_118),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_107),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_131),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_127),
.B1(n_128),
.B2(n_123),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_131),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_135),
.C(n_125),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.C(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_125),
.C(n_134),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_126),
.C(n_22),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_20),
.C(n_26),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_28),
.B(n_33),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_108),
.Y(n_148)
);


endmodule