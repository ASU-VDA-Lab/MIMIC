module fake_jpeg_29996_n_370 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_370);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_370;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_55),
.Y(n_84)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_21),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_47),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_28),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_93),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_28),
.B1(n_32),
.B2(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_103),
.B1(n_112),
.B2(n_106),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_44),
.B1(n_37),
.B2(n_32),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_36),
.B1(n_38),
.B2(n_22),
.Y(n_121)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_24),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_28),
.B1(n_32),
.B2(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_58),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_48),
.A2(n_38),
.B1(n_37),
.B2(n_46),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_134),
.Y(n_151)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_126),
.B1(n_140),
.B2(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_35),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_129),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_59),
.B1(n_66),
.B2(n_22),
.Y(n_126)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_75),
.B(n_24),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_49),
.B1(n_78),
.B2(n_99),
.Y(n_152)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_81),
.B(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_141),
.Y(n_161)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_91),
.A2(n_58),
.B1(n_49),
.B2(n_34),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_34),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_33),
.B1(n_43),
.B2(n_40),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_29),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_29),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_97),
.B1(n_103),
.B2(n_100),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_121),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_153),
.B1(n_119),
.B2(n_97),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_78),
.B1(n_73),
.B2(n_99),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_87),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_116),
.B(n_106),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_140),
.C(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_113),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_157),
.Y(n_199)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_125),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_188),
.CI(n_166),
.CON(n_193),
.SN(n_193)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_185),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_166),
.B1(n_162),
.B2(n_157),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_183),
.B(n_142),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_123),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_131),
.B(n_113),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_167),
.B1(n_165),
.B2(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_146),
.B(n_150),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_202),
.C(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_178),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_146),
.B(n_161),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_206),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_204),
.B1(n_180),
.B2(n_181),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_184),
.B1(n_187),
.B2(n_175),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_158),
.C(n_143),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_148),
.B1(n_168),
.B2(n_163),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_215),
.B1(n_200),
.B2(n_175),
.Y(n_247)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_224),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_180),
.B1(n_183),
.B2(n_179),
.Y(n_215)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_216),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_221),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_198),
.B(n_191),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_178),
.C(n_188),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_199),
.C(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_187),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_227),
.B1(n_197),
.B2(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_175),
.B1(n_173),
.B2(n_172),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_191),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_240),
.B(n_156),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_189),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_235),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_232),
.A2(n_213),
.B1(n_175),
.B2(n_208),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_192),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_248),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_191),
.B(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_221),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_169),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_226),
.B1(n_218),
.B2(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_168),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_143),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_159),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_262),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_252),
.A2(n_228),
.B1(n_234),
.B2(n_244),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_222),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_215),
.C(n_207),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_265),
.C(n_272),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_222),
.B1(n_213),
.B2(n_203),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_264),
.B1(n_238),
.B2(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_235),
.A2(n_216),
.B1(n_208),
.B2(n_124),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_158),
.C(n_156),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_43),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_176),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_27),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_164),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_160),
.C(n_134),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_160),
.C(n_155),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_274),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_228),
.B1(n_234),
.B2(n_238),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_281),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_272),
.B1(n_257),
.B2(n_268),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_253),
.B(n_216),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_273),
.C(n_258),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_117),
.B(n_136),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_255),
.B(n_252),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_124),
.B1(n_128),
.B2(n_87),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_30),
.B1(n_40),
.B2(n_125),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_144),
.B1(n_3),
.B2(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_266),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_176),
.Y(n_291)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_257),
.B(n_176),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_294),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_304),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_265),
.C(n_260),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_308),
.C(n_311),
.Y(n_325)
);

BUFx12_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_139),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_127),
.C(n_115),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_127),
.C(n_115),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_282),
.A2(n_288),
.B(n_289),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_128),
.C(n_73),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_316),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_284),
.B1(n_283),
.B2(n_307),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_275),
.Y(n_319)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_322),
.B(n_323),
.Y(n_333)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_301),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_328),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_283),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_274),
.B(n_301),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_329),
.A2(n_79),
.B(n_88),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_292),
.B(n_306),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_330),
.B(n_335),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_306),
.B1(n_281),
.B2(n_294),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_331),
.A2(n_334),
.B1(n_312),
.B2(n_133),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_82),
.B1(n_89),
.B2(n_100),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_2),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_2),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_336),
.B(n_7),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_318),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_339),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_312),
.C(n_88),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_342),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_79),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_344)
);

AO21x1_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_8),
.B(n_10),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_345),
.A2(n_69),
.B(n_9),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_346),
.B(n_347),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_331),
.A2(n_110),
.B(n_36),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_348),
.A2(n_334),
.B(n_9),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_354),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_352),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_343),
.B(n_8),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_341),
.B(n_342),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_353),
.B(n_356),
.Y(n_358)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_349),
.A2(n_345),
.B(n_344),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_361),
.B(n_11),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_69),
.C(n_10),
.Y(n_361)
);

AOI322xp5_ASAP7_75t_L g363 ( 
.A1(n_360),
.A2(n_8),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_363),
.A2(n_12),
.B(n_13),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_357),
.Y(n_365)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_365),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_362),
.B(n_366),
.Y(n_368)
);

OAI321xp33_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_13),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g370 ( 
.A(n_369),
.B(n_16),
.CI(n_17),
.CON(n_370),
.SN(n_370)
);


endmodule