module fake_jpeg_11640_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_12),
.B(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_4),
.Y(n_71)
);

BUFx6f_ASAP7_75t_SL g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_21),
.B(n_46),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_53),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_3),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_51),
.B1(n_57),
.B2(n_52),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_93),
.B1(n_24),
.B2(n_44),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_63),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_51),
.B1(n_57),
.B2(n_61),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_60),
.CI(n_64),
.CON(n_94),
.SN(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_98),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_54),
.B(n_75),
.C(n_62),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_54),
.B(n_61),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_1),
.C(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_59),
.B1(n_68),
.B2(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_27),
.B1(n_43),
.B2(n_41),
.Y(n_118)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_81),
.B(n_58),
.C(n_70),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_114),
.B1(n_109),
.B2(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_65),
.B1(n_59),
.B2(n_67),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_108),
.B(n_110),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_68),
.B1(n_69),
.B2(n_83),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_83),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_47),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_13),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_86),
.B(n_20),
.C(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_5),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_123),
.B1(n_36),
.B2(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_14),
.B1(n_45),
.B2(n_19),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_29),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_14),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_16),
.B1(n_25),
.B2(n_30),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_13),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_140),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_131),
.B(n_129),
.C(n_133),
.D(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_126),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_147),
.C(n_120),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_31),
.B(n_33),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_124),
.B(n_134),
.C(n_125),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_152),
.C(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_139),
.B(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_138),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_150),
.B1(n_149),
.B2(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_143),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_151),
.C(n_157),
.Y(n_163)
);


endmodule