module fake_ariane_2149_n_2770 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2770);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2770;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2662;
wire n_1259;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_727;
wire n_699;
wire n_2075;
wire n_1726;
wire n_590;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_545;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_640;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_649;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_586;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_2647;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_1968;
wire n_918;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_820;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_969;
wire n_2028;
wire n_1663;
wire n_919;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_1720;
wire n_663;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_2212;
wire n_761;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1806;
wire n_1533;
wire n_671;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_1474;
wire n_2081;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_803;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_333),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_390),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_105),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_98),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_363),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_77),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_364),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_301),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_185),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_176),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_240),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_490),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_98),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_388),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_314),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_499),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_392),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_246),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_299),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_457),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_410),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_524),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_363),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_206),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_246),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_407),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_519),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_227),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_451),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_476),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_404),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_403),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_298),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_78),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_387),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_279),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_72),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_329),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_222),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_447),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_430),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_391),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_518),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_238),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_527),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_69),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_494),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_195),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_107),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_220),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_508),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_426),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_503),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_137),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_415),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_485),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_338),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_487),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_107),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_486),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_269),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_211),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_42),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_90),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_129),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_509),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_496),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_233),
.Y(n_606)
);

BUFx5_ASAP7_75t_L g607 ( 
.A(n_139),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_86),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_28),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_330),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_358),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_231),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_223),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_505),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_429),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_336),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_386),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_437),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_70),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_406),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_319),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_445),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_421),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_338),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_368),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_341),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_169),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_419),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_401),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_381),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_214),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_72),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_13),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_216),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_492),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_149),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_475),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_459),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_378),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_8),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_399),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_153),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_4),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_229),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_192),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_166),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_84),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_177),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_121),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_477),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_10),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_44),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_242),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_145),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_89),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_78),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_469),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_303),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_69),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_264),
.Y(n_662)
);

BUFx5_ASAP7_75t_L g663 ( 
.A(n_428),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_131),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_237),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_22),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_83),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_431),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_454),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_179),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_257),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_204),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_215),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_247),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

CKINVDCx14_ASAP7_75t_R g676 ( 
.A(n_121),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_56),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_77),
.Y(n_678)
);

BUFx5_ASAP7_75t_L g679 ( 
.A(n_265),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_89),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_389),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_438),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_52),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_136),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_34),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_309),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_167),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_335),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_320),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_434),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_0),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_177),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_235),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_423),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_156),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_308),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_33),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_215),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_464),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_317),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_144),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_506),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_45),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_52),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_59),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_218),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_396),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_452),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_374),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_319),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_328),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_424),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_307),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_71),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_465),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_372),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_263),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_495),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_456),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_258),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_308),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_224),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_29),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_332),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_479),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_383),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_317),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_60),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_207),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_478),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_153),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_17),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_234),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_483),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_39),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_432),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_141),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_500),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_122),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_420),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_279),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_37),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_412),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_409),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_336),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_513),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_346),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_288),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_23),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_525),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_144),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_425),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_74),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_191),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_474),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_236),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_214),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_1),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_507),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_470),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_446),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_201),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_112),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_247),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_297),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_229),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_448),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_209),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_71),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_230),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_39),
.Y(n_772)
);

CKINVDCx14_ASAP7_75t_R g773 ( 
.A(n_473),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_160),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_28),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_481),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_329),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_161),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_271),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_510),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_193),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_161),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_439),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_228),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_472),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_44),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_13),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_123),
.Y(n_788)
);

BUFx2_ASAP7_75t_SL g789 ( 
.A(n_461),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_480),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_263),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_440),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_463),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_436),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_123),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_255),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_100),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_284),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_211),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_414),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_29),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_332),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_294),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_417),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_427),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_45),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_408),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_295),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_405),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_383),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_258),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_367),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_398),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_491),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_6),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_66),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_166),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_26),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_366),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_143),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_493),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_130),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_262),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_318),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_250),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_160),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_42),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_325),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_344),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_195),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_369),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_93),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_411),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_30),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_523),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_170),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_146),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_112),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_12),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_75),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_218),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_86),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_394),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_148),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_441),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_341),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_416),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_450),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_462),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_88),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_393),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_364),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_489),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_289),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_276),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_362),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_198),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_163),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_471),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_488),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_1),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_129),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_455),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_512),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_349),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_32),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_118),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_442),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_94),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_520),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_402),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_68),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_453),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_178),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_307),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_502),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_422),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_119),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_435),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_122),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_35),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_444),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_296),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_413),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_515),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_235),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_516),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_273),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_326),
.Y(n_889)
);

CKINVDCx14_ASAP7_75t_R g890 ( 
.A(n_382),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_131),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_243),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_221),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_369),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_498),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_397),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_270),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_400),
.Y(n_898)
);

CKINVDCx14_ASAP7_75t_R g899 ( 
.A(n_356),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_55),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_68),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_191),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_257),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_208),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_384),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_312),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_193),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_283),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_347),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_517),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_379),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_224),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_282),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_497),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_74),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_528),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_351),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_183),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_482),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_222),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_315),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_342),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_271),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_276),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_178),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_377),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_204),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_262),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_128),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_466),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_449),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_282),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_511),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_325),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_24),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_179),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_187),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_82),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_468),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_504),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_14),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_348),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_281),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_365),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_175),
.Y(n_945)
);

BUFx10_ASAP7_75t_L g946 ( 
.A(n_186),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_49),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_360),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_385),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_199),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_333),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_165),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_395),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_142),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_484),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_458),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_635),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_635),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_635),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_826),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_826),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_659),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_676),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_826),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_842),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_842),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_641),
.Y(n_968)
);

CKINVDCx14_ASAP7_75t_R g969 ( 
.A(n_890),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_641),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_899),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_842),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_667),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_536),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_680),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_680),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_696),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_696),
.Y(n_978)
);

INVxp33_ASAP7_75t_L g979 ( 
.A(n_585),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_766),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_667),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_655),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_718),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_607),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_549),
.Y(n_985)
);

INVxp33_ASAP7_75t_SL g986 ( 
.A(n_572),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_718),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_561),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_754),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_674),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_754),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_786),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_786),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_837),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_837),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_674),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_846),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_724),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_578),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_648),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_694),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_629),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_854),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_607),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_607),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_724),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_607),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_607),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_729),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_549),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_629),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_847),
.Y(n_1014)
);

INVxp33_ASAP7_75t_SL g1015 ( 
.A(n_681),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_558),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_607),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_659),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_648),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_729),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_742),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_847),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_660),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_742),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_607),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_679),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_558),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_679),
.Y(n_1028)
);

CKINVDCx16_ASAP7_75t_R g1029 ( 
.A(n_538),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_679),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_679),
.Y(n_1031)
);

OAI22x1_ASAP7_75t_R g1032 ( 
.A1(n_968),
.A2(n_839),
.B1(n_904),
.B2(n_806),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_984),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_984),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_964),
.B(n_594),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_982),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_974),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_985),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_963),
.B(n_660),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_963),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_985),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1026),
.Y(n_1042)
);

BUFx8_ASAP7_75t_L g1043 ( 
.A(n_1018),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1026),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_1004),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_974),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_974),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_974),
.Y(n_1048)
);

OA21x2_ASAP7_75t_L g1049 ( 
.A1(n_1006),
.A2(n_550),
.B(n_541),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1007),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_985),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_1002),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1009),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_986),
.A2(n_839),
.B1(n_904),
.B2(n_806),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1010),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_986),
.B(n_813),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_958),
.B(n_773),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1017),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1015),
.A2(n_929),
.B1(n_938),
.B2(n_920),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_957),
.B(n_885),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1025),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1028),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1030),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_959),
.B(n_625),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1031),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_960),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_961),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_965),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1018),
.B(n_672),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_966),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1012),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_967),
.B(n_679),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_972),
.B(n_625),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_987),
.B(n_679),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_975),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_976),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_977),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_978),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_983),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_991),
.B(n_679),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_989),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_R g1082 ( 
.A1(n_968),
.A2(n_929),
.B1(n_938),
.B2(n_920),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_995),
.B(n_631),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_992),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_980),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_997),
.B(n_672),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_993),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_994),
.B(n_851),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1001),
.B(n_953),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1003),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_969),
.B(n_538),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1005),
.B(n_551),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_999),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1045),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_1043),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1040),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_1032),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1043),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_1056),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1079),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1085),
.B(n_979),
.Y(n_1101)
);

BUFx10_ASAP7_75t_L g1102 ( 
.A(n_1086),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1085),
.B(n_1029),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1076),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1043),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1043),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_1032),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_1093),
.B(n_988),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1076),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1054),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1081),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1054),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1059),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1059),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1081),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1075),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1075),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1036),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1082),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1036),
.B(n_988),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_R g1121 ( 
.A(n_1093),
.B(n_1004),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1052),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_1093),
.B(n_1013),
.Y(n_1123)
);

XOR2xp5_ASAP7_75t_L g1124 ( 
.A(n_1052),
.B(n_1013),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1093),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_1040),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1075),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1091),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1033),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1040),
.Y(n_1130)
);

NAND2xp33_ASAP7_75t_R g1131 ( 
.A(n_1091),
.B(n_1014),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1079),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1079),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1079),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1057),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1078),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1079),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1078),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_1082),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1033),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1035),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_1077),
.B(n_1000),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1057),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1078),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1057),
.Y(n_1145)
);

OR2x2_ASAP7_75t_SL g1146 ( 
.A(n_1088),
.B(n_962),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1087),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1079),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1087),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1033),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1084),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1135),
.B(n_1083),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1104),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_1135),
.B(n_1084),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1129),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1125),
.B(n_1071),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1094),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1101),
.B(n_996),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1125),
.B(n_1086),
.Y(n_1159)
);

CKINVDCx8_ASAP7_75t_R g1160 ( 
.A(n_1097),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1096),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1121),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1102),
.B(n_1086),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1109),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1129),
.B(n_1060),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1126),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1140),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1111),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1143),
.B(n_1071),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1140),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1150),
.Y(n_1171)
);

AND2x6_ASAP7_75t_L g1172 ( 
.A(n_1150),
.B(n_1060),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1130),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1110),
.A2(n_1015),
.B1(n_1086),
.B2(n_1049),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1103),
.B(n_998),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1128),
.B(n_1083),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1102),
.B(n_1060),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1112),
.A2(n_1049),
.B1(n_942),
.B2(n_1083),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1118),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1116),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1143),
.A2(n_942),
.B1(n_1022),
.B2(n_1014),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1142),
.B(n_1039),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1096),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1117),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1115),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1145),
.A2(n_896),
.B1(n_933),
.B2(n_898),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1102),
.B(n_1053),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1100),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1120),
.B(n_1008),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1100),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1127),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1136),
.Y(n_1192)
);

AND2x6_ASAP7_75t_L g1193 ( 
.A(n_1138),
.B(n_1039),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1122),
.B(n_1022),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1145),
.B(n_1016),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1098),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1123),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1144),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1147),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1100),
.Y(n_1200)
);

AND2x6_ASAP7_75t_L g1201 ( 
.A(n_1149),
.B(n_1100),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1132),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1098),
.B(n_1039),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1099),
.B(n_1074),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1133),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1124),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1134),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1108),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1137),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1095),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1105),
.B(n_1039),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1106),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1148),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_SL g1214 ( 
.A(n_1141),
.B(n_563),
.C(n_560),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1131),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1151),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1099),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1099),
.B(n_1074),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1141),
.B(n_1080),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1146),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1113),
.B(n_1069),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1114),
.Y(n_1222)
);

BUFx4f_ASAP7_75t_L g1223 ( 
.A(n_1139),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1107),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1107),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1119),
.B(n_1080),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1119),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1100),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1104),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1153),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1186),
.B(n_970),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1164),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1168),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1155),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1173),
.B(n_1064),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1204),
.B(n_1053),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1155),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1158),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1167),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1189),
.B(n_1027),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1216),
.B(n_896),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1157),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1183),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1185),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1229),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1191),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1192),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1198),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1199),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1216),
.B(n_1084),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1222),
.A2(n_973),
.B1(n_981),
.B2(n_970),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1204),
.B(n_1058),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1218),
.B(n_898),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1167),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_L g1255 ( 
.A(n_1201),
.B(n_1058),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1190),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1170),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1190),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1175),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1173),
.B(n_1064),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1169),
.Y(n_1261)
);

AO22x2_ASAP7_75t_L g1262 ( 
.A1(n_1222),
.A2(n_981),
.B1(n_990),
.B2(n_973),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1157),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1195),
.B(n_999),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1162),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1180),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1176),
.B(n_1221),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1170),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1209),
.B(n_1084),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1184),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1197),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1194),
.B(n_990),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1184),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_L g1274 ( 
.A(n_1201),
.B(n_1061),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1152),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1176),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1209),
.B(n_1084),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1171),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1221),
.B(n_1069),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1152),
.Y(n_1280)
);

AO22x2_ASAP7_75t_L g1281 ( 
.A1(n_1178),
.A2(n_1020),
.B1(n_1021),
.B2(n_1011),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1179),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1159),
.B(n_933),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1166),
.B(n_956),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1171),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1154),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1166),
.B(n_956),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1219),
.B(n_1061),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1219),
.B(n_1011),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1154),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1160),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1200),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1169),
.A2(n_1069),
.B1(n_971),
.B2(n_964),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1215),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1163),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1225),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1226),
.B(n_1203),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1174),
.B(n_1062),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1223),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1203),
.B(n_1064),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1196),
.B(n_1073),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1223),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1182),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1211),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1182),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1174),
.B(n_1062),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1165),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1178),
.A2(n_1020),
.B1(n_1024),
.B2(n_1021),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1165),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1211),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1165),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1208),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1165),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1196),
.B(n_1069),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1220),
.A2(n_1024),
.B1(n_1049),
.B2(n_971),
.Y(n_1316)
);

NAND2x1_ASAP7_75t_L g1317 ( 
.A(n_1201),
.B(n_1050),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1183),
.B(n_1084),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1156),
.B(n_1063),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1156),
.A2(n_1077),
.B(n_1065),
.C(n_1063),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1206),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1206),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1172),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1210),
.B(n_1019),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1187),
.B(n_1077),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1177),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1172),
.Y(n_1327)
);

AO22x2_ASAP7_75t_L g1328 ( 
.A1(n_1214),
.A2(n_1088),
.B1(n_656),
.B2(n_693),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1172),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1225),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1172),
.B(n_1065),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1077),
.B1(n_552),
.B2(n_714),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1264),
.B(n_1224),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1261),
.A2(n_1181),
.B(n_1214),
.C(n_1217),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1256),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1261),
.B(n_1172),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_R g1337 ( 
.A(n_1265),
.B(n_1210),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1236),
.A2(n_1161),
.B(n_1188),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1236),
.A2(n_1161),
.B(n_1188),
.Y(n_1339)
);

AND2x2_ASAP7_75t_SL g1340 ( 
.A(n_1231),
.B(n_1227),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1234),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1289),
.B(n_1212),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1326),
.B(n_1207),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1252),
.A2(n_1187),
.B(n_1200),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1230),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1252),
.A2(n_1228),
.B(n_1190),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1272),
.B(n_1181),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1319),
.A2(n_559),
.B(n_1023),
.C(n_1202),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1281),
.A2(n_1225),
.B1(n_1212),
.B2(n_1213),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1319),
.A2(n_1228),
.B(n_1190),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1256),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1237),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1263),
.B(n_1242),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1288),
.A2(n_1228),
.B(n_1213),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1326),
.B(n_1207),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1276),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1288),
.A2(n_1205),
.B(n_717),
.C(n_721),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1239),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1255),
.A2(n_1228),
.B(n_1055),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1295),
.A2(n_563),
.B1(n_569),
.B2(n_560),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1238),
.B(n_1193),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1295),
.A2(n_574),
.B1(n_575),
.B2(n_569),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1267),
.B(n_1073),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1238),
.B(n_1259),
.Y(n_1364)
);

NOR3xp33_ASAP7_75t_L g1365 ( 
.A(n_1284),
.B(n_1287),
.C(n_1324),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1320),
.B(n_1055),
.C(n_1050),
.Y(n_1366)
);

AOI221xp5_ASAP7_75t_L g1367 ( 
.A1(n_1281),
.A2(n_819),
.B1(n_932),
.B2(n_769),
.C(n_712),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1274),
.A2(n_1055),
.B(n_1050),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1297),
.A2(n_1193),
.B1(n_1201),
.B2(n_936),
.Y(n_1370)
);

AND2x6_ASAP7_75t_L g1371 ( 
.A(n_1307),
.B(n_1193),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1294),
.B(n_1068),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1254),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_SL g1374 ( 
.A1(n_1317),
.A2(n_1072),
.B(n_853),
.C(n_703),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_L g1375 ( 
.A(n_1271),
.B(n_1201),
.Y(n_1375)
);

AND2x6_ASAP7_75t_SL g1376 ( 
.A(n_1235),
.B(n_1072),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1330),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1232),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1275),
.B(n_1073),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1280),
.B(n_1087),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1300),
.B(n_1090),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1331),
.A2(n_1042),
.B(n_1034),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1233),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1282),
.B(n_1068),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1331),
.A2(n_1042),
.B(n_1034),
.Y(n_1385)
);

AO32x2_ASAP7_75t_L g1386 ( 
.A1(n_1251),
.A2(n_853),
.A3(n_703),
.B1(n_1049),
.B2(n_1089),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1332),
.A2(n_1067),
.B(n_1070),
.C(n_1066),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1298),
.A2(n_1049),
.B(n_1042),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1299),
.B(n_594),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1303),
.B(n_1090),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1256),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1253),
.A2(n_533),
.B1(n_535),
.B2(n_531),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1312),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1300),
.B(n_1090),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1279),
.B(n_1066),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1291),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1309),
.A2(n_1067),
.B(n_1070),
.C(n_1066),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1240),
.B(n_1304),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1243),
.A2(n_1044),
.B(n_1034),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1235),
.B(n_1067),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1325),
.A2(n_1044),
.B(n_1070),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1311),
.A2(n_1092),
.B(n_1089),
.C(n_556),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1260),
.B(n_1068),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1318),
.A2(n_1044),
.B(n_1046),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1260),
.B(n_1092),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1243),
.A2(n_554),
.B(n_542),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1257),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1301),
.B(n_1068),
.Y(n_1408)
);

CKINVDCx10_ASAP7_75t_R g1409 ( 
.A(n_1302),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1301),
.B(n_1068),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1292),
.A2(n_554),
.B(n_542),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1283),
.A2(n_537),
.B(n_540),
.C(n_534),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1318),
.A2(n_739),
.B(n_708),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1244),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1310),
.B(n_538),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1245),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1305),
.B(n_1068),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1246),
.A2(n_739),
.B(n_708),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1315),
.B(n_595),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1258),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1241),
.A2(n_547),
.B1(n_553),
.B2(n_544),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1247),
.A2(n_835),
.B(n_807),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1248),
.A2(n_835),
.B(n_807),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1293),
.B(n_573),
.C(n_549),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1249),
.B(n_1038),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1308),
.B(n_595),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1325),
.A2(n_545),
.B(n_568),
.C(n_543),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1296),
.B(n_539),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1322),
.B(n_574),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1313),
.A2(n_562),
.B(n_566),
.C(n_555),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1347),
.B(n_1321),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1398),
.B(n_1316),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1340),
.B(n_1258),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1338),
.A2(n_1258),
.B(n_1298),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_R g1435 ( 
.A(n_1409),
.B(n_1312),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1367),
.A2(n_1262),
.B1(n_1328),
.B2(n_1266),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1351),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1363),
.B(n_1328),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1345),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1336),
.A2(n_1269),
.B1(n_1277),
.B2(n_1306),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1328),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1337),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1339),
.A2(n_1306),
.B(n_1277),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1351),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1334),
.A2(n_571),
.B(n_584),
.C(n_582),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1342),
.B(n_1270),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_SL g1447 ( 
.A(n_1348),
.B(n_580),
.C(n_575),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1333),
.B(n_1273),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1419),
.B(n_1262),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1364),
.B(n_1285),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_R g1451 ( 
.A(n_1396),
.B(n_1393),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1370),
.A2(n_1269),
.B1(n_1250),
.B2(n_1314),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1356),
.B(n_1268),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1377),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1388),
.A2(n_1250),
.B(n_1278),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1357),
.A2(n_1327),
.B(n_1329),
.C(n_1323),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1429),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1343),
.A2(n_1286),
.B1(n_1290),
.B2(n_894),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1351),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1360),
.A2(n_603),
.B(n_608),
.C(n_588),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1424),
.A2(n_877),
.B(n_579),
.C(n_586),
.Y(n_1461)
);

NOR2xp67_ASAP7_75t_L g1462 ( 
.A(n_1355),
.B(n_1038),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1365),
.B(n_580),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_L g1464 ( 
.A1(n_1372),
.A2(n_1354),
.B(n_1350),
.C(n_1346),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1426),
.B(n_592),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1349),
.A2(n_597),
.B1(n_599),
.B2(n_592),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1335),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1378),
.B(n_597),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1424),
.A2(n_877),
.B(n_593),
.C(n_596),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1344),
.A2(n_587),
.B(n_949),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1359),
.A2(n_587),
.B(n_949),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1375),
.A2(n_587),
.B(n_570),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_SL g1473 ( 
.A(n_1353),
.B(n_1361),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1369),
.A2(n_615),
.B(n_614),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1383),
.B(n_599),
.Y(n_1475)
);

OA22x2_ASAP7_75t_L g1476 ( 
.A1(n_1421),
.A2(n_1392),
.B1(n_1416),
.B2(n_1414),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1341),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1427),
.A2(n_621),
.B(n_623),
.C(n_619),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1374),
.A2(n_675),
.B(n_645),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1368),
.A2(n_881),
.B1(n_891),
.B2(n_872),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_R g1481 ( 
.A(n_1415),
.B(n_539),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1428),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1401),
.A2(n_713),
.B(n_682),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1400),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1352),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1358),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1401),
.A2(n_720),
.B(n_719),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1366),
.A2(n_768),
.B(n_756),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1373),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1407),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1389),
.B(n_1335),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1389),
.B(n_600),
.Y(n_1492)
);

OA22x2_ASAP7_75t_L g1493 ( 
.A1(n_1379),
.A2(n_764),
.B1(n_872),
.B2(n_600),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1390),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_R g1495 ( 
.A(n_1390),
.B(n_557),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1391),
.B(n_564),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1366),
.A2(n_792),
.B(n_780),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1381),
.B(n_764),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1394),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1391),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1399),
.A2(n_809),
.B(n_804),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1362),
.A2(n_951),
.B1(n_950),
.B2(n_883),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1382),
.A2(n_833),
.B(n_821),
.Y(n_1503)
);

AO32x2_ASAP7_75t_L g1504 ( 
.A1(n_1386),
.A2(n_595),
.A3(n_775),
.B1(n_725),
.B2(n_722),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1385),
.A2(n_863),
.B(n_843),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_SL g1506 ( 
.A(n_1371),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1395),
.B(n_881),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1408),
.A2(n_886),
.B1(n_888),
.B2(n_883),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1420),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1376),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1380),
.Y(n_1511)
);

AOI222xp33_ASAP7_75t_L g1512 ( 
.A1(n_1403),
.A2(n_908),
.B1(n_725),
.B2(n_946),
.C1(n_775),
.C2(n_722),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1376),
.B(n_886),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1420),
.B(n_564),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1410),
.B(n_888),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1412),
.B(n_889),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1425),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1417),
.B(n_565),
.Y(n_1518)
);

AND2x6_ASAP7_75t_L g1519 ( 
.A(n_1371),
.B(n_873),
.Y(n_1519)
);

NOR3xp33_ASAP7_75t_SL g1520 ( 
.A(n_1384),
.B(n_891),
.C(n_889),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1418),
.B(n_892),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1402),
.A2(n_613),
.B(n_617),
.C(n_612),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_SL g1523 ( 
.A1(n_1413),
.A2(n_627),
.B(n_634),
.C(n_626),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1430),
.B(n_565),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_SL g1525 ( 
.A(n_1406),
.B(n_892),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1371),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1422),
.B(n_894),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1397),
.A2(n_882),
.B(n_876),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1371),
.B(n_1038),
.Y(n_1529)
);

OR2x6_ASAP7_75t_L g1530 ( 
.A(n_1423),
.B(n_1411),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1386),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1386),
.Y(n_1532)
);

BUFx4_ASAP7_75t_SL g1533 ( 
.A(n_1482),
.Y(n_1533)
);

BUFx4_ASAP7_75t_SL g1534 ( 
.A(n_1454),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1476),
.A2(n_725),
.B1(n_775),
.B2(n_722),
.Y(n_1535)
);

BUFx12f_ASAP7_75t_L g1536 ( 
.A(n_1457),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1437),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1457),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1439),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1526),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1455),
.Y(n_1541)
);

CKINVDCx6p67_ASAP7_75t_R g1542 ( 
.A(n_1459),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1442),
.Y(n_1543)
);

BUFx5_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1437),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1435),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1485),
.Y(n_1547)
);

INVx8_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_SL g1549 ( 
.A(n_1467),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1509),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1431),
.B(n_908),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1510),
.A2(n_1481),
.B1(n_1484),
.B2(n_1495),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1448),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1451),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1446),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1450),
.B(n_637),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1477),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1437),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1444),
.Y(n_1559)
);

INVx5_ASAP7_75t_L g1560 ( 
.A(n_1526),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1499),
.B(n_643),
.Y(n_1561)
);

CKINVDCx16_ASAP7_75t_R g1562 ( 
.A(n_1466),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1526),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1444),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1433),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1453),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1494),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1500),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1532),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1489),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1500),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1432),
.B(n_646),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1529),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1486),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1491),
.Y(n_1575)
);

NAND2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1473),
.B(n_1404),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1490),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1517),
.Y(n_1578)
);

INVx5_ASAP7_75t_L g1579 ( 
.A(n_1519),
.Y(n_1579)
);

BUFx2_ASAP7_75t_SL g1580 ( 
.A(n_1519),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1529),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1519),
.B(n_1387),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1511),
.B(n_1462),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1530),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1493),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1530),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1447),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1436),
.A2(n_946),
.B1(n_908),
.B2(n_631),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1438),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1449),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1441),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1456),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1531),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1464),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1468),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1521),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1513),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1498),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1520),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1492),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1504),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1525),
.B(n_1038),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1475),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1463),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1496),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1515),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1480),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1452),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1507),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1514),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1465),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1516),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1504),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1504),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_R g1615 ( 
.A(n_1546),
.B(n_897),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1594),
.A2(n_1470),
.B(n_1434),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1536),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1594),
.A2(n_1443),
.B(n_1471),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1592),
.A2(n_1527),
.B1(n_1458),
.B2(n_946),
.Y(n_1619)
);

OAI22x1_ASAP7_75t_L g1620 ( 
.A1(n_1552),
.A2(n_1604),
.B1(n_1555),
.B2(n_1611),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1550),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1551),
.A2(n_1445),
.B(n_1478),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1539),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1578),
.B(n_1440),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1593),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1553),
.B(n_1483),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1576),
.A2(n_1584),
.B(n_1583),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1612),
.A2(n_1487),
.B(n_1488),
.Y(n_1628)
);

INVx8_ASAP7_75t_L g1629 ( 
.A(n_1548),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1601),
.A2(n_1479),
.B(n_1497),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1578),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1472),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1613),
.A2(n_1505),
.B(n_1503),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1575),
.B(n_1512),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1547),
.Y(n_1635)
);

OAI211xp5_ASAP7_75t_L g1636 ( 
.A1(n_1607),
.A2(n_1502),
.B(n_1460),
.C(n_926),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1536),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1571),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1576),
.A2(n_1474),
.B(n_1528),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1568),
.A2(n_1522),
.B(n_1501),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1584),
.A2(n_1524),
.B(n_1518),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1550),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1583),
.A2(n_1047),
.B(n_1046),
.Y(n_1643)
);

NOR2x1p5_ASAP7_75t_L g1644 ( 
.A(n_1538),
.B(n_895),
.Y(n_1644)
);

AOI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1535),
.A2(n_1523),
.B(n_1469),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1607),
.A2(n_1608),
.B1(n_1535),
.B2(n_1588),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1538),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_SL g1648 ( 
.A1(n_1554),
.A2(n_653),
.B(n_664),
.C(n_647),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1649)
);

AO31x2_ASAP7_75t_L g1650 ( 
.A1(n_1613),
.A2(n_1461),
.A3(n_1508),
.B(n_910),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1608),
.A2(n_926),
.B1(n_950),
.B2(n_897),
.Y(n_1651)
);

CKINVDCx6p67_ASAP7_75t_R g1652 ( 
.A(n_1554),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1570),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1566),
.B(n_677),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1589),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1541),
.A2(n_1047),
.B(n_1046),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1562),
.B(n_951),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1586),
.B(n_789),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1557),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1545),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1565),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1541),
.A2(n_1048),
.B(n_1047),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_SL g1663 ( 
.A1(n_1608),
.A2(n_765),
.B(n_763),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1612),
.A2(n_1048),
.B(n_1051),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1603),
.B(n_678),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1609),
.B(n_685),
.Y(n_1666)
);

AO31x2_ASAP7_75t_L g1667 ( 
.A1(n_1614),
.A2(n_916),
.A3(n_931),
.B(n_905),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1564),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1593),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1577),
.Y(n_1670)
);

AO221x1_ASAP7_75t_L g1671 ( 
.A1(n_1596),
.A2(n_573),
.B1(n_810),
.B2(n_549),
.C(n_690),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1586),
.B(n_848),
.Y(n_1672)
);

NAND2x1_ASAP7_75t_L g1673 ( 
.A(n_1537),
.B(n_1051),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1569),
.A2(n_1048),
.B(n_939),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1646),
.A2(n_1596),
.B1(n_1572),
.B2(n_1603),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1618),
.A2(n_1569),
.B(n_1537),
.Y(n_1676)
);

BUFx8_ASAP7_75t_SL g1677 ( 
.A(n_1617),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1627),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1635),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1646),
.A2(n_1580),
.B1(n_1544),
.B2(n_1579),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1653),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1625),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1631),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1619),
.A2(n_1597),
.B1(n_1585),
.B2(n_1591),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1625),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1622),
.A2(n_1579),
.B1(n_1597),
.B2(n_1609),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1623),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1659),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1670),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1624),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1624),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1669),
.Y(n_1693)
);

INVx8_ASAP7_75t_L g1694 ( 
.A(n_1629),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

INVx6_ASAP7_75t_L g1696 ( 
.A(n_1629),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1667),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1652),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1616),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1616),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1674),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1674),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1638),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1642),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1660),
.B(n_1591),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1630),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1630),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1633),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1619),
.A2(n_1598),
.B1(n_1606),
.B2(n_1611),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1633),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1649),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1656),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1649),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1634),
.A2(n_1598),
.B1(n_1606),
.B2(n_1588),
.Y(n_1719)
);

INVxp33_ASAP7_75t_L g1720 ( 
.A(n_1615),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1661),
.B(n_1595),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1666),
.B(n_1556),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1651),
.A2(n_1600),
.B1(n_1587),
.B2(n_1599),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1690),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1637),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1690),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1679),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1705),
.B(n_1626),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1705),
.B(n_1654),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1686),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1714),
.A2(n_1651),
.B1(n_1622),
.B2(n_1636),
.Y(n_1732)
);

BUFx5_ASAP7_75t_L g1733 ( 
.A(n_1710),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1699),
.B(n_1587),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1675),
.A2(n_1620),
.B1(n_1671),
.B2(n_1600),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1677),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_R g1738 ( 
.A(n_1694),
.B(n_1629),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1680),
.B(n_1658),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1694),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1679),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1682),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1684),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1685),
.A2(n_1636),
.B1(n_1628),
.B2(n_1657),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1680),
.B(n_1647),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1675),
.A2(n_1644),
.B1(n_1645),
.B2(n_1665),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1691),
.B(n_1632),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1682),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1692),
.B(n_1632),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1560),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1687),
.B(n_1668),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1723),
.A2(n_1548),
.B(n_1610),
.C(n_1645),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1708),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1697),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1692),
.B(n_1658),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1709),
.B(n_1668),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1684),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1688),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1695),
.B(n_1628),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1711),
.B(n_1543),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1689),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_R g1764 ( 
.A(n_1722),
.B(n_1672),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1719),
.A2(n_1582),
.B1(n_1579),
.B2(n_1672),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1706),
.B(n_1543),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1693),
.B(n_1683),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1721),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1688),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1681),
.A2(n_1640),
.B(n_1639),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1706),
.Y(n_1771)
);

AOI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1716),
.A2(n_1648),
.B1(n_1582),
.B2(n_1672),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1698),
.A2(n_1574),
.B1(n_1582),
.B2(n_1704),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1693),
.B(n_1650),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1683),
.Y(n_1775)
);

CKINVDCx16_ASAP7_75t_R g1776 ( 
.A(n_1716),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1771),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1734),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1771),
.B(n_1678),
.Y(n_1781)
);

NAND2x1_ASAP7_75t_L g1782 ( 
.A(n_1740),
.B(n_1696),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1776),
.B(n_1718),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1724),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1727),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1761),
.B(n_1718),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1744),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1725),
.Y(n_1789)
);

OA21x2_ASAP7_75t_L g1790 ( 
.A1(n_1761),
.A2(n_1712),
.B(n_1774),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1775),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1676),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1729),
.B(n_1712),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1751),
.B(n_1678),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1767),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1751),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1728),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1748),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1742),
.B(n_1678),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1726),
.B(n_1676),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1740),
.B(n_1678),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1749),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1774),
.B(n_1698),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1746),
.B(n_1756),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1730),
.B(n_1704),
.Y(n_1807)
);

AOI33xp33_ASAP7_75t_L g1808 ( 
.A1(n_1747),
.A2(n_831),
.A3(n_765),
.B1(n_838),
.B2(n_828),
.B3(n_763),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1791),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1796),
.B(n_1769),
.Y(n_1810)
);

OAI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1787),
.A2(n_1736),
.B1(n_1745),
.B2(n_1732),
.C(n_1754),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1779),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1779),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1792),
.B(n_1800),
.Y(n_1814)
);

AOI211x1_ASAP7_75t_L g1815 ( 
.A1(n_1792),
.A2(n_1732),
.B(n_1745),
.C(n_1753),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1790),
.B(n_1757),
.C(n_1770),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1801),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1795),
.Y(n_1818)
);

AND2x4_ASAP7_75t_SL g1819 ( 
.A(n_1806),
.B(n_1758),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1800),
.B(n_1758),
.Y(n_1820)
);

INVx4_ASAP7_75t_SL g1821 ( 
.A(n_1803),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1797),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1797),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1806),
.B(n_1737),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1804),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1766),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1804),
.Y(n_1828)
);

INVx5_ASAP7_75t_L g1829 ( 
.A(n_1781),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_SL g1830 ( 
.A(n_1783),
.B(n_1750),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1778),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1803),
.A2(n_1765),
.B1(n_1707),
.B2(n_1704),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1788),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1784),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1784),
.Y(n_1835)
);

AO21x1_ASAP7_75t_L g1836 ( 
.A1(n_1799),
.A2(n_1765),
.B(n_1772),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1777),
.B(n_1768),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1798),
.A2(n_1764),
.B1(n_1750),
.B2(n_1773),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1811),
.A2(n_702),
.B1(n_705),
.B2(n_692),
.C(n_688),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1809),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1820),
.B(n_1777),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1822),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1824),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1818),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1820),
.B(n_1777),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1826),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1815),
.B(n_1790),
.C(n_1794),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1817),
.B(n_1790),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1828),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1836),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_L g1851 ( 
.A(n_1816),
.B(n_1790),
.C(n_1780),
.Y(n_1851)
);

NAND4xp25_ASAP7_75t_L g1852 ( 
.A(n_1817),
.B(n_1780),
.C(n_1808),
.D(n_1777),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1827),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1810),
.B(n_1805),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1834),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1835),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1827),
.B(n_1781),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1812),
.A2(n_1823),
.B(n_1813),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1814),
.B(n_1781),
.Y(n_1860)
);

AO21x2_ASAP7_75t_L g1861 ( 
.A1(n_1836),
.A2(n_1785),
.B(n_1805),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1830),
.A2(n_1782),
.B(n_1750),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1812),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1783),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1837),
.Y(n_1865)
);

INVx4_ASAP7_75t_L g1866 ( 
.A(n_1829),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1831),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1837),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1813),
.B(n_1785),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1846),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1854),
.B(n_1760),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1854),
.B(n_1793),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1861),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1865),
.B(n_1819),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1840),
.B(n_1755),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1840),
.B(n_1829),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1865),
.B(n_1829),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1846),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1850),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1851),
.A2(n_1720),
.B(n_710),
.C(n_723),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1855),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_SL g1882 ( 
.A(n_1839),
.B(n_1838),
.C(n_1832),
.D(n_1534),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1855),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1861),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1866),
.B(n_1829),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1864),
.B(n_1829),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1844),
.B(n_1867),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1864),
.B(n_1830),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1853),
.B(n_1793),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1853),
.B(n_1823),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1852),
.B(n_1833),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1868),
.Y(n_1892)
);

OR2x6_ASAP7_75t_L g1893 ( 
.A(n_1862),
.B(n_1548),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1857),
.B(n_1821),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1861),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1857),
.B(n_1825),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1866),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1866),
.B(n_1821),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1842),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1870),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1841),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1892),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1874),
.B(n_1841),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1874),
.B(n_1845),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1888),
.B(n_1845),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1878),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1881),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1879),
.B(n_1856),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1879),
.B(n_1843),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1880),
.B(n_1849),
.Y(n_1911)
);

OR2x6_ASAP7_75t_L g1912 ( 
.A(n_1893),
.B(n_1694),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1877),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1888),
.B(n_1859),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1883),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1899),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1887),
.B(n_1847),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1892),
.B(n_1848),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1891),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1875),
.B(n_1848),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1871),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1873),
.B(n_1869),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1894),
.B(n_1859),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1872),
.B(n_1869),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1890),
.Y(n_1925)
);

O2A1O1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1873),
.A2(n_727),
.B(n_730),
.C(n_707),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1889),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1884),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1884),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1894),
.B(n_1886),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1895),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1895),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1876),
.B(n_1860),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1897),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1886),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1898),
.B(n_1863),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1885),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1898),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1898),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1885),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1893),
.Y(n_1941)
);

OAI21xp33_ASAP7_75t_L g1942 ( 
.A1(n_1893),
.A2(n_1860),
.B(n_1780),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1930),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1939),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1901),
.B(n_1821),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1923),
.B(n_1735),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1939),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1938),
.B(n_1882),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1914),
.B(n_1821),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1920),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1904),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1902),
.B(n_1858),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1929),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1931),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1932),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1913),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1909),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1909),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1921),
.B(n_1858),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1924),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1919),
.B(n_1833),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1910),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1910),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1906),
.B(n_1741),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1911),
.A2(n_1782),
.B(n_831),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1911),
.B(n_750),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1900),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1905),
.B(n_1738),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1935),
.B(n_1741),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1907),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1918),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1934),
.B(n_1696),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1927),
.B(n_740),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1908),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1937),
.B(n_1696),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1937),
.B(n_1696),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1915),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1933),
.B(n_1803),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1922),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1936),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1917),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1941),
.B(n_1803),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1922),
.Y(n_1984)
);

INVx4_ASAP7_75t_L g1985 ( 
.A(n_1912),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1925),
.B(n_752),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1936),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1940),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1916),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1912),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1912),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1942),
.B(n_755),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1926),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1926),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1924),
.B(n_770),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1919),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1902),
.B(n_772),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1939),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1934),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1930),
.B(n_828),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1930),
.B(n_1694),
.Y(n_2001)
);

INVx3_ASAP7_75t_SL g2002 ( 
.A(n_1912),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1928),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1943),
.B(n_774),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1996),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1946),
.B(n_2001),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1944),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1944),
.B(n_782),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1945),
.B(n_1694),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1996),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1950),
.A2(n_866),
.B(n_838),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1945),
.B(n_784),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1998),
.B(n_787),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1969),
.B(n_796),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1998),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_2000),
.B(n_811),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1961),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1982),
.A2(n_1678),
.B1(n_1707),
.B2(n_1605),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1961),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1952),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1985),
.B(n_1549),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_2002),
.B(n_818),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1947),
.B(n_827),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1949),
.B(n_836),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1995),
.Y(n_2025)
);

OAI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1950),
.A2(n_874),
.B(n_866),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1965),
.B(n_850),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1963),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1997),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1974),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1986),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1965),
.B(n_852),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1963),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1982),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1952),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1987),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1952),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1987),
.Y(n_2038)
);

NAND2x1p5_ASAP7_75t_L g2039 ( 
.A(n_1985),
.B(n_1533),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2000),
.B(n_855),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2000),
.B(n_856),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1999),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1972),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1981),
.B(n_867),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1999),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1951),
.B(n_875),
.Y(n_2046)
);

INVx1_ASAP7_75t_SL g2047 ( 
.A(n_2002),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1951),
.B(n_878),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1957),
.B(n_880),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1976),
.Y(n_2050)
);

NAND2x1p5_ASAP7_75t_L g2051 ( 
.A(n_1985),
.B(n_1533),
.Y(n_2051)
);

CKINVDCx16_ASAP7_75t_R g2052 ( 
.A(n_1990),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1972),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1976),
.B(n_1977),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1957),
.B(n_893),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1977),
.B(n_901),
.Y(n_2056)
);

NOR2xp67_ASAP7_75t_L g2057 ( 
.A(n_1988),
.B(n_0),
.Y(n_2057)
);

NOR2xp67_ASAP7_75t_L g2058 ( 
.A(n_1988),
.B(n_2),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1991),
.B(n_902),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1954),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_1958),
.B(n_1959),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1955),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1964),
.B(n_906),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1980),
.B(n_907),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1994),
.A2(n_1678),
.B1(n_1707),
.B2(n_1605),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1956),
.Y(n_2066)
);

BUFx2_ASAP7_75t_L g2067 ( 
.A(n_1973),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1973),
.B(n_912),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1979),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1984),
.B(n_921),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1991),
.B(n_922),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1970),
.B(n_923),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1962),
.B(n_927),
.Y(n_2073)
);

INVxp33_ASAP7_75t_L g2074 ( 
.A(n_1948),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2003),
.Y(n_2075)
);

AND2x2_ASAP7_75t_SL g2076 ( 
.A(n_1948),
.B(n_1534),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1953),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1992),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1967),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1967),
.B(n_928),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1989),
.B(n_934),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1960),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1968),
.B(n_941),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1971),
.B(n_1975),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1983),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1983),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2034),
.A2(n_1966),
.B1(n_1993),
.B2(n_1978),
.Y(n_2087)
);

OAI21xp33_ASAP7_75t_L g2088 ( 
.A1(n_2074),
.A2(n_1983),
.B(n_1993),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2067),
.B(n_943),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2034),
.Y(n_2090)
);

OAI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2054),
.A2(n_900),
.B(n_874),
.Y(n_2091)
);

A2O1A1Ixp33_ASAP7_75t_SL g2092 ( 
.A1(n_2042),
.A2(n_945),
.B(n_918),
.C(n_924),
.Y(n_2092)
);

OAI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_2053),
.A2(n_1752),
.B1(n_1579),
.B2(n_1605),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_2085),
.A2(n_918),
.B(n_900),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2037),
.B(n_924),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2052),
.B(n_952),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2045),
.B(n_2),
.Y(n_2097)
);

AOI21xp33_ASAP7_75t_SL g2098 ( 
.A1(n_2039),
.A2(n_3),
.B(n_5),
.Y(n_2098)
);

A2O1A1Ixp33_ASAP7_75t_L g2099 ( 
.A1(n_2082),
.A2(n_952),
.B(n_602),
.C(n_606),
.Y(n_2099)
);

O2A1O1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_2028),
.A2(n_1561),
.B(n_1663),
.C(n_1602),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2017),
.A2(n_1605),
.B1(n_1549),
.B2(n_1542),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_2076),
.B(n_1733),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2019),
.A2(n_2021),
.B1(n_2047),
.B2(n_2043),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2051),
.B(n_601),
.Y(n_2104)
);

NOR4xp25_ASAP7_75t_L g2105 ( 
.A(n_2028),
.B(n_2033),
.C(n_2005),
.D(n_2010),
.Y(n_2105)
);

OAI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2050),
.A2(n_610),
.B(n_609),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2006),
.B(n_611),
.Y(n_2107)
);

A2O1A1Ixp33_ASAP7_75t_L g2108 ( 
.A1(n_2077),
.A2(n_622),
.B(n_628),
.C(n_620),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2069),
.B(n_632),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2005),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2037),
.B(n_633),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2010),
.Y(n_2112)
);

OAI21xp5_ASAP7_75t_SL g2113 ( 
.A1(n_2020),
.A2(n_573),
.B(n_549),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2007),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2048),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2015),
.Y(n_2116)
);

A2O1A1Ixp33_ASAP7_75t_L g2117 ( 
.A1(n_2057),
.A2(n_640),
.B(n_649),
.C(n_644),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2009),
.B(n_650),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2027),
.B(n_651),
.Y(n_2119)
);

AO22x1_ASAP7_75t_L g2120 ( 
.A1(n_2035),
.A2(n_654),
.B1(n_658),
.B2(n_657),
.Y(n_2120)
);

AOI21xp33_ASAP7_75t_SL g2121 ( 
.A1(n_2086),
.A2(n_3),
.B(n_5),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2068),
.Y(n_2122)
);

AOI31xp33_ASAP7_75t_L g2123 ( 
.A1(n_2061),
.A2(n_662),
.A3(n_665),
.B(n_661),
.Y(n_2123)
);

OAI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2036),
.A2(n_1752),
.B1(n_1807),
.B2(n_1802),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2008),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_2084),
.B(n_1571),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2032),
.B(n_666),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2013),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2013),
.Y(n_2129)
);

INVx2_ASAP7_75t_SL g2130 ( 
.A(n_2024),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2004),
.A2(n_1789),
.B1(n_1807),
.B2(n_670),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_SL g2132 ( 
.A1(n_2084),
.A2(n_671),
.B1(n_684),
.B2(n_673),
.Y(n_2132)
);

NOR3xp33_ASAP7_75t_L g2133 ( 
.A(n_2022),
.B(n_687),
.C(n_686),
.Y(n_2133)
);

OAI33xp33_ASAP7_75t_L g2134 ( 
.A1(n_2060),
.A2(n_699),
.A3(n_697),
.B1(n_701),
.B2(n_698),
.B3(n_689),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2023),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2080),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2014),
.A2(n_704),
.B1(n_711),
.B2(n_706),
.Y(n_2137)
);

NOR3xp33_ASAP7_75t_L g2138 ( 
.A(n_2044),
.B(n_728),
.C(n_715),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2012),
.Y(n_2139)
);

AOI31xp33_ASAP7_75t_L g2140 ( 
.A1(n_2062),
.A2(n_733),
.A3(n_734),
.B(n_732),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2038),
.A2(n_1560),
.B1(n_1564),
.B2(n_1713),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2072),
.B(n_736),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2066),
.B(n_738),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2029),
.A2(n_1733),
.B1(n_743),
.B2(n_746),
.Y(n_2144)
);

OA21x2_ASAP7_75t_L g2145 ( 
.A1(n_2075),
.A2(n_2058),
.B(n_2026),
.Y(n_2145)
);

AOI21xp33_ASAP7_75t_R g2146 ( 
.A1(n_2079),
.A2(n_7),
.B(n_9),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2046),
.A2(n_749),
.B(n_748),
.Y(n_2147)
);

OAI332xp33_ASAP7_75t_L g2148 ( 
.A1(n_2025),
.A2(n_776),
.A3(n_767),
.B1(n_758),
.B2(n_771),
.B3(n_777),
.C1(n_759),
.C2(n_757),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2073),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_2056),
.Y(n_2150)
);

INVx1_ASAP7_75t_SL g2151 ( 
.A(n_2081),
.Y(n_2151)
);

NOR3xp33_ASAP7_75t_L g2152 ( 
.A(n_2071),
.B(n_779),
.C(n_778),
.Y(n_2152)
);

OAI21xp33_ASAP7_75t_SL g2153 ( 
.A1(n_2064),
.A2(n_1641),
.B(n_7),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2055),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2048),
.Y(n_2155)
);

OAI32xp33_ASAP7_75t_L g2156 ( 
.A1(n_2063),
.A2(n_791),
.A3(n_795),
.B1(n_788),
.B2(n_781),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2083),
.B(n_2030),
.Y(n_2157)
);

AOI21xp33_ASAP7_75t_L g2158 ( 
.A1(n_2031),
.A2(n_798),
.B(n_797),
.Y(n_2158)
);

OAI21xp33_ASAP7_75t_L g2159 ( 
.A1(n_2070),
.A2(n_801),
.B(n_799),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_2083),
.Y(n_2160)
);

OAI32xp33_ASAP7_75t_L g2161 ( 
.A1(n_2078),
.A2(n_808),
.A3(n_812),
.B1(n_803),
.B2(n_802),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2049),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2016),
.B(n_9),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2049),
.Y(n_2164)
);

NAND2x1p5_ASAP7_75t_L g2165 ( 
.A(n_2059),
.B(n_1560),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2040),
.Y(n_2166)
);

OA21x2_ASAP7_75t_L g2167 ( 
.A1(n_2011),
.A2(n_816),
.B(n_815),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2041),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2059),
.B(n_817),
.Y(n_2169)
);

OAI21xp33_ASAP7_75t_L g2170 ( 
.A1(n_2065),
.A2(n_822),
.B(n_820),
.Y(n_2170)
);

OAI211xp5_ASAP7_75t_L g2171 ( 
.A1(n_2018),
.A2(n_823),
.B(n_825),
.C(n_824),
.Y(n_2171)
);

OAI21xp33_ASAP7_75t_L g2172 ( 
.A1(n_2074),
.A2(n_830),
.B(n_829),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_2074),
.B(n_832),
.Y(n_2173)
);

O2A1O1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_2074),
.A2(n_840),
.B(n_844),
.C(n_841),
.Y(n_2174)
);

OAI22xp33_ASAP7_75t_L g2175 ( 
.A1(n_2034),
.A2(n_1560),
.B1(n_1715),
.B2(n_1713),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2034),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2034),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2067),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2034),
.Y(n_2179)
);

INVxp67_ASAP7_75t_L g2180 ( 
.A(n_2067),
.Y(n_2180)
);

AOI211xp5_ASAP7_75t_L g2181 ( 
.A1(n_2074),
.A2(n_857),
.B(n_858),
.C(n_834),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2052),
.B(n_861),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_2067),
.Y(n_2183)
);

OAI321xp33_ASAP7_75t_L g2184 ( 
.A1(n_2034),
.A2(n_573),
.A3(n_810),
.B1(n_1563),
.B2(n_1540),
.C(n_1558),
.Y(n_2184)
);

AOI32xp33_ASAP7_75t_L g2185 ( 
.A1(n_2074),
.A2(n_869),
.A3(n_903),
.B1(n_865),
.B2(n_862),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2034),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2074),
.A2(n_911),
.B1(n_913),
.B2(n_909),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2067),
.B(n_10),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2034),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_2067),
.Y(n_2190)
);

INVxp67_ASAP7_75t_L g2191 ( 
.A(n_2067),
.Y(n_2191)
);

OAI21xp5_ASAP7_75t_SL g2192 ( 
.A1(n_2039),
.A2(n_810),
.B(n_573),
.Y(n_2192)
);

OAI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2034),
.A2(n_917),
.B1(n_935),
.B2(n_925),
.C(n_915),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_2067),
.B(n_11),
.Y(n_2194)
);

AOI322xp5_ASAP7_75t_L g2195 ( 
.A1(n_2034),
.A2(n_1715),
.A3(n_947),
.B1(n_948),
.B2(n_937),
.C1(n_944),
.C2(n_1703),
.Y(n_2195)
);

INVx2_ASAP7_75t_SL g2196 ( 
.A(n_2076),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2067),
.B(n_11),
.Y(n_2197)
);

AOI221xp5_ASAP7_75t_L g2198 ( 
.A1(n_2034),
.A2(n_810),
.B1(n_567),
.B2(n_577),
.C(n_576),
.Y(n_2198)
);

OAI31xp33_ASAP7_75t_L g2199 ( 
.A1(n_2034),
.A2(n_1702),
.A3(n_1559),
.B(n_1574),
.Y(n_2199)
);

CKINVDCx20_ASAP7_75t_R g2200 ( 
.A(n_2052),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2037),
.Y(n_2201)
);

OAI322xp33_ASAP7_75t_L g2202 ( 
.A1(n_2034),
.A2(n_589),
.A3(n_581),
.B1(n_590),
.B2(n_591),
.C1(n_583),
.C2(n_557),
.Y(n_2202)
);

OAI32xp33_ASAP7_75t_L g2203 ( 
.A1(n_2074),
.A2(n_15),
.A3(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_2203)
);

AOI21xp33_ASAP7_75t_SL g2204 ( 
.A1(n_2052),
.A2(n_15),
.B(n_16),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2034),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2052),
.B(n_1733),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2034),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2034),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2037),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2074),
.B(n_17),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2034),
.Y(n_2211)
);

NAND2x1p5_ASAP7_75t_L g2212 ( 
.A(n_2047),
.B(n_1540),
.Y(n_2212)
);

A2O1A1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_2074),
.A2(n_590),
.B(n_591),
.C(n_589),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2067),
.B(n_18),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2052),
.B(n_1733),
.Y(n_2215)
);

AOI222xp33_ASAP7_75t_L g2216 ( 
.A1(n_2034),
.A2(n_744),
.B1(n_700),
.B2(n_849),
.C1(n_594),
.C2(n_1700),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2074),
.B(n_18),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2067),
.B(n_19),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_L g2219 ( 
.A1(n_2074),
.A2(n_870),
.B(n_598),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2052),
.B(n_19),
.Y(n_2220)
);

OAI222xp33_ASAP7_75t_L g2221 ( 
.A1(n_2034),
.A2(n_1701),
.B1(n_1700),
.B2(n_1763),
.C1(n_1673),
.C2(n_1689),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2074),
.A2(n_1581),
.B1(n_1573),
.B2(n_1563),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2034),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2034),
.A2(n_879),
.B1(n_884),
.B2(n_870),
.C(n_598),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2052),
.B(n_20),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2105),
.B(n_20),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_2220),
.Y(n_2227)
);

NOR2x1_ASAP7_75t_L g2228 ( 
.A(n_2200),
.B(n_21),
.Y(n_2228)
);

INVx1_ASAP7_75t_SL g2229 ( 
.A(n_2190),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2107),
.B(n_21),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2197),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2146),
.B(n_22),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2214),
.Y(n_2233)
);

NOR2xp67_ASAP7_75t_L g2234 ( 
.A(n_2178),
.B(n_24),
.Y(n_2234)
);

NAND2x1_ASAP7_75t_L g2235 ( 
.A(n_2201),
.B(n_1540),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2188),
.B(n_25),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2218),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2225),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2180),
.B(n_25),
.Y(n_2239)
);

NAND2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2209),
.B(n_1540),
.Y(n_2240)
);

NAND2x1_ASAP7_75t_L g2241 ( 
.A(n_2188),
.B(n_1563),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2135),
.A2(n_1544),
.B1(n_700),
.B2(n_849),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2089),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2183),
.B(n_26),
.Y(n_2244)
);

INVxp67_ASAP7_75t_L g2245 ( 
.A(n_2142),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2096),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2194),
.B(n_2130),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2157),
.Y(n_2248)
);

INVx2_ASAP7_75t_SL g2249 ( 
.A(n_2104),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2191),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2119),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_2196),
.Y(n_2252)
);

AOI21xp33_ASAP7_75t_SL g2253 ( 
.A1(n_2123),
.A2(n_27),
.B(n_30),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2127),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2090),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2204),
.B(n_31),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2118),
.B(n_31),
.Y(n_2257)
);

BUFx2_ASAP7_75t_L g2258 ( 
.A(n_2114),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2176),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_L g2260 ( 
.A(n_2182),
.B(n_32),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2177),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2160),
.B(n_33),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2210),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2120),
.B(n_34),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2139),
.B(n_2132),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2140),
.A2(n_884),
.B(n_879),
.Y(n_2266)
);

NOR2x1_ASAP7_75t_L g2267 ( 
.A(n_2179),
.B(n_35),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_SL g2268 ( 
.A(n_2217),
.B(n_700),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2150),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2126),
.B(n_36),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_2169),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2126),
.B(n_36),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2186),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2189),
.Y(n_2274)
);

INVxp67_ASAP7_75t_L g2275 ( 
.A(n_2145),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2205),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2207),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2208),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2121),
.B(n_37),
.Y(n_2279)
);

NAND2x1_ASAP7_75t_L g2280 ( 
.A(n_2103),
.B(n_1563),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2211),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2109),
.B(n_38),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2097),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_L g2284 ( 
.A(n_2148),
.B(n_38),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2145),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2151),
.B(n_40),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2185),
.B(n_40),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2223),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2143),
.B(n_41),
.Y(n_2289)
);

NOR3xp33_ASAP7_75t_L g2290 ( 
.A(n_2192),
.B(n_955),
.C(n_887),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2163),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2098),
.B(n_41),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2111),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2122),
.B(n_43),
.Y(n_2294)
);

INVxp67_ASAP7_75t_L g2295 ( 
.A(n_2173),
.Y(n_2295)
);

NAND3xp33_ASAP7_75t_L g2296 ( 
.A(n_2110),
.B(n_955),
.C(n_887),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2181),
.B(n_744),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2149),
.A2(n_1544),
.B1(n_744),
.B2(n_849),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2095),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2133),
.B(n_43),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2134),
.B(n_46),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_2116),
.B(n_46),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2206),
.B(n_47),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2095),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2112),
.B(n_47),
.Y(n_2305)
);

AOI22x1_ASAP7_75t_L g2306 ( 
.A1(n_2212),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2088),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_2137),
.B(n_2156),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2136),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2106),
.B(n_50),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2138),
.B(n_51),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2125),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2152),
.B(n_51),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2187),
.B(n_53),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2108),
.B(n_2099),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2213),
.B(n_53),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2172),
.B(n_2159),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2195),
.B(n_54),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2215),
.B(n_54),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2144),
.B(n_55),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_2153),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2128),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2129),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_2102),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2147),
.B(n_57),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2174),
.B(n_57),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2166),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2219),
.B(n_58),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2101),
.B(n_58),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_SL g2330 ( 
.A(n_2115),
.B(n_59),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2164),
.B(n_60),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2203),
.B(n_61),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2087),
.B(n_2117),
.Y(n_2333)
);

INVxp67_ASAP7_75t_L g2334 ( 
.A(n_2167),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2167),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2224),
.B(n_61),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2229),
.B(n_2168),
.Y(n_2337)
);

AOI32xp33_ASAP7_75t_L g2338 ( 
.A1(n_2226),
.A2(n_2198),
.A3(n_2162),
.B1(n_2193),
.B2(n_2184),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2234),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2248),
.B(n_2094),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2234),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2252),
.B(n_2161),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2228),
.B(n_2091),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2335),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2253),
.B(n_2249),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2306),
.Y(n_2346)
);

INVx1_ASAP7_75t_SL g2347 ( 
.A(n_2321),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2253),
.B(n_2158),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2269),
.B(n_2155),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2257),
.B(n_2230),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2289),
.B(n_2113),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2307),
.B(n_2154),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2258),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2285),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2267),
.Y(n_2355)
);

NAND2xp33_ASAP7_75t_L g2356 ( 
.A(n_2247),
.B(n_2170),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2239),
.B(n_2131),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2331),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2244),
.B(n_2092),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2305),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2275),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2302),
.Y(n_2362)
);

NAND3xp33_ASAP7_75t_L g2363 ( 
.A(n_2290),
.B(n_2216),
.C(n_2171),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2232),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_R g2365 ( 
.A(n_2250),
.B(n_2202),
.Y(n_2365)
);

NAND2x1_ASAP7_75t_L g2366 ( 
.A(n_2231),
.B(n_2222),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2236),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2233),
.B(n_2100),
.Y(n_2368)
);

AOI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2332),
.A2(n_2141),
.B1(n_2165),
.B2(n_2175),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2303),
.B(n_2199),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2237),
.B(n_2124),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2309),
.B(n_2093),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2256),
.Y(n_2373)
);

NAND2x1p5_ASAP7_75t_L g2374 ( 
.A(n_2283),
.B(n_1643),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2243),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2284),
.B(n_62),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2241),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2294),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2279),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2286),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2245),
.B(n_62),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2319),
.B(n_2221),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2265),
.B(n_663),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2262),
.Y(n_2384)
);

AND2x4_ASAP7_75t_SL g2385 ( 
.A(n_2270),
.B(n_1573),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2291),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2251),
.B(n_63),
.Y(n_2387)
);

INVxp67_ASAP7_75t_L g2388 ( 
.A(n_2268),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2260),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2272),
.B(n_63),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2292),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2271),
.B(n_64),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2327),
.B(n_64),
.Y(n_2393)
);

NAND2xp33_ASAP7_75t_L g2394 ( 
.A(n_2324),
.B(n_1544),
.Y(n_2394)
);

INVxp33_ASAP7_75t_L g2395 ( 
.A(n_2301),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2255),
.B(n_65),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2254),
.Y(n_2397)
);

NAND4xp25_ASAP7_75t_L g2398 ( 
.A(n_2238),
.B(n_70),
.C(n_66),
.D(n_67),
.Y(n_2398)
);

INVx1_ASAP7_75t_SL g2399 ( 
.A(n_2330),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2227),
.B(n_67),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2235),
.Y(n_2401)
);

INVxp67_ASAP7_75t_L g2402 ( 
.A(n_2268),
.Y(n_2402)
);

NAND2x1_ASAP7_75t_SL g2403 ( 
.A(n_2259),
.B(n_2261),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2273),
.B(n_73),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2325),
.Y(n_2405)
);

OAI21xp33_ASAP7_75t_L g2406 ( 
.A1(n_2308),
.A2(n_1581),
.B(n_1573),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2333),
.B(n_663),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2263),
.B(n_73),
.Y(n_2408)
);

INVx1_ASAP7_75t_SL g2409 ( 
.A(n_2282),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2274),
.B(n_75),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2276),
.B(n_76),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2314),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2334),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2318),
.A2(n_1544),
.B1(n_663),
.B2(n_1567),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2328),
.B(n_76),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_2264),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2277),
.B(n_79),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2315),
.Y(n_2418)
);

OAI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2280),
.A2(n_546),
.B1(n_604),
.B2(n_548),
.C(n_532),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2311),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2300),
.Y(n_2421)
);

HB1xp67_ASAP7_75t_L g2422 ( 
.A(n_2278),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2313),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2310),
.B(n_2312),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2326),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2287),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2322),
.B(n_79),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2323),
.B(n_80),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_SL g2429 ( 
.A(n_2297),
.B(n_616),
.C(n_605),
.Y(n_2429)
);

INVxp33_ASAP7_75t_L g2430 ( 
.A(n_2317),
.Y(n_2430)
);

INVxp67_ASAP7_75t_SL g2431 ( 
.A(n_2266),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2320),
.B(n_81),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2281),
.B(n_663),
.Y(n_2433)
);

CKINVDCx14_ASAP7_75t_R g2434 ( 
.A(n_2293),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2296),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2288),
.B(n_81),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2299),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2296),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2336),
.B(n_82),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2295),
.A2(n_1717),
.B1(n_1567),
.B2(n_1689),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2316),
.Y(n_2441)
);

NAND3xp33_ASAP7_75t_L g2442 ( 
.A(n_2246),
.B(n_691),
.C(n_536),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2329),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_2240),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2304),
.B(n_83),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_2242),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2298),
.B(n_663),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2228),
.B(n_84),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2253),
.B(n_85),
.Y(n_2449)
);

OAI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2275),
.A2(n_624),
.B1(n_636),
.B2(n_630),
.C(n_618),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2228),
.B(n_85),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2253),
.B(n_87),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2306),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2306),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2234),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2229),
.B(n_87),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2228),
.B(n_90),
.Y(n_2457)
);

OR2x2_ASAP7_75t_L g2458 ( 
.A(n_2229),
.B(n_91),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2229),
.B(n_91),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2226),
.A2(n_1664),
.B(n_92),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2234),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2234),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2234),
.Y(n_2463)
);

INVx5_ASAP7_75t_L g2464 ( 
.A(n_2269),
.Y(n_2464)
);

INVx3_ASAP7_75t_L g2465 ( 
.A(n_2226),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2228),
.B(n_93),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2253),
.B(n_94),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2234),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2234),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2234),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2347),
.B(n_95),
.Y(n_2471)
);

NOR2x1p5_ASAP7_75t_L g2472 ( 
.A(n_2346),
.B(n_95),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2353),
.B(n_96),
.Y(n_2473)
);

NOR3xp33_ASAP7_75t_L g2474 ( 
.A(n_2429),
.B(n_639),
.C(n_638),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2390),
.B(n_96),
.Y(n_2475)
);

AOI222xp33_ASAP7_75t_L g2476 ( 
.A1(n_2361),
.A2(n_2344),
.B1(n_2354),
.B2(n_2413),
.C1(n_2389),
.C2(n_2341),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_SL g2477 ( 
.A(n_2386),
.B(n_97),
.C(n_99),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2350),
.Y(n_2478)
);

NOR2xp67_ASAP7_75t_L g2479 ( 
.A(n_2464),
.B(n_97),
.Y(n_2479)
);

NAND3xp33_ASAP7_75t_L g2480 ( 
.A(n_2464),
.B(n_691),
.C(n_536),
.Y(n_2480)
);

AOI221xp5_ASAP7_75t_SL g2481 ( 
.A1(n_2434),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.C(n_102),
.Y(n_2481)
);

NAND3xp33_ASAP7_75t_L g2482 ( 
.A(n_2464),
.B(n_691),
.C(n_536),
.Y(n_2482)
);

NOR4xp25_ASAP7_75t_L g2483 ( 
.A(n_2355),
.B(n_103),
.C(n_101),
.D(n_102),
.Y(n_2483)
);

XNOR2xp5_ASAP7_75t_L g2484 ( 
.A(n_2430),
.B(n_103),
.Y(n_2484)
);

AOI222xp33_ASAP7_75t_L g2485 ( 
.A1(n_2339),
.A2(n_848),
.B1(n_691),
.B2(n_871),
.C1(n_741),
.C2(n_536),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2456),
.B(n_104),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2459),
.Y(n_2487)
);

NAND4xp25_ASAP7_75t_L g2488 ( 
.A(n_2337),
.B(n_106),
.C(n_104),
.D(n_105),
.Y(n_2488)
);

OAI31xp33_ASAP7_75t_L g2489 ( 
.A1(n_2465),
.A2(n_109),
.A3(n_106),
.B(n_108),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2449),
.B(n_108),
.Y(n_2490)
);

NOR3xp33_ASAP7_75t_L g2491 ( 
.A(n_2465),
.B(n_652),
.C(n_642),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2452),
.B(n_109),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2467),
.B(n_110),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_SL g2494 ( 
.A(n_2398),
.B(n_1544),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2445),
.B(n_111),
.Y(n_2495)
);

AOI211xp5_ASAP7_75t_L g2496 ( 
.A1(n_2422),
.A2(n_114),
.B(n_111),
.C(n_113),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2358),
.B(n_2399),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2345),
.B(n_113),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2448),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2352),
.B(n_114),
.Y(n_2500)
);

OAI211xp5_ASAP7_75t_L g2501 ( 
.A1(n_2403),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2396),
.B(n_115),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2451),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2404),
.B(n_116),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2342),
.B(n_117),
.Y(n_2505)
);

NAND3xp33_ASAP7_75t_SL g2506 ( 
.A(n_2365),
.B(n_669),
.C(n_668),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2457),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2410),
.B(n_118),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2466),
.Y(n_2509)
);

O2A1O1Ixp33_ASAP7_75t_L g2510 ( 
.A1(n_2376),
.A2(n_124),
.B(n_119),
.C(n_120),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2349),
.B(n_120),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_L g2512 ( 
.A(n_2338),
.B(n_741),
.C(n_691),
.Y(n_2512)
);

XNOR2x1_ASAP7_75t_L g2513 ( 
.A(n_2409),
.B(n_124),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2397),
.B(n_125),
.Y(n_2514)
);

AOI21xp33_ASAP7_75t_L g2515 ( 
.A1(n_2395),
.A2(n_695),
.B(n_683),
.Y(n_2515)
);

NOR3xp33_ASAP7_75t_L g2516 ( 
.A(n_2388),
.B(n_716),
.C(n_709),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2458),
.B(n_125),
.Y(n_2517)
);

OR2x2_ASAP7_75t_L g2518 ( 
.A(n_2427),
.B(n_126),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2411),
.B(n_126),
.Y(n_2519)
);

NAND2x1_ASAP7_75t_L g2520 ( 
.A(n_2453),
.B(n_127),
.Y(n_2520)
);

NAND3xp33_ASAP7_75t_L g2521 ( 
.A(n_2338),
.B(n_848),
.C(n_741),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2417),
.Y(n_2522)
);

NAND4xp75_ASAP7_75t_L g2523 ( 
.A(n_2424),
.B(n_130),
.C(n_127),
.D(n_128),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2454),
.B(n_132),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_SL g2525 ( 
.A1(n_2375),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2525)
);

NOR4xp25_ASAP7_75t_SL g2526 ( 
.A(n_2360),
.B(n_136),
.C(n_133),
.D(n_135),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2436),
.B(n_135),
.Y(n_2527)
);

NAND3xp33_ASAP7_75t_L g2528 ( 
.A(n_2356),
.B(n_848),
.C(n_741),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_2402),
.B(n_731),
.C(n_726),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2405),
.B(n_137),
.Y(n_2530)
);

NOR2xp67_ASAP7_75t_L g2531 ( 
.A(n_2377),
.B(n_138),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2366),
.A2(n_737),
.B1(n_745),
.B2(n_735),
.Y(n_2532)
);

NOR3xp33_ASAP7_75t_L g2533 ( 
.A(n_2416),
.B(n_751),
.C(n_747),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2364),
.A2(n_1557),
.B1(n_663),
.B2(n_848),
.Y(n_2534)
);

NOR2xp67_ASAP7_75t_L g2535 ( 
.A(n_2428),
.B(n_138),
.Y(n_2535)
);

INVxp67_ASAP7_75t_SL g2536 ( 
.A(n_2348),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_2437),
.B(n_139),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2444),
.B(n_140),
.Y(n_2538)
);

AOI221xp5_ASAP7_75t_L g2539 ( 
.A1(n_2425),
.A2(n_871),
.B1(n_741),
.B2(n_760),
.C(n_761),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2455),
.Y(n_2540)
);

AOI21xp33_ASAP7_75t_L g2541 ( 
.A1(n_2461),
.A2(n_2463),
.B(n_2462),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_2387),
.A2(n_2381),
.B(n_2450),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2373),
.A2(n_871),
.B1(n_783),
.B2(n_785),
.C(n_762),
.Y(n_2543)
);

NAND4xp25_ASAP7_75t_L g2544 ( 
.A(n_2371),
.B(n_143),
.C(n_141),
.D(n_142),
.Y(n_2544)
);

NOR4xp25_ASAP7_75t_L g2545 ( 
.A(n_2418),
.B(n_149),
.C(n_147),
.D(n_148),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2468),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2401),
.B(n_871),
.Y(n_2547)
);

OAI211xp5_ASAP7_75t_SL g2548 ( 
.A1(n_2476),
.A2(n_2379),
.B(n_2438),
.C(n_2435),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2479),
.Y(n_2549)
);

AOI322xp5_ASAP7_75t_L g2550 ( 
.A1(n_2536),
.A2(n_2391),
.A3(n_2441),
.B1(n_2470),
.B2(n_2469),
.C1(n_2423),
.C2(n_2421),
.Y(n_2550)
);

OAI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2501),
.A2(n_2363),
.B(n_2460),
.Y(n_2551)
);

AOI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2532),
.A2(n_2392),
.B(n_2400),
.Y(n_2552)
);

OAI21x1_ASAP7_75t_L g2553 ( 
.A1(n_2520),
.A2(n_2359),
.B(n_2343),
.Y(n_2553)
);

OAI321xp33_ASAP7_75t_L g2554 ( 
.A1(n_2497),
.A2(n_2369),
.A3(n_2368),
.B1(n_2426),
.B2(n_2372),
.C(n_2362),
.Y(n_2554)
);

AOI221xp5_ASAP7_75t_L g2555 ( 
.A1(n_2541),
.A2(n_2420),
.B1(n_2431),
.B2(n_2367),
.C(n_2378),
.Y(n_2555)
);

AOI211x1_ASAP7_75t_L g2556 ( 
.A1(n_2542),
.A2(n_2382),
.B(n_2406),
.C(n_2384),
.Y(n_2556)
);

AOI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2499),
.A2(n_2380),
.B1(n_2414),
.B2(n_2412),
.Y(n_2557)
);

OAI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2540),
.A2(n_2393),
.B1(n_2369),
.B2(n_2419),
.C(n_2340),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2506),
.B(n_2407),
.C(n_2408),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_SL g2560 ( 
.A1(n_2478),
.A2(n_2370),
.B1(n_2443),
.B2(n_2385),
.Y(n_2560)
);

OAI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2538),
.A2(n_2357),
.B(n_2351),
.Y(n_2561)
);

AOI221x1_ASAP7_75t_L g2562 ( 
.A1(n_2491),
.A2(n_2439),
.B1(n_2415),
.B2(n_2442),
.C(n_2432),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2472),
.Y(n_2563)
);

AOI221xp5_ASAP7_75t_L g2564 ( 
.A1(n_2546),
.A2(n_2383),
.B1(n_2433),
.B2(n_2446),
.C(n_2447),
.Y(n_2564)
);

OAI32xp33_ASAP7_75t_L g2565 ( 
.A1(n_2498),
.A2(n_2374),
.A3(n_2440),
.B1(n_2394),
.B2(n_2414),
.Y(n_2565)
);

AOI211xp5_ASAP7_75t_SL g2566 ( 
.A1(n_2471),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_2566)
);

NAND3xp33_ASAP7_75t_L g2567 ( 
.A(n_2481),
.B(n_2477),
.C(n_2496),
.Y(n_2567)
);

INVx1_ASAP7_75t_SL g2568 ( 
.A(n_2500),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_R g2569 ( 
.A(n_2473),
.B(n_2484),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2483),
.B(n_2545),
.Y(n_2570)
);

NAND4xp25_ASAP7_75t_L g2571 ( 
.A(n_2524),
.B(n_152),
.C(n_150),
.D(n_151),
.Y(n_2571)
);

NOR2x1_ASAP7_75t_L g2572 ( 
.A(n_2488),
.B(n_154),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2537),
.B(n_154),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2537),
.B(n_2511),
.Y(n_2574)
);

AOI211xp5_ASAP7_75t_SL g2575 ( 
.A1(n_2487),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2575)
);

XNOR2xp5_ASAP7_75t_L g2576 ( 
.A(n_2513),
.B(n_155),
.Y(n_2576)
);

AOI221xp5_ASAP7_75t_L g2577 ( 
.A1(n_2503),
.A2(n_2509),
.B1(n_2507),
.B2(n_2522),
.C(n_2517),
.Y(n_2577)
);

O2A1O1Ixp33_ASAP7_75t_L g2578 ( 
.A1(n_2525),
.A2(n_162),
.B(n_158),
.C(n_159),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2514),
.B(n_162),
.Y(n_2579)
);

INVxp33_ASAP7_75t_SL g2580 ( 
.A(n_2505),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2527),
.B(n_164),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2496),
.B(n_871),
.C(n_790),
.Y(n_2582)
);

NOR3xp33_ASAP7_75t_L g2583 ( 
.A(n_2544),
.B(n_793),
.C(n_753),
.Y(n_2583)
);

AOI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2533),
.A2(n_805),
.B1(n_814),
.B2(n_800),
.C(n_794),
.Y(n_2584)
);

OAI221xp5_ASAP7_75t_L g2585 ( 
.A1(n_2530),
.A2(n_860),
.B1(n_864),
.B2(n_859),
.C(n_845),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2535),
.A2(n_914),
.B1(n_919),
.B2(n_868),
.Y(n_2586)
);

INVx3_ASAP7_75t_L g2587 ( 
.A(n_2518),
.Y(n_2587)
);

INVx1_ASAP7_75t_SL g2588 ( 
.A(n_2486),
.Y(n_2588)
);

A2O1A1Ixp33_ASAP7_75t_SL g2589 ( 
.A1(n_2516),
.A2(n_2529),
.B(n_2474),
.C(n_2489),
.Y(n_2589)
);

OAI221xp5_ASAP7_75t_L g2590 ( 
.A1(n_2490),
.A2(n_940),
.B1(n_930),
.B2(n_170),
.C(n_168),
.Y(n_2590)
);

NAND4xp25_ASAP7_75t_L g2591 ( 
.A(n_2510),
.B(n_172),
.C(n_169),
.D(n_171),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2502),
.A2(n_171),
.B(n_172),
.Y(n_2592)
);

AOI221xp5_ASAP7_75t_L g2593 ( 
.A1(n_2539),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.C(n_176),
.Y(n_2593)
);

NOR2x1p5_ASAP7_75t_L g2594 ( 
.A(n_2523),
.B(n_173),
.Y(n_2594)
);

OAI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2492),
.A2(n_1051),
.B1(n_1041),
.B2(n_181),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2526),
.B(n_180),
.Y(n_2596)
);

OAI211xp5_ASAP7_75t_L g2597 ( 
.A1(n_2543),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2597)
);

AOI222xp33_ASAP7_75t_L g2598 ( 
.A1(n_2531),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.C1(n_186),
.C2(n_188),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2475),
.B(n_188),
.Y(n_2599)
);

OAI221xp5_ASAP7_75t_SL g2600 ( 
.A1(n_2550),
.A2(n_2534),
.B1(n_2493),
.B2(n_2482),
.C(n_2480),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2576),
.Y(n_2601)
);

OAI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2548),
.A2(n_2494),
.B1(n_2508),
.B2(n_2519),
.C(n_2504),
.Y(n_2602)
);

AOI221x1_ASAP7_75t_SL g2603 ( 
.A1(n_2567),
.A2(n_2512),
.B1(n_2521),
.B2(n_2495),
.C(n_2528),
.Y(n_2603)
);

OAI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2555),
.A2(n_2515),
.B1(n_2547),
.B2(n_2485),
.C(n_192),
.Y(n_2604)
);

BUFx2_ASAP7_75t_L g2605 ( 
.A(n_2569),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2549),
.A2(n_2580),
.B1(n_2563),
.B2(n_2587),
.Y(n_2606)
);

OAI221xp5_ASAP7_75t_SL g2607 ( 
.A1(n_2558),
.A2(n_194),
.B1(n_189),
.B2(n_190),
.C(n_196),
.Y(n_2607)
);

AOI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2587),
.A2(n_1051),
.B1(n_1041),
.B2(n_1662),
.Y(n_2608)
);

BUFx12f_ASAP7_75t_L g2609 ( 
.A(n_2594),
.Y(n_2609)
);

AOI222xp33_ASAP7_75t_L g2610 ( 
.A1(n_2570),
.A2(n_189),
.B1(n_190),
.B2(n_194),
.C1(n_196),
.C2(n_197),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2554),
.B(n_197),
.Y(n_2611)
);

AOI221xp5_ASAP7_75t_L g2612 ( 
.A1(n_2565),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_201),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2588),
.A2(n_1037),
.B1(n_1650),
.B2(n_203),
.Y(n_2613)
);

AOI221x1_ASAP7_75t_SL g2614 ( 
.A1(n_2574),
.A2(n_203),
.B1(n_200),
.B2(n_202),
.C(n_205),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2566),
.B(n_202),
.Y(n_2615)
);

NAND3xp33_ASAP7_75t_SL g2616 ( 
.A(n_2568),
.B(n_206),
.C(n_207),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2596),
.Y(n_2617)
);

AOI211xp5_ASAP7_75t_L g2618 ( 
.A1(n_2578),
.A2(n_213),
.B(n_210),
.C(n_212),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2579),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2589),
.A2(n_212),
.B(n_213),
.Y(n_2620)
);

AOI222xp33_ASAP7_75t_L g2621 ( 
.A1(n_2551),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.C1(n_220),
.C2(n_221),
.Y(n_2621)
);

AOI211xp5_ASAP7_75t_L g2622 ( 
.A1(n_2595),
.A2(n_223),
.B(n_217),
.C(n_219),
.Y(n_2622)
);

NAND4xp25_ASAP7_75t_L g2623 ( 
.A(n_2556),
.B(n_227),
.C(n_225),
.D(n_226),
.Y(n_2623)
);

OAI211xp5_ASAP7_75t_L g2624 ( 
.A1(n_2560),
.A2(n_228),
.B(n_225),
.C(n_226),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2577),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_2625)
);

AOI211xp5_ASAP7_75t_L g2626 ( 
.A1(n_2590),
.A2(n_236),
.B(n_232),
.C(n_234),
.Y(n_2626)
);

INVx1_ASAP7_75t_SL g2627 ( 
.A(n_2573),
.Y(n_2627)
);

NAND4xp25_ASAP7_75t_SL g2628 ( 
.A(n_2572),
.B(n_239),
.C(n_237),
.D(n_238),
.Y(n_2628)
);

NOR2x1_ASAP7_75t_L g2629 ( 
.A(n_2571),
.B(n_240),
.Y(n_2629)
);

XNOR2x1_ASAP7_75t_L g2630 ( 
.A(n_2553),
.B(n_241),
.Y(n_2630)
);

AOI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2585),
.A2(n_241),
.B(n_242),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2559),
.A2(n_248),
.B1(n_244),
.B2(n_245),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2599),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2605),
.B(n_2561),
.Y(n_2634)
);

AOI222xp33_ASAP7_75t_L g2635 ( 
.A1(n_2617),
.A2(n_2564),
.B1(n_2582),
.B2(n_2586),
.C1(n_2581),
.C2(n_2593),
.Y(n_2635)
);

NOR3xp33_ASAP7_75t_SL g2636 ( 
.A(n_2623),
.B(n_2552),
.C(n_2597),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2630),
.Y(n_2637)
);

O2A1O1Ixp33_ASAP7_75t_L g2638 ( 
.A1(n_2611),
.A2(n_2620),
.B(n_2601),
.C(n_2624),
.Y(n_2638)
);

NAND3xp33_ASAP7_75t_L g2639 ( 
.A(n_2606),
.B(n_2557),
.C(n_2575),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_L g2640 ( 
.A1(n_2627),
.A2(n_2591),
.B1(n_2583),
.B2(n_2592),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2614),
.B(n_2598),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2619),
.Y(n_2642)
);

NAND3xp33_ASAP7_75t_L g2643 ( 
.A(n_2612),
.B(n_2562),
.C(n_2584),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2629),
.Y(n_2644)
);

XNOR2xp5_ASAP7_75t_L g2645 ( 
.A(n_2618),
.B(n_251),
.Y(n_2645)
);

OAI21xp33_ASAP7_75t_SL g2646 ( 
.A1(n_2628),
.A2(n_251),
.B(n_252),
.Y(n_2646)
);

AOI221xp5_ASAP7_75t_L g2647 ( 
.A1(n_2602),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.C(n_255),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2625),
.A2(n_253),
.B(n_254),
.Y(n_2648)
);

OAI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2616),
.A2(n_256),
.B(n_259),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2615),
.Y(n_2650)
);

O2A1O1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2607),
.A2(n_260),
.B(n_256),
.C(n_259),
.Y(n_2651)
);

INVx1_ASAP7_75t_SL g2652 ( 
.A(n_2634),
.Y(n_2652)
);

OR4x2_ASAP7_75t_L g2653 ( 
.A(n_2634),
.B(n_2609),
.C(n_2626),
.D(n_2610),
.Y(n_2653)
);

AND3x2_ASAP7_75t_L g2654 ( 
.A(n_2644),
.B(n_2622),
.C(n_2621),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2641),
.B(n_2627),
.Y(n_2655)
);

CKINVDCx16_ASAP7_75t_R g2656 ( 
.A(n_2637),
.Y(n_2656)
);

NAND5xp2_ASAP7_75t_L g2657 ( 
.A(n_2638),
.B(n_2600),
.C(n_2604),
.D(n_2631),
.E(n_2632),
.Y(n_2657)
);

OAI221xp5_ASAP7_75t_L g2658 ( 
.A1(n_2639),
.A2(n_2603),
.B1(n_2633),
.B2(n_2608),
.C(n_2613),
.Y(n_2658)
);

AOI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2650),
.A2(n_264),
.B1(n_260),
.B2(n_261),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2642),
.B(n_261),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2646),
.B(n_265),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2645),
.Y(n_2662)
);

NOR2x1_ASAP7_75t_L g2663 ( 
.A(n_2643),
.B(n_266),
.Y(n_2663)
);

NOR3xp33_ASAP7_75t_L g2664 ( 
.A(n_2647),
.B(n_267),
.C(n_268),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2636),
.Y(n_2665)
);

AND2x2_ASAP7_75t_SL g2666 ( 
.A(n_2640),
.B(n_269),
.Y(n_2666)
);

OAI221xp5_ASAP7_75t_L g2667 ( 
.A1(n_2652),
.A2(n_2649),
.B1(n_2651),
.B2(n_2648),
.C(n_2635),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_2656),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2660),
.Y(n_2669)
);

CKINVDCx20_ASAP7_75t_R g2670 ( 
.A(n_2655),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2661),
.Y(n_2671)
);

AO221x1_ASAP7_75t_L g2672 ( 
.A1(n_2665),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.C(n_274),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2662),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_L g2674 ( 
.A(n_2666),
.Y(n_2674)
);

CKINVDCx20_ASAP7_75t_R g2675 ( 
.A(n_2659),
.Y(n_2675)
);

OAI22xp33_ASAP7_75t_SL g2676 ( 
.A1(n_2663),
.A2(n_275),
.B1(n_272),
.B2(n_274),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2653),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2654),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2658),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2657),
.Y(n_2680)
);

INVx6_ASAP7_75t_L g2681 ( 
.A(n_2664),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2652),
.B(n_275),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2652),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2668),
.B(n_277),
.Y(n_2684)
);

OAI22xp5_ASAP7_75t_L g2685 ( 
.A1(n_2670),
.A2(n_281),
.B1(n_278),
.B2(n_280),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2682),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_SL g2687 ( 
.A(n_2677),
.B(n_283),
.Y(n_2687)
);

AO21x2_ASAP7_75t_L g2688 ( 
.A1(n_2683),
.A2(n_284),
.B(n_285),
.Y(n_2688)
);

XOR2xp5_ASAP7_75t_L g2689 ( 
.A(n_2680),
.B(n_286),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2672),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2678),
.A2(n_2673),
.B1(n_2667),
.B2(n_2679),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2674),
.Y(n_2692)
);

OAI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2675),
.A2(n_2681),
.B1(n_2671),
.B2(n_2669),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2674),
.Y(n_2694)
);

XNOR2xp5_ASAP7_75t_L g2695 ( 
.A(n_2676),
.B(n_286),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2674),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2681),
.A2(n_1037),
.B1(n_289),
.B2(n_287),
.Y(n_2697)
);

XOR2xp5_ASAP7_75t_L g2698 ( 
.A(n_2668),
.B(n_287),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2668),
.A2(n_1037),
.B1(n_291),
.B2(n_288),
.Y(n_2699)
);

OAI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2668),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_2700)
);

NAND3xp33_ASAP7_75t_L g2701 ( 
.A(n_2691),
.B(n_1037),
.C(n_294),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2690),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2688),
.Y(n_2703)
);

OAI22xp5_ASAP7_75t_SL g2704 ( 
.A1(n_2689),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2686),
.Y(n_2705)
);

CKINVDCx20_ASAP7_75t_R g2706 ( 
.A(n_2693),
.Y(n_2706)
);

OAI22x1_ASAP7_75t_L g2707 ( 
.A1(n_2695),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_2707)
);

HB1xp67_ASAP7_75t_L g2708 ( 
.A(n_2698),
.Y(n_2708)
);

OR3x2_ASAP7_75t_L g2709 ( 
.A(n_2692),
.B(n_302),
.C(n_303),
.Y(n_2709)
);

OAI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2694),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_2710)
);

NOR3xp33_ASAP7_75t_L g2711 ( 
.A(n_2696),
.B(n_304),
.C(n_305),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2684),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2687),
.B(n_2697),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2705),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_2703),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2709),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2706),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2707),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2704),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2708),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2712),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2713),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2702),
.Y(n_2723)
);

INVxp67_ASAP7_75t_SL g2724 ( 
.A(n_2711),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2710),
.B(n_2700),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2714),
.A2(n_2720),
.B1(n_2717),
.B2(n_2722),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2715),
.A2(n_2701),
.B1(n_2699),
.B2(n_2685),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2721),
.A2(n_306),
.B(n_310),
.Y(n_2728)
);

HB1xp67_ASAP7_75t_L g2729 ( 
.A(n_2716),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2718),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2719),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2724),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2723),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_2733)
);

AO22x1_ASAP7_75t_L g2734 ( 
.A1(n_2725),
.A2(n_316),
.B1(n_320),
.B2(n_321),
.Y(n_2734)
);

INVx4_ASAP7_75t_L g2735 ( 
.A(n_2714),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2714),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_SL g2737 ( 
.A1(n_2714),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2735),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_2738)
);

AOI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2732),
.A2(n_327),
.B1(n_328),
.B2(n_330),
.C(n_331),
.Y(n_2739)
);

OR2x2_ASAP7_75t_L g2740 ( 
.A(n_2729),
.B(n_331),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2726),
.Y(n_2741)
);

OAI21x1_ASAP7_75t_L g2742 ( 
.A1(n_2736),
.A2(n_334),
.B(n_335),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2731),
.A2(n_334),
.B1(n_337),
.B2(n_339),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2730),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2727),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_2745)
);

OAI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2728),
.A2(n_343),
.B(n_344),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2734),
.A2(n_345),
.B(n_346),
.Y(n_2747)
);

OAI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2733),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2740),
.Y(n_2749)
);

INVxp67_ASAP7_75t_SL g2750 ( 
.A(n_2742),
.Y(n_2750)
);

HB1xp67_ASAP7_75t_L g2751 ( 
.A(n_2746),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2745),
.A2(n_2738),
.B1(n_2748),
.B2(n_2743),
.Y(n_2752)
);

O2A1O1Ixp33_ASAP7_75t_L g2753 ( 
.A1(n_2747),
.A2(n_2737),
.B(n_351),
.C(n_352),
.Y(n_2753)
);

OAI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_2744),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_2754)
);

NAND5xp2_ASAP7_75t_L g2755 ( 
.A(n_2739),
.B(n_354),
.C(n_355),
.D(n_356),
.E(n_357),
.Y(n_2755)
);

OAI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2741),
.A2(n_354),
.B1(n_355),
.B2(n_357),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2741),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2749),
.Y(n_2758)
);

OA22x2_ASAP7_75t_L g2759 ( 
.A1(n_2750),
.A2(n_359),
.B1(n_361),
.B2(n_362),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2751),
.Y(n_2760)
);

AOI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_2755),
.A2(n_367),
.B1(n_368),
.B2(n_370),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2754),
.A2(n_2752),
.B1(n_2756),
.B2(n_2753),
.Y(n_2762)
);

OAI222xp33_ASAP7_75t_L g2763 ( 
.A1(n_2757),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.C1(n_373),
.C2(n_374),
.Y(n_2763)
);

OAI21xp5_ASAP7_75t_SL g2764 ( 
.A1(n_2757),
.A2(n_371),
.B(n_373),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2760),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_2765)
);

OAI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2758),
.A2(n_375),
.B1(n_376),
.B2(n_378),
.Y(n_2766)
);

NAND3xp33_ASAP7_75t_L g2767 ( 
.A(n_2762),
.B(n_379),
.C(n_380),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2767),
.B(n_2761),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2768),
.A2(n_2764),
.B(n_2759),
.Y(n_2769)
);

AOI211xp5_ASAP7_75t_L g2770 ( 
.A1(n_2769),
.A2(n_2766),
.B(n_2763),
.C(n_2765),
.Y(n_2770)
);


endmodule