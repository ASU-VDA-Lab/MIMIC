module fake_jpeg_31583_n_493 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_493);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_493;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_16),
.B(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_4),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_85),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_76),
.Y(n_140)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_82),
.Y(n_133)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_7),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_37),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_7),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_93),
.Y(n_113)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

BUFx6f_ASAP7_75t_SL g92 ( 
.A(n_44),
.Y(n_92)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_3),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_29),
.CON(n_105),
.SN(n_105)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_95),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_128),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_112),
.B(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_36),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_34),
.B(n_40),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_125),
.A2(n_40),
.B(n_38),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_41),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_52),
.B(n_36),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_76),
.B(n_41),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_46),
.Y(n_192)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_46),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_44),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_163),
.Y(n_210)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_154),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_15),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_160),
.Y(n_201)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_110),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_47),
.B(n_39),
.Y(n_162)
);

NOR2x1_ASAP7_75t_R g219 ( 
.A(n_162),
.B(n_184),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_32),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_168),
.A2(n_177),
.B1(n_190),
.B2(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_15),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_46),
.Y(n_209)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_176),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_191),
.Y(n_220)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_175),
.Y(n_218)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_121),
.A2(n_82),
.B1(n_86),
.B2(n_40),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_181),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_140),
.B(n_148),
.Y(n_225)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_94),
.C(n_69),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_103),
.C(n_135),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_111),
.B(n_42),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_188),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_113),
.A2(n_47),
.B(n_42),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_132),
.A2(n_73),
.B1(n_77),
.B2(n_75),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_189),
.B1(n_195),
.B2(n_119),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_63),
.B1(n_56),
.B2(n_54),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_101),
.A2(n_51),
.B1(n_79),
.B2(n_38),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_196),
.B1(n_147),
.B2(n_118),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_101),
.A2(n_38),
.B1(n_37),
.B2(n_32),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_26),
.B1(n_37),
.B2(n_32),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_98),
.B1(n_147),
.B2(n_148),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_152),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_204),
.A2(n_165),
.B1(n_173),
.B2(n_178),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_156),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_97),
.B1(n_152),
.B2(n_140),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_142),
.B1(n_97),
.B2(n_151),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_216),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_151),
.B1(n_119),
.B2(n_150),
.Y(n_216)
);

AND2x4_ASAP7_75t_SL g224 ( 
.A(n_153),
.B(n_120),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_225),
.A2(n_170),
.B(n_133),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_231),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_150),
.B1(n_141),
.B2(n_135),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_237),
.B1(n_161),
.B2(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_153),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_153),
.A2(n_141),
.B1(n_102),
.B2(n_109),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_235),
.B1(n_195),
.B2(n_187),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_158),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_133),
.B1(n_118),
.B2(n_45),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_239),
.B(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_248),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_255),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_242),
.A2(n_232),
.B1(n_221),
.B2(n_222),
.Y(n_300)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_160),
.C(n_182),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_262),
.C(n_247),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_210),
.C(n_224),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_186),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_198),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_166),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_185),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_167),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_205),
.B(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_201),
.B(n_163),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_257),
.B(n_273),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_207),
.B1(n_228),
.B2(n_193),
.Y(n_304)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_212),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_263),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_191),
.C(n_174),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_230),
.Y(n_263)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_267),
.Y(n_297)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_217),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_219),
.B(n_238),
.Y(n_266)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_225),
.B(n_210),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_212),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_272),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_214),
.B1(n_207),
.B2(n_226),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_179),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_268),
.B(n_244),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_285),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_204),
.B1(n_234),
.B2(n_216),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_291),
.B1(n_296),
.B2(n_303),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_210),
.B(n_215),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_283),
.A2(n_286),
.B(n_306),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_245),
.A2(n_211),
.B(n_224),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_236),
.B1(n_223),
.B2(n_224),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_219),
.C(n_227),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_305),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_256),
.B1(n_270),
.B2(n_261),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_221),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_304),
.B1(n_253),
.B2(n_263),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_239),
.B(n_226),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_301),
.Y(n_336)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_256),
.A2(n_176),
.B1(n_181),
.B2(n_159),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_250),
.B(n_228),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_155),
.B(n_157),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_314),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_249),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_311),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_312),
.A2(n_274),
.B(n_284),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_241),
.B1(n_244),
.B2(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_322),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_292),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_326),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_258),
.B1(n_242),
.B2(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_318),
.A2(n_320),
.B1(n_321),
.B2(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_271),
.B1(n_251),
.B2(n_254),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_271),
.B1(n_266),
.B2(n_240),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_248),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_283),
.A2(n_271),
.B1(n_255),
.B2(n_272),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_263),
.B1(n_273),
.B2(n_269),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_324),
.A2(n_318),
.B1(n_323),
.B2(n_313),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_306),
.A2(n_265),
.B(n_269),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_332),
.B(n_294),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_287),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_328),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_299),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_330),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_267),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_335),
.Y(n_369)
);

A2O1A1O1Ixp25_ASAP7_75t_L g332 ( 
.A1(n_290),
.A2(n_267),
.B(n_264),
.C(n_260),
.D(n_243),
.Y(n_332)
);

INVx11_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_337),
.Y(n_354)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_339),
.B(n_295),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_275),
.C(n_298),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_349),
.C(n_364),
.Y(n_375)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_343),
.A2(n_348),
.B(n_351),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_345),
.A2(n_307),
.B1(n_312),
.B2(n_310),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_289),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_350),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_329),
.C(n_275),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_289),
.Y(n_350)
);

XNOR2x2_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_282),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_294),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_353),
.A2(n_341),
.B(n_324),
.Y(n_380)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_276),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_360),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_276),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_SL g362 ( 
.A(n_331),
.B(n_290),
.C(n_294),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_363),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_327),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_298),
.C(n_293),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_315),
.B(n_305),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_370),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_314),
.B(n_293),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_285),
.C(n_326),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_294),
.B1(n_304),
.B2(n_282),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_313),
.B1(n_310),
.B2(n_319),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_373),
.A2(n_381),
.B1(n_384),
.B2(n_388),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_368),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_377),
.A2(n_393),
.B1(n_369),
.B2(n_352),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_385),
.B(n_386),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_334),
.B1(n_333),
.B2(n_337),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_333),
.C(n_339),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_389),
.C(n_391),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_338),
.B1(n_330),
.B2(n_308),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_332),
.B(n_308),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_353),
.A2(n_280),
.B(n_288),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_366),
.A2(n_288),
.B1(n_277),
.B2(n_281),
.Y(n_387)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_358),
.A2(n_277),
.B1(n_303),
.B2(n_213),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_259),
.C(n_208),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_351),
.A2(n_347),
.B(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_395),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_208),
.C(n_229),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_366),
.A2(n_213),
.B1(n_190),
.B2(n_164),
.Y(n_392)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_345),
.A2(n_213),
.B1(n_202),
.B2(n_154),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_202),
.C(n_264),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_397),
.C(n_355),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_202),
.B1(n_18),
.B2(n_260),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_197),
.C(n_133),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_400),
.A2(n_388),
.B1(n_384),
.B2(n_352),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_408),
.C(n_416),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_371),
.B(n_368),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_406),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_383),
.B(n_361),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_413),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_407),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_371),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_369),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_361),
.C(n_370),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_372),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_415),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_348),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_348),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_370),
.C(n_340),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_340),
.C(n_365),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_417),
.B(n_381),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_354),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_405),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_427),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_378),
.B(n_382),
.Y(n_422)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_422),
.Y(n_443)
);

FAx1_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_390),
.CI(n_378),
.CON(n_424),
.SN(n_424)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_428),
.Y(n_438)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_399),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_414),
.A2(n_380),
.B(n_385),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_418),
.A2(n_377),
.B1(n_379),
.B2(n_393),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_429),
.A2(n_408),
.B1(n_407),
.B2(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_432),
.Y(n_451)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_418),
.A2(n_379),
.B1(n_373),
.B2(n_404),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_436),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_398),
.C(n_402),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_424),
.C(n_422),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_398),
.C(n_416),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_442),
.B(n_444),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_417),
.C(n_397),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_429),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_448),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_396),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_446),
.B(n_450),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_386),
.C(n_354),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_396),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_437),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_355),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_436),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_457),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_456),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_426),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_451),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_443),
.A2(n_433),
.B(n_424),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_458),
.A2(n_461),
.B(n_463),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_464),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_449),
.A2(n_428),
.B(n_434),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_438),
.C(n_453),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_438),
.A2(n_440),
.B(n_448),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_466),
.A2(n_465),
.B(n_462),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_197),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_467),
.B(n_18),
.Y(n_471)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_468),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_470),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_464),
.B(n_243),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_175),
.C(n_46),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_472),
.B(n_8),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_465),
.A2(n_3),
.B1(n_8),
.B2(n_11),
.Y(n_473)
);

AOI322xp5_ASAP7_75t_L g478 ( 
.A1(n_473),
.A2(n_475),
.A3(n_457),
.B1(n_3),
.B2(n_8),
.C1(n_13),
.C2(n_2),
.Y(n_478)
);

OAI321xp33_ASAP7_75t_L g485 ( 
.A1(n_478),
.A2(n_483),
.A3(n_0),
.B1(n_1),
.B2(n_2),
.C(n_13),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_474),
.B1(n_472),
.B2(n_477),
.Y(n_484)
);

A2O1A1O1Ixp25_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_13),
.B(n_1),
.C(n_2),
.D(n_0),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_485),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_479),
.A2(n_469),
.B(n_470),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_486),
.B(n_482),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_480),
.C(n_1),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_488),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_490),
.B(n_0),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_0),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_1),
.B(n_2),
.Y(n_493)
);


endmodule