module fake_jpeg_19567_n_229 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_21),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_32),
.B1(n_20),
.B2(n_13),
.Y(n_38)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_30),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_31),
.B(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_28),
.B1(n_27),
.B2(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_29),
.B1(n_32),
.B2(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_38),
.B(n_40),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_27),
.B1(n_31),
.B2(n_20),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_33),
.B1(n_41),
.B2(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_19),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_51),
.B1(n_53),
.B2(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_13),
.B1(n_32),
.B2(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_71),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_44),
.B(n_49),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_48),
.B(n_43),
.Y(n_76)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_75),
.B1(n_34),
.B2(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_48),
.B1(n_55),
.B2(n_43),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_72),
.B1(n_61),
.B2(n_65),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_55),
.C(n_45),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_39),
.C(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_89),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_54),
.B(n_52),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_50),
.B(n_47),
.C(n_51),
.D(n_34),
.Y(n_86)
);

XOR2x2_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_76),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_61),
.B1(n_69),
.B2(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_74),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_94),
.B(n_98),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_11),
.B1(n_18),
.B2(n_46),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_106),
.B1(n_108),
.B2(n_77),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_58),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_17),
.B1(n_15),
.B2(n_18),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_72),
.B1(n_42),
.B2(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_57),
.B1(n_41),
.B2(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_78),
.C(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_118),
.C(n_120),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_86),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_125),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_78),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_96),
.C(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_39),
.C(n_79),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_126),
.B1(n_105),
.B2(n_93),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_77),
.B(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_109),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_41),
.B1(n_73),
.B2(n_67),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_39),
.C(n_73),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_46),
.C(n_67),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_108),
.B1(n_100),
.B2(n_102),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_46),
.C(n_23),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_145),
.B1(n_154),
.B2(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_103),
.B1(n_97),
.B2(n_46),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_97),
.B1(n_23),
.B2(n_16),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_12),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_0),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_124),
.B1(n_130),
.B2(n_112),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_115),
.B(n_12),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_12),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_23),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_120),
.C(n_127),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_162),
.C(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_131),
.C(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_147),
.B1(n_142),
.B2(n_156),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_117),
.A3(n_136),
.B1(n_23),
.B2(n_16),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_0),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_0),
.B(n_1),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_151),
.B(n_141),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_138),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_16),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_145),
.B(n_137),
.C(n_143),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_174),
.B(n_164),
.C(n_162),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_182),
.C(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_183),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_179),
.A2(n_180),
.B1(n_173),
.B2(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_148),
.C(n_16),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_1),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_9),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_196),
.C(n_9),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_192),
.B1(n_174),
.B2(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_161),
.B1(n_2),
.B2(n_3),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_161),
.B(n_2),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_3),
.C(n_4),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_195),
.B(n_4),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_1),
.C(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_201),
.C(n_205),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_202),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_3),
.C(n_4),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_201),
.B(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_5),
.B(n_6),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_190),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_213),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_189),
.C(n_6),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_209),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_6),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_215),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_212),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_217),
.B(n_7),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.B(n_221),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_220),
.B(n_6),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_8),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_8),
.Y(n_229)
);


endmodule