module fake_jpeg_4205_n_309 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_54),
.Y(n_104)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_19),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_64),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_32),
.Y(n_99)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_67),
.Y(n_103)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_83),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_64),
.B(n_60),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_32),
.B1(n_36),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_78),
.B1(n_92),
.B2(n_108),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_39),
.B1(n_26),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_68),
.B1(n_31),
.B2(n_25),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_27),
.B1(n_39),
.B2(n_26),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_106),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_99),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_39),
.B1(n_26),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_97),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_56),
.B(n_23),
.CI(n_41),
.CON(n_97),
.SN(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_45),
.A2(n_43),
.B1(n_25),
.B2(n_28),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_110),
.B1(n_1),
.B2(n_3),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_4),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_36),
.B1(n_29),
.B2(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_46),
.A2(n_29),
.B1(n_42),
.B2(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_23),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_23),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_146),
.B1(n_74),
.B2(n_107),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_123),
.Y(n_154)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_27),
.B1(n_39),
.B2(n_20),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_74),
.B1(n_82),
.B2(n_89),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_23),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_0),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_41),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_41),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_41),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_148),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_41),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_144),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_141),
.B1(n_147),
.B2(n_86),
.Y(n_155)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_147),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_78),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_97),
.A2(n_4),
.B(n_7),
.C(n_10),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_17),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_158),
.B1(n_121),
.B2(n_137),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_172),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_162),
.B1(n_169),
.B2(n_91),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_83),
.B1(n_70),
.B2(n_86),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_115),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_165),
.Y(n_210)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_92),
.B1(n_70),
.B2(n_109),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_81),
.C(n_85),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_181),
.C(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_85),
.C(n_69),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_114),
.C(n_113),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_129),
.B(n_125),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_204),
.C(n_167),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_113),
.B(n_142),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_193),
.B(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_118),
.B1(n_145),
.B2(n_69),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_214),
.B1(n_158),
.B2(n_180),
.Y(n_217)
);

BUFx8_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_118),
.B(n_122),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_135),
.B(n_140),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_143),
.C(n_122),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_197),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_148),
.C(n_136),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_199),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_82),
.B1(n_96),
.B2(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_203),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_131),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_171),
.C(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_164),
.B1(n_182),
.B2(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_140),
.B(n_138),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_121),
.B(n_75),
.Y(n_212)
);

OAI211xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_160),
.B(n_169),
.C(n_161),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_233),
.B1(n_200),
.B2(n_194),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_190),
.C(n_144),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_156),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_156),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_229),
.B(n_217),
.Y(n_247)
);

AOI221xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_193),
.B1(n_189),
.B2(n_195),
.C(n_212),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_163),
.A3(n_91),
.B1(n_75),
.B2(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_235),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_163),
.B1(n_133),
.B2(n_165),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_170),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_238),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_191),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_196),
.C(n_184),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_243),
.C(n_151),
.Y(n_273)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_245),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_218),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_202),
.C(n_185),
.Y(n_243)
);

AO221x1_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_205),
.B1(n_192),
.B2(n_190),
.C(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_225),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_207),
.B(n_209),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_216),
.B(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_200),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_224),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

OAI321xp33_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_214),
.A3(n_208),
.B1(n_194),
.B2(n_197),
.C(n_186),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_219),
.B(n_227),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_271),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_240),
.B(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_249),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_231),
.B1(n_216),
.B2(n_232),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_257),
.B1(n_248),
.B2(n_246),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_228),
.B1(n_229),
.B2(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_220),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_151),
.B1(n_192),
.B2(n_220),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_239),
.C(n_243),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_265),
.B(n_269),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_279),
.B(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_282),
.C(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_259),
.B(n_255),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_285),
.Y(n_291)
);

OAI22x1_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_247),
.B1(n_251),
.B2(n_256),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_260),
.B1(n_253),
.B2(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_245),
.C(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_260),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_246),
.C(n_250),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_292),
.C(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_288),
.B(n_289),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_262),
.B(n_259),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_255),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_252),
.C(n_241),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_290),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_280),
.B(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_12),
.B(n_14),
.Y(n_304)
);

OAI221xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_277),
.B1(n_284),
.B2(n_192),
.C(n_16),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_298),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.C(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_300),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_301),
.C(n_14),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_305),
.Y(n_309)
);


endmodule