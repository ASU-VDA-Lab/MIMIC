module fake_jpeg_23213_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx2_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_40),
.B1(n_19),
.B2(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_20),
.B1(n_26),
.B2(n_14),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_21),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_60),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_31),
.B2(n_41),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_45),
.B1(n_39),
.B2(n_44),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_0),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_64),
.B1(n_49),
.B2(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_66),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_50),
.B1(n_33),
.B2(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_83),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_75),
.B(n_64),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_48),
.B(n_39),
.C(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_51),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_91),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_97),
.B(n_21),
.Y(n_114)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_98),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_58),
.C(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_58),
.C(n_60),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_76),
.B(n_91),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_70),
.B1(n_75),
.B2(n_73),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_57),
.B1(n_95),
.B2(n_74),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_46),
.A3(n_81),
.B1(n_70),
.B2(n_15),
.C1(n_25),
.C2(n_7),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_97),
.C(n_86),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_123),
.C(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_124),
.B1(n_128),
.B2(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_47),
.C(n_55),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_15),
.B1(n_25),
.B2(n_22),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_24),
.C(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_136),
.B1(n_141),
.B2(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_114),
.B1(n_104),
.B2(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_123),
.B1(n_112),
.B2(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_128),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_116),
.C(n_126),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_13),
.C(n_3),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_106),
.B(n_118),
.C(n_105),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_16),
.B(n_14),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_100),
.B1(n_16),
.B2(n_14),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_1),
.C(n_2),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_2),
.C(n_3),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_1),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_130),
.B(n_136),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_143),
.B(n_148),
.Y(n_162)
);

OAI21x1_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_156),
.B(n_5),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_147),
.C(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_153),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_150),
.B(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_5),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_169),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_9),
.B(n_11),
.C(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_173),
.C(n_10),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);


endmodule