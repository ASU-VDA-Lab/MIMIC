module fake_jpeg_17859_n_294 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_294);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_23),
.B1(n_16),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_23),
.B1(n_25),
.B2(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_68),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_32),
.CI(n_27),
.CON(n_53),
.SN(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_15),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_13),
.CON(n_67),
.SN(n_67)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_16),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_13),
.B(n_1),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_45),
.C(n_47),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_81),
.Y(n_101)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_85),
.B1(n_23),
.B2(n_25),
.Y(n_100)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_16),
.B1(n_48),
.B2(n_25),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_55),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_54),
.B1(n_53),
.B2(n_51),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_100),
.B1(n_107),
.B2(n_89),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_55),
.C(n_61),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_18),
.C(n_21),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_79),
.B(n_75),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_101),
.B(n_105),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_110),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_16),
.B1(n_67),
.B2(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_64),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_74),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_123),
.B(n_21),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_87),
.B(n_70),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_117),
.B1(n_58),
.B2(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_74),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_60),
.B1(n_82),
.B2(n_76),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_121),
.B1(n_39),
.B2(n_44),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_82),
.B1(n_37),
.B2(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2x1p5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_45),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_18),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_132),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_52),
.B1(n_58),
.B2(n_77),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_96),
.B1(n_88),
.B2(n_72),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_21),
.A3(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_14),
.A3(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_28),
.CI(n_29),
.CON(n_132),
.SN(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_155),
.B1(n_129),
.B2(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_115),
.C(n_123),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_97),
.C(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_43),
.B1(n_108),
.B2(n_39),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_157),
.B1(n_158),
.B2(n_17),
.Y(n_174)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_159),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_122),
.B(n_116),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_131),
.B(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_93),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_160),
.B(n_22),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_118),
.B1(n_29),
.B2(n_28),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_83),
.C(n_93),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_114),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_124),
.B1(n_132),
.B2(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_18),
.C(n_17),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_0),
.B(n_2),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_167),
.B(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_129),
.B(n_130),
.Y(n_167)
);

AOI22x1_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_118),
.B1(n_62),
.B2(n_36),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_34),
.B(n_30),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_167),
.B(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_159),
.B1(n_36),
.B2(n_34),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_19),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_179)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_138),
.B1(n_143),
.B2(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_151),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_135),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_19),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_10),
.B(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_190),
.Y(n_226)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_197),
.B1(n_206),
.B2(n_208),
.Y(n_214)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_0),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_2),
.Y(n_225)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_181),
.C(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_181),
.C(n_182),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_166),
.C(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_169),
.B1(n_166),
.B2(n_171),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_187),
.B1(n_190),
.B2(n_199),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_177),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_196),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_173),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_193),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_169),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_224),
.A2(n_208),
.B1(n_196),
.B2(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_33),
.C(n_13),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_204),
.C(n_200),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_203),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_236),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_199),
.C(n_194),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_238),
.C(n_241),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_193),
.B1(n_205),
.B2(n_201),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_219),
.B1(n_214),
.B2(n_227),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_205),
.C(n_197),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_218),
.B1(n_212),
.B2(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_8),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_8),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_241),
.B(n_230),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_217),
.B(n_209),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_225),
.B(n_9),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_254),
.B1(n_236),
.B2(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_9),
.B1(n_11),
.B2(n_7),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

XOR2x1_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_9),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_228),
.B(n_11),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_249),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_19),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_268),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_3),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_5),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_255),
.C(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_251),
.C(n_19),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_5),
.B(n_6),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_259),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_268),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_270),
.C(n_271),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_267),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_282),
.B(n_269),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_264),
.B1(n_6),
.B2(n_5),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_18),
.C(n_19),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_278),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_290),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_288),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_33),
.C(n_13),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_13),
.B(n_134),
.Y(n_294)
);


endmodule