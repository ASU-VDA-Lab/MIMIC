module real_aes_12035_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_1932, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_1932;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_351;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1914;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1802;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_1496;
wire n_524;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1889;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_1352;
wire n_729;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1623 ( .A1(n_0), .A2(n_139), .B1(n_1578), .B2(n_1624), .C(n_1626), .Y(n_1623) );
AOI22xp5_ASAP7_75t_L g1612 ( .A1(n_1), .A2(n_123), .B1(n_1578), .B2(n_1582), .Y(n_1612) );
CKINVDCx5p33_ASAP7_75t_R g1476 ( .A(n_2), .Y(n_1476) );
INVx1_ASAP7_75t_L g759 ( .A(n_3), .Y(n_759) );
INVx1_ASAP7_75t_L g1477 ( .A(n_4), .Y(n_1477) );
INVx1_ASAP7_75t_L g869 ( .A(n_5), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g1466 ( .A1(n_6), .A2(n_91), .B1(n_604), .B2(n_1467), .C(n_1468), .Y(n_1466) );
INVx1_ASAP7_75t_L g1484 ( .A(n_6), .Y(n_1484) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_7), .A2(n_156), .B1(n_699), .B2(n_710), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_7), .A2(n_50), .B1(n_588), .B2(n_1312), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g1234 ( .A1(n_8), .A2(n_266), .B1(n_394), .B2(n_1002), .C(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1267 ( .A(n_8), .Y(n_1267) );
INVx1_ASAP7_75t_L g1627 ( .A(n_9), .Y(n_1627) );
INVx1_ASAP7_75t_L g1184 ( .A(n_10), .Y(n_1184) );
XNOR2x2_ASAP7_75t_L g1368 ( .A(n_11), .B(n_1369), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_12), .Y(n_1532) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_13), .A2(n_50), .B1(n_624), .B2(n_694), .Y(n_1376) );
AOI21xp33_ASAP7_75t_L g1397 ( .A1(n_13), .A2(n_601), .B(n_1059), .Y(n_1397) );
OAI22xp5_ASAP7_75t_L g1881 ( .A1(n_14), .A2(n_239), .B1(n_1191), .B2(n_1882), .Y(n_1881) );
CKINVDCx5p33_ASAP7_75t_R g1924 ( .A(n_14), .Y(n_1924) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_15), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_16), .A2(n_289), .B1(n_411), .B2(n_802), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g1217 ( .A(n_16), .Y(n_1217) );
INVxp33_ASAP7_75t_L g769 ( .A(n_17), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_17), .A2(n_73), .B1(n_701), .B2(n_818), .C(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g1846 ( .A(n_18), .Y(n_1846) );
AOI22xp33_ASAP7_75t_SL g1863 ( .A1(n_18), .A2(n_204), .B1(n_601), .B2(n_1061), .Y(n_1863) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_19), .A2(n_63), .B1(n_985), .B2(n_986), .C(n_987), .Y(n_984) );
INVx1_ASAP7_75t_L g1022 ( .A(n_19), .Y(n_1022) );
INVx1_ASAP7_75t_L g1388 ( .A(n_20), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_20), .A2(n_298), .B1(n_588), .B2(n_601), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_21), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_22), .A2(n_342), .B1(n_861), .B2(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1253 ( .A(n_22), .Y(n_1253) );
INVx1_ASAP7_75t_L g926 ( .A(n_23), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_23), .A2(n_48), .B1(n_969), .B2(n_970), .Y(n_968) );
INVxp67_ASAP7_75t_SL g1289 ( .A(n_24), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_24), .A2(n_325), .B1(n_393), .B2(n_399), .C(n_566), .Y(n_1308) );
INVxp33_ASAP7_75t_L g914 ( .A(n_25), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_25), .A2(n_77), .B1(n_588), .B2(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_26), .A2(n_329), .B1(n_794), .B2(n_796), .Y(n_793) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_26), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_27), .A2(n_230), .B1(n_399), .B2(n_1148), .C(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1495 ( .A(n_27), .Y(n_1495) );
OAI211xp5_ASAP7_75t_SL g1168 ( .A1(n_28), .A2(n_433), .B(n_1169), .C(n_1177), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1211 ( .A1(n_28), .A2(n_188), .B1(n_694), .B2(n_1212), .C(n_1214), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g1511 ( .A(n_29), .Y(n_1511) );
INVx1_ASAP7_75t_L g1005 ( .A(n_30), .Y(n_1005) );
INVx1_ASAP7_75t_L g350 ( .A(n_31), .Y(n_350) );
INVx1_ASAP7_75t_L g1241 ( .A(n_32), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_32), .A2(n_313), .B1(n_818), .B2(n_1262), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_33), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_34), .A2(n_192), .B1(n_516), .B2(n_921), .C(n_922), .Y(n_920) );
OAI33xp33_ASAP7_75t_L g960 ( .A1(n_34), .A2(n_192), .A3(n_418), .B1(n_578), .B2(n_787), .B3(n_1932), .Y(n_960) );
INVx1_ASAP7_75t_L g371 ( .A(n_35), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g1577 ( .A1(n_35), .A2(n_147), .B1(n_1578), .B2(n_1582), .Y(n_1577) );
INVx1_ASAP7_75t_L g1514 ( .A(n_36), .Y(n_1514) );
AOI221xp5_ASAP7_75t_L g1539 ( .A1(n_36), .A2(n_182), .B1(n_451), .B2(n_1540), .C(n_1542), .Y(n_1539) );
OAI221xp5_ASAP7_75t_L g1886 ( .A1(n_37), .A2(n_64), .B1(n_884), .B2(n_921), .C(n_922), .Y(n_1886) );
OAI222xp33_ASAP7_75t_L g1911 ( .A1(n_37), .A2(n_64), .B1(n_226), .B2(n_1004), .C1(n_1912), .C2(n_1913), .Y(n_1911) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_38), .A2(n_57), .B1(n_861), .B2(n_862), .Y(n_860) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_38), .A2(n_57), .B1(n_504), .B2(n_511), .C(n_884), .Y(n_883) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_39), .A2(n_591), .B(n_593), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_39), .A2(n_84), .B1(n_498), .B2(n_632), .C(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g778 ( .A(n_40), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_41), .A2(n_328), .B1(n_494), .B2(n_1127), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_41), .A2(n_248), .B1(n_563), .B2(n_1154), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1170 ( .A1(n_42), .A2(n_102), .B1(n_411), .B2(n_855), .Y(n_1170) );
AOI22xp33_ASAP7_75t_SL g1193 ( .A1(n_42), .A2(n_175), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_43), .A2(n_199), .B1(n_855), .B2(n_856), .C(n_1176), .Y(n_1175) );
OAI21xp33_ASAP7_75t_SL g1190 ( .A1(n_43), .A2(n_1191), .B(n_1192), .Y(n_1190) );
INVx1_ASAP7_75t_L g1248 ( .A(n_44), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_44), .A2(n_318), .B1(n_1194), .B2(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1851 ( .A1(n_45), .A2(n_201), .B1(n_488), .B2(n_1122), .Y(n_1851) );
AOI22xp33_ASAP7_75t_L g1856 ( .A1(n_45), .A2(n_201), .B1(n_1451), .B2(n_1467), .Y(n_1856) );
OAI222xp33_ASAP7_75t_L g1337 ( .A1(n_46), .A2(n_171), .B1(n_270), .B2(n_1338), .C1(n_1340), .C2(n_1341), .Y(n_1337) );
AOI221xp5_ASAP7_75t_L g1362 ( .A1(n_46), .A2(n_171), .B1(n_1363), .B2(n_1364), .C(n_1366), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g1373 ( .A(n_47), .Y(n_1373) );
INVx1_ASAP7_75t_L g932 ( .A(n_48), .Y(n_932) );
INVxp67_ASAP7_75t_SL g1288 ( .A(n_49), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_49), .A2(n_213), .B1(n_858), .B2(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g938 ( .A(n_51), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1895 ( .A(n_52), .Y(n_1895) );
AO221x2_ASAP7_75t_L g1710 ( .A1(n_53), .A2(n_263), .B1(n_1624), .B2(n_1711), .C(n_1713), .Y(n_1710) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_54), .A2(n_200), .B1(n_411), .B2(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_54), .A2(n_200), .B1(n_844), .B2(n_845), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_55), .A2(n_93), .B1(n_393), .B2(n_394), .C(n_399), .Y(n_392) );
INVxp67_ASAP7_75t_L g539 ( .A(n_55), .Y(n_539) );
INVxp67_ASAP7_75t_L g1410 ( .A(n_56), .Y(n_1410) );
INVx1_ASAP7_75t_L g1117 ( .A(n_58), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_59), .A2(n_154), .B1(n_1013), .B2(n_1122), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_59), .A2(n_217), .B1(n_1130), .B2(n_1131), .C(n_1133), .Y(n_1129) );
XNOR2xp5_ASAP7_75t_L g1876 ( .A(n_60), .B(n_1877), .Y(n_1876) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_61), .A2(n_143), .B1(n_570), .B2(n_578), .C(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g639 ( .A(n_61), .Y(n_639) );
INVxp67_ASAP7_75t_L g1429 ( .A(n_62), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_62), .A2(n_99), .B1(n_603), .B2(n_1130), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_63), .A2(n_207), .B1(n_1017), .B2(n_1019), .C(n_1021), .Y(n_1016) );
INVx1_ASAP7_75t_L g909 ( .A(n_65), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_65), .A2(n_290), .B1(n_1578), .B2(n_1582), .Y(n_1585) );
AOI22xp5_ASAP7_75t_L g1611 ( .A1(n_66), .A2(n_324), .B1(n_1566), .B2(n_1574), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_67), .Y(n_1529) );
CKINVDCx5p33_ASAP7_75t_R g1893 ( .A(n_68), .Y(n_1893) );
AOI21xp33_ASAP7_75t_L g1047 ( .A1(n_69), .A2(n_406), .B(n_856), .Y(n_1047) );
INVxp33_ASAP7_75t_L g1073 ( .A(n_69), .Y(n_1073) );
XOR2x2_ASAP7_75t_L g754 ( .A(n_70), .B(n_755), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g1470 ( .A1(n_71), .A2(n_214), .B1(n_1317), .B2(n_1447), .Y(n_1470) );
OAI221xp5_ASAP7_75t_L g1489 ( .A1(n_71), .A2(n_214), .B1(n_922), .B2(n_1282), .C(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g431 ( .A(n_72), .Y(n_431) );
INVxp33_ASAP7_75t_L g773 ( .A(n_73), .Y(n_773) );
INVxp33_ASAP7_75t_L g917 ( .A(n_74), .Y(n_917) );
AOI21xp33_ASAP7_75t_L g955 ( .A1(n_74), .A2(n_603), .B(n_604), .Y(n_955) );
INVx1_ASAP7_75t_L g1434 ( .A(n_75), .Y(n_1434) );
AOI22x1_ASAP7_75t_L g1165 ( .A1(n_76), .A2(n_1166), .B1(n_1218), .B2(n_1219), .Y(n_1165) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_76), .Y(n_1218) );
AO22x1_ASAP7_75t_L g1588 ( .A1(n_76), .A2(n_252), .B1(n_1582), .B2(n_1589), .Y(n_1588) );
INVxp33_ASAP7_75t_L g918 ( .A(n_77), .Y(n_918) );
INVx1_ASAP7_75t_L g1109 ( .A(n_78), .Y(n_1109) );
AO22x1_ASAP7_75t_L g1590 ( .A1(n_79), .A2(n_249), .B1(n_1566), .B2(n_1574), .Y(n_1590) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_80), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_81), .Y(n_1386) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_82), .A2(n_332), .B1(n_854), .B2(n_855), .C(n_856), .Y(n_853) );
INVxp33_ASAP7_75t_L g879 ( .A(n_82), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_83), .A2(n_177), .B1(n_632), .B2(n_1378), .Y(n_1377) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_83), .A2(n_177), .B1(n_750), .B2(n_1141), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_84), .A2(n_234), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_85), .A2(n_176), .B1(n_795), .B2(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1030 ( .A(n_85), .Y(n_1030) );
OAI221xp5_ASAP7_75t_L g1515 ( .A1(n_86), .A2(n_159), .B1(n_511), .B2(n_515), .C(n_921), .Y(n_1515) );
OAI22xp33_ASAP7_75t_L g1537 ( .A1(n_86), .A2(n_159), .B1(n_1233), .B2(n_1538), .Y(n_1537) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_87), .A2(n_291), .B1(n_451), .B2(n_868), .Y(n_867) );
INVxp67_ASAP7_75t_SL g897 ( .A(n_87), .Y(n_897) );
INVx1_ASAP7_75t_L g1319 ( .A(n_88), .Y(n_1319) );
AOI22xp33_ASAP7_75t_SL g857 ( .A1(n_89), .A2(n_224), .B1(n_447), .B2(n_858), .Y(n_857) );
INVxp33_ASAP7_75t_SL g882 ( .A(n_89), .Y(n_882) );
BUFx2_ASAP7_75t_L g378 ( .A(n_90), .Y(n_378) );
OR2x2_ASAP7_75t_L g467 ( .A(n_90), .B(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g471 ( .A(n_90), .Y(n_471) );
INVx1_ASAP7_75t_L g483 ( .A(n_90), .Y(n_483) );
INVx1_ASAP7_75t_L g1486 ( .A(n_91), .Y(n_1486) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_92), .A2(n_294), .B1(n_494), .B2(n_519), .C(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g738 ( .A(n_92), .Y(n_738) );
INVxp33_ASAP7_75t_SL g531 ( .A(n_93), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g1379 ( .A1(n_94), .A2(n_109), .B1(n_699), .B2(n_710), .Y(n_1379) );
INVx1_ASAP7_75t_L g1405 ( .A(n_94), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_95), .Y(n_1036) );
INVx1_ASAP7_75t_L g1813 ( .A(n_96), .Y(n_1813) );
AOI22xp33_ASAP7_75t_L g1853 ( .A1(n_96), .A2(n_335), .B1(n_498), .B2(n_632), .Y(n_1853) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_97), .A2(n_227), .B1(n_1052), .B2(n_1054), .C(n_1057), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1083 ( .A(n_97), .Y(n_1083) );
AOI221xp5_ASAP7_75t_SL g993 ( .A1(n_98), .A2(n_103), .B1(n_856), .B2(n_994), .C(n_996), .Y(n_993) );
INVx1_ASAP7_75t_L g1012 ( .A(n_98), .Y(n_1012) );
INVxp33_ASAP7_75t_L g1423 ( .A(n_99), .Y(n_1423) );
INVx1_ASAP7_75t_L g989 ( .A(n_100), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g1505 ( .A1(n_101), .A2(n_1506), .B1(n_1553), .B2(n_1554), .Y(n_1505) );
INVx1_ASAP7_75t_L g1553 ( .A(n_101), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_102), .A2(n_119), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g1011 ( .A(n_103), .Y(n_1011) );
XOR2x2_ASAP7_75t_L g558 ( .A(n_104), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g453 ( .A(n_105), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_106), .Y(n_721) );
INVxp67_ASAP7_75t_SL g933 ( .A(n_107), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_107), .A2(n_300), .B1(n_593), .B2(n_965), .C(n_967), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1818 ( .A1(n_108), .A2(n_115), .B1(n_1819), .B2(n_1822), .Y(n_1818) );
OAI22xp5_ASAP7_75t_L g1830 ( .A1(n_108), .A2(n_115), .B1(n_1831), .B2(n_1833), .Y(n_1830) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_109), .B(n_427), .Y(n_1391) );
AO221x1_ASAP7_75t_L g1595 ( .A1(n_110), .A2(n_126), .B1(n_1578), .B2(n_1582), .C(n_1596), .Y(n_1595) );
OAI22xp5_ASAP7_75t_L g1883 ( .A1(n_111), .A2(n_226), .B1(n_466), .B2(n_1884), .Y(n_1883) );
CKINVDCx5p33_ASAP7_75t_R g1922 ( .A(n_111), .Y(n_1922) );
AO221x1_ASAP7_75t_L g1603 ( .A1(n_112), .A2(n_314), .B1(n_1578), .B2(n_1582), .C(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1606 ( .A(n_113), .Y(n_1606) );
INVx1_ASAP7_75t_L g1440 ( .A(n_114), .Y(n_1440) );
INVxp67_ASAP7_75t_L g1419 ( .A(n_116), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_116), .A2(n_149), .B1(n_954), .B2(n_1002), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_117), .A2(n_259), .B1(n_413), .B2(n_601), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_117), .A2(n_606), .B(n_608), .C(n_614), .Y(n_605) );
INVx1_ASAP7_75t_L g659 ( .A(n_118), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_118), .A2(n_136), .B1(n_498), .B2(n_694), .C(n_695), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g1171 ( .A1(n_119), .A2(n_175), .B1(n_393), .B2(n_1172), .C(n_1173), .Y(n_1171) );
INVx1_ASAP7_75t_L g1456 ( .A(n_120), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1465 ( .A(n_121), .Y(n_1465) );
INVx1_ASAP7_75t_L g1600 ( .A(n_122), .Y(n_1600) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_124), .A2(n_186), .B1(n_393), .B2(n_399), .C(n_1000), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_124), .A2(n_176), .B1(n_1026), .B2(n_1028), .C(n_1029), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g1565 ( .A1(n_125), .A2(n_153), .B1(n_1566), .B2(n_1574), .Y(n_1565) );
INVx1_ASAP7_75t_L g1151 ( .A(n_127), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g1531 ( .A(n_128), .Y(n_1531) );
OAI222xp33_ASAP7_75t_L g1342 ( .A1(n_129), .A2(n_195), .B1(n_327), .B2(n_1004), .C1(n_1317), .C2(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1354 ( .A(n_129), .Y(n_1354) );
INVx1_ASAP7_75t_L g1714 ( .A(n_130), .Y(n_1714) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_131), .A2(n_308), .B1(n_568), .B2(n_570), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_131), .A2(n_184), .B1(n_626), .B2(n_628), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_132), .A2(n_303), .B1(n_1059), .B2(n_1172), .C(n_1243), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_132), .A2(n_221), .B1(n_901), .B2(n_1194), .Y(n_1257) );
INVxp67_ASAP7_75t_L g1418 ( .A(n_133), .Y(n_1418) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_133), .A2(n_189), .B1(n_406), .B2(n_854), .C(n_856), .Y(n_1444) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_134), .A2(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g615 ( .A(n_134), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_135), .A2(n_184), .B1(n_563), .B2(n_565), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_135), .A2(n_308), .B1(n_478), .B2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g680 ( .A(n_136), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_137), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_138), .A2(n_169), .B1(n_504), .B2(n_512), .C(n_1282), .Y(n_1281) );
OAI22xp33_ASAP7_75t_L g1316 ( .A1(n_138), .A2(n_169), .B1(n_1041), .B2(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1111 ( .A(n_140), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_141), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g1420 ( .A1(n_142), .A2(n_180), .B1(n_884), .B2(n_921), .C(n_922), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_142), .A2(n_180), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
INVx1_ASAP7_75t_L g610 ( .A(n_143), .Y(n_610) );
INVx1_ASAP7_75t_L g991 ( .A(n_144), .Y(n_991) );
AOI221xp5_ASAP7_75t_L g1329 ( .A1(n_145), .A2(n_299), .B1(n_1059), .B2(n_1148), .C(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1361 ( .A(n_145), .Y(n_1361) );
CKINVDCx5p33_ASAP7_75t_R g1898 ( .A(n_146), .Y(n_1898) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_148), .Y(n_1534) );
INVxp67_ASAP7_75t_L g1415 ( .A(n_149), .Y(n_1415) );
INVx1_ASAP7_75t_L g1570 ( .A(n_150), .Y(n_1570) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_151), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g1811 ( .A(n_152), .Y(n_1811) );
INVx1_ASAP7_75t_L g1136 ( .A(n_154), .Y(n_1136) );
INVx1_ASAP7_75t_L g1605 ( .A(n_155), .Y(n_1605) );
INVx1_ASAP7_75t_L g1394 ( .A(n_156), .Y(n_1394) );
INVx1_ASAP7_75t_L g915 ( .A(n_157), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_157), .B(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g784 ( .A(n_158), .Y(n_784) );
INVx1_ASAP7_75t_L g1571 ( .A(n_160), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_160), .B(n_1569), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_161), .A2(n_243), .B1(n_447), .B2(n_451), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_161), .A2(n_243), .B1(n_815), .B2(n_1009), .C(n_1010), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_162), .A2(n_190), .B1(n_741), .B2(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_SL g829 ( .A(n_162), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_163), .A2(n_221), .B1(n_455), .B2(n_1245), .Y(n_1244) );
AOI22xp33_ASAP7_75t_SL g1255 ( .A1(n_163), .A2(n_303), .B1(n_626), .B2(n_1256), .Y(n_1255) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_164), .A2(n_406), .B(n_458), .Y(n_1237) );
INVx1_ASAP7_75t_L g1266 ( .A(n_164), .Y(n_1266) );
INVx2_ASAP7_75t_L g362 ( .A(n_165), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_166), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_167), .A2(n_319), .B1(n_399), .B2(n_448), .C(n_865), .Y(n_864) );
INVxp33_ASAP7_75t_SL g890 ( .A(n_167), .Y(n_890) );
BUFx3_ASAP7_75t_L g386 ( .A(n_168), .Y(n_386) );
INVx1_ASAP7_75t_L g415 ( .A(n_168), .Y(n_415) );
INVx1_ASAP7_75t_L g1178 ( .A(n_170), .Y(n_1178) );
INVx1_ASAP7_75t_L g1518 ( .A(n_172), .Y(n_1518) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_172), .A2(n_282), .B1(n_796), .B2(n_969), .Y(n_1550) );
AOI22xp33_ASAP7_75t_SL g1850 ( .A1(n_173), .A2(n_241), .B1(n_632), .B2(n_1378), .Y(n_1850) );
AOI22xp33_ASAP7_75t_SL g1857 ( .A1(n_173), .A2(n_241), .B1(n_413), .B2(n_601), .Y(n_1857) );
INVx1_ASAP7_75t_L g764 ( .A(n_174), .Y(n_764) );
INVx1_ASAP7_75t_L g940 ( .A(n_178), .Y(n_940) );
INVxp33_ASAP7_75t_L g1279 ( .A(n_179), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g1314 ( .A1(n_179), .A2(n_225), .B1(n_603), .B2(n_604), .C(n_1148), .Y(n_1314) );
INVx1_ASAP7_75t_L g1809 ( .A(n_181), .Y(n_1809) );
AOI22xp33_ASAP7_75t_L g1854 ( .A1(n_181), .A2(n_297), .B1(n_488), .B2(n_1122), .Y(n_1854) );
INVx1_ASAP7_75t_L g1510 ( .A(n_182), .Y(n_1510) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_183), .A2(n_311), .B1(n_541), .B2(n_624), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_183), .A2(n_311), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_185), .Y(n_463) );
INVx1_ASAP7_75t_L g1031 ( .A(n_186), .Y(n_1031) );
OAI221xp5_ASAP7_75t_SL g1040 ( .A1(n_187), .A2(n_331), .B1(n_862), .B2(n_1041), .C(n_1043), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1075 ( .A1(n_187), .A2(n_331), .B1(n_512), .B2(n_515), .C(n_921), .Y(n_1075) );
INVxp67_ASAP7_75t_SL g1179 ( .A(n_188), .Y(n_1179) );
INVxp67_ASAP7_75t_L g1416 ( .A(n_189), .Y(n_1416) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_190), .Y(n_837) );
INVx1_ASAP7_75t_L g990 ( .A(n_191), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g1896 ( .A(n_193), .Y(n_1896) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_194), .Y(n_808) );
INVx1_ASAP7_75t_L g1347 ( .A(n_195), .Y(n_1347) );
INVxp33_ASAP7_75t_SL g1104 ( .A(n_196), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1139 ( .A1(n_196), .A2(n_253), .B1(n_1130), .B2(n_1140), .C(n_1142), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_197), .A2(n_287), .B1(n_802), .B2(n_1245), .Y(n_1328) );
INVx1_ASAP7_75t_L g1352 ( .A(n_197), .Y(n_1352) );
INVx1_ASAP7_75t_L g1628 ( .A(n_198), .Y(n_1628) );
INVxp33_ASAP7_75t_SL g1208 ( .A(n_199), .Y(n_1208) );
INVx1_ASAP7_75t_L g1716 ( .A(n_202), .Y(n_1716) );
INVx1_ASAP7_75t_L g1064 ( .A(n_203), .Y(n_1064) );
INVx1_ASAP7_75t_L g1839 ( .A(n_204), .Y(n_1839) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_205), .A2(n_305), .B1(n_393), .B2(n_455), .C(n_458), .Y(n_454) );
INVxp33_ASAP7_75t_SL g492 ( .A(n_205), .Y(n_492) );
INVx1_ASAP7_75t_L g390 ( .A(n_206), .Y(n_390) );
INVx1_ASAP7_75t_L g402 ( .A(n_206), .Y(n_402) );
INVx1_ASAP7_75t_L g988 ( .A(n_207), .Y(n_988) );
INVxp33_ASAP7_75t_SL g1276 ( .A(n_208), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_208), .A2(n_215), .B1(n_1000), .B2(n_1155), .Y(n_1315) );
INVx1_ASAP7_75t_L g669 ( .A(n_209), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_209), .A2(n_233), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g937 ( .A(n_210), .Y(n_937) );
INVx1_ASAP7_75t_L g436 ( .A(n_211), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_211), .A2(n_245), .B1(n_504), .B2(n_511), .C(n_515), .Y(n_503) );
INVx1_ASAP7_75t_L g859 ( .A(n_212), .Y(n_859) );
INVx1_ASAP7_75t_L g1293 ( .A(n_213), .Y(n_1293) );
INVxp33_ASAP7_75t_SL g1280 ( .A(n_215), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_216), .Y(n_597) );
INVx1_ASAP7_75t_L g1120 ( .A(n_217), .Y(n_1120) );
INVx1_ASAP7_75t_L g1597 ( .A(n_218), .Y(n_1597) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_219), .A2(n_279), .B1(n_791), .B2(n_799), .Y(n_798) );
OAI211xp5_ASAP7_75t_SL g812 ( .A1(n_219), .A2(n_813), .B(n_814), .C(n_820), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g1586 ( .A1(n_220), .A2(n_343), .B1(n_1566), .B2(n_1574), .Y(n_1586) );
INVx1_ASAP7_75t_L g1269 ( .A(n_222), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_223), .A2(n_306), .B1(n_856), .B2(n_994), .C(n_996), .Y(n_1327) );
INVx1_ASAP7_75t_L g1350 ( .A(n_223), .Y(n_1350) );
INVxp33_ASAP7_75t_L g877 ( .A(n_224), .Y(n_877) );
INVxp33_ASAP7_75t_L g1277 ( .A(n_225), .Y(n_1277) );
INVx1_ASAP7_75t_L g1080 ( .A(n_227), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_228), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_229), .A2(n_235), .B1(n_742), .B2(n_1172), .Y(n_1469) );
INVx1_ASAP7_75t_L g1482 ( .A(n_229), .Y(n_1482) );
INVx1_ASAP7_75t_L g1497 ( .A(n_230), .Y(n_1497) );
INVxp67_ASAP7_75t_L g1426 ( .A(n_231), .Y(n_1426) );
AOI221xp5_ASAP7_75t_L g1450 ( .A1(n_231), .A2(n_244), .B1(n_396), .B2(n_1451), .C(n_1452), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_232), .A2(n_292), .B1(n_405), .B2(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1079 ( .A(n_232), .Y(n_1079) );
INVx1_ASAP7_75t_L g674 ( .A(n_233), .Y(n_674) );
INVx1_ASAP7_75t_L g634 ( .A(n_234), .Y(n_634) );
INVx1_ASAP7_75t_L g1487 ( .A(n_235), .Y(n_1487) );
XNOR2xp5_ASAP7_75t_L g1457 ( .A(n_236), .B(n_1458), .Y(n_1457) );
OAI211xp5_ASAP7_75t_SL g1180 ( .A1(n_237), .A2(n_1181), .B(n_1182), .C(n_1187), .Y(n_1180) );
INVx1_ASAP7_75t_L g1215 ( .A(n_237), .Y(n_1215) );
INVx1_ASAP7_75t_L g1389 ( .A(n_238), .Y(n_1389) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_238), .A2(n_1004), .B(n_1404), .C(n_1407), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g1921 ( .A(n_239), .Y(n_1921) );
CKINVDCx5p33_ASAP7_75t_R g1899 ( .A(n_240), .Y(n_1899) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_242), .A2(n_285), .B1(n_405), .B2(n_411), .Y(n_404) );
INVxp67_ASAP7_75t_L g524 ( .A(n_242), .Y(n_524) );
INVxp33_ASAP7_75t_L g1424 ( .A(n_244), .Y(n_1424) );
INVx1_ASAP7_75t_L g441 ( .A(n_245), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_246), .A2(n_256), .B1(n_396), .B2(n_413), .Y(n_1046) );
INVxp33_ASAP7_75t_L g1074 ( .A(n_246), .Y(n_1074) );
INVx1_ASAP7_75t_L g1523 ( .A(n_247), .Y(n_1523) );
AOI221xp5_ASAP7_75t_L g1546 ( .A1(n_247), .A2(n_261), .B1(n_591), .B2(n_1452), .C(n_1547), .Y(n_1546) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_248), .Y(n_1125) );
XNOR2x1_ASAP7_75t_L g1323 ( .A(n_250), .B(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g425 ( .A(n_251), .Y(n_425) );
INVxp33_ASAP7_75t_SL g1108 ( .A(n_253), .Y(n_1108) );
BUFx3_ASAP7_75t_L g387 ( .A(n_254), .Y(n_387) );
INVx1_ASAP7_75t_L g398 ( .A(n_254), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g1892 ( .A(n_255), .Y(n_1892) );
INVxp33_ASAP7_75t_L g1070 ( .A(n_256), .Y(n_1070) );
INVx1_ASAP7_75t_L g1094 ( .A(n_257), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_258), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_258), .B(n_323), .Y(n_468) );
AND2x2_ASAP7_75t_L g484 ( .A(n_258), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g556 ( .A(n_258), .Y(n_556) );
INVx1_ASAP7_75t_L g618 ( .A(n_259), .Y(n_618) );
OAI332xp33_ASAP7_75t_L g1887 ( .A1(n_260), .A2(n_518), .A3(n_552), .B1(n_1888), .B2(n_1891), .B3(n_1894), .C1(n_1897), .C2(n_1900), .Y(n_1887) );
INVx1_ASAP7_75t_L g1925 ( .A(n_260), .Y(n_1925) );
INVx1_ASAP7_75t_L g1521 ( .A(n_261), .Y(n_1521) );
INVx1_ASAP7_75t_L g871 ( .A(n_262), .Y(n_871) );
INVx1_ASAP7_75t_L g1150 ( .A(n_264), .Y(n_1150) );
OR2x2_ASAP7_75t_L g389 ( .A(n_265), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g403 ( .A(n_265), .Y(n_403) );
INVx1_ASAP7_75t_L g1264 ( .A(n_266), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g1890 ( .A(n_267), .Y(n_1890) );
INVx1_ASAP7_75t_L g1432 ( .A(n_268), .Y(n_1432) );
INVx1_ASAP7_75t_L g461 ( .A(n_269), .Y(n_461) );
INVx1_ASAP7_75t_L g1367 ( .A(n_270), .Y(n_1367) );
CKINVDCx16_ASAP7_75t_R g980 ( .A(n_271), .Y(n_980) );
INVx1_ASAP7_75t_L g1296 ( .A(n_272), .Y(n_1296) );
INVx1_ASAP7_75t_L g1249 ( .A(n_273), .Y(n_1249) );
INVx1_ASAP7_75t_L g872 ( .A(n_274), .Y(n_872) );
INVxp67_ASAP7_75t_SL g1183 ( .A(n_275), .Y(n_1183) );
OAI211xp5_ASAP7_75t_SL g1201 ( .A1(n_275), .A2(n_928), .B(n_1202), .C(n_1205), .Y(n_1201) );
INVx1_ASAP7_75t_L g391 ( .A(n_276), .Y(n_391) );
INVx1_ASAP7_75t_L g726 ( .A(n_277), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_277), .A2(n_304), .B1(n_741), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g1050 ( .A(n_278), .Y(n_1050) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_279), .A2(n_825), .B1(n_826), .B2(n_833), .C(n_842), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_280), .A2(n_301), .B1(n_858), .B2(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1360 ( .A(n_280), .Y(n_1360) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_281), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g1526 ( .A(n_282), .Y(n_1526) );
INVx1_ASAP7_75t_L g449 ( .A(n_283), .Y(n_449) );
INVx1_ASAP7_75t_L g907 ( .A(n_284), .Y(n_907) );
INVxp67_ASAP7_75t_L g543 ( .A(n_285), .Y(n_543) );
INVx1_ASAP7_75t_L g1382 ( .A(n_286), .Y(n_1382) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_286), .A2(n_587), .B(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1349 ( .A(n_287), .Y(n_1349) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_288), .Y(n_1513) );
INVxp33_ASAP7_75t_L g1209 ( .A(n_289), .Y(n_1209) );
INVxp33_ASAP7_75t_L g887 ( .A(n_291), .Y(n_887) );
INVx1_ASAP7_75t_L g1086 ( .A(n_292), .Y(n_1086) );
INVx1_ASAP7_75t_L g1836 ( .A(n_293), .Y(n_1836) );
AOI22xp33_ASAP7_75t_L g1862 ( .A1(n_293), .A2(n_326), .B1(n_792), .B2(n_1467), .Y(n_1862) );
INVx1_ASAP7_75t_L g739 ( .A(n_294), .Y(n_739) );
INVx1_ASAP7_75t_L g942 ( .A(n_295), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_296), .Y(n_1528) );
INVx1_ASAP7_75t_L g1817 ( .A(n_297), .Y(n_1817) );
INVx1_ASAP7_75t_L g1385 ( .A(n_298), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_299), .A2(n_301), .B1(n_1017), .B2(n_1358), .C(n_1359), .Y(n_1357) );
INVxp33_ASAP7_75t_L g927 ( .A(n_300), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_302), .A2(n_333), .B1(n_855), .B2(n_1155), .Y(n_1474) );
INVx1_ASAP7_75t_L g1499 ( .A(n_302), .Y(n_1499) );
INVx1_ASAP7_75t_L g724 ( .A(n_304), .Y(n_724) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_305), .Y(n_486) );
INVx1_ASAP7_75t_L g1356 ( .A(n_306), .Y(n_1356) );
CKINVDCx5p33_ASAP7_75t_R g1336 ( .A(n_307), .Y(n_1336) );
INVx1_ASAP7_75t_L g1439 ( .A(n_309), .Y(n_1439) );
INVx1_ASAP7_75t_L g873 ( .A(n_310), .Y(n_873) );
INVx1_ASAP7_75t_L g1044 ( .A(n_312), .Y(n_1044) );
INVx1_ASAP7_75t_L g1247 ( .A(n_313), .Y(n_1247) );
INVx1_ASAP7_75t_L g1271 ( .A(n_314), .Y(n_1271) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_315), .B(n_350), .Y(n_1573) );
AND3x2_ASAP7_75t_L g1581 ( .A(n_315), .B(n_350), .C(n_1570), .Y(n_1581) );
INVx2_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
XNOR2x2_ASAP7_75t_L g1100 ( .A(n_317), .B(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1231 ( .A(n_318), .Y(n_1231) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_319), .Y(n_893) );
INVx1_ASAP7_75t_L g1106 ( .A(n_320), .Y(n_1106) );
CKINVDCx5p33_ASAP7_75t_R g1889 ( .A(n_321), .Y(n_1889) );
INVx1_ASAP7_75t_L g1299 ( .A(n_322), .Y(n_1299) );
INVx1_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
INVx2_ASAP7_75t_L g485 ( .A(n_323), .Y(n_485) );
XNOR2xp5_ASAP7_75t_L g1805 ( .A(n_324), .B(n_1806), .Y(n_1805) );
AOI22xp33_ASAP7_75t_L g1871 ( .A1(n_324), .A2(n_1872), .B1(n_1875), .B2(n_1927), .Y(n_1871) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_325), .Y(n_1292) );
INVx1_ASAP7_75t_L g1826 ( .A(n_326), .Y(n_1826) );
INVx1_ASAP7_75t_L g1346 ( .A(n_327), .Y(n_1346) );
OAI22xp33_ASAP7_75t_L g1156 ( .A1(n_328), .A2(n_337), .B1(n_395), .B2(n_570), .Y(n_1156) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_329), .Y(n_841) );
INVx1_ASAP7_75t_L g1297 ( .A(n_330), .Y(n_1297) );
INVxp33_ASAP7_75t_L g881 ( .A(n_332), .Y(n_881) );
INVx1_ASAP7_75t_L g1494 ( .A(n_333), .Y(n_1494) );
INVx1_ASAP7_75t_L g1185 ( .A(n_334), .Y(n_1185) );
INVx1_ASAP7_75t_L g1814 ( .A(n_335), .Y(n_1814) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_336), .Y(n_1463) );
INVxp67_ASAP7_75t_SL g1124 ( .A(n_337), .Y(n_1124) );
INVx1_ASAP7_75t_L g677 ( .A(n_338), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_338), .A2(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g1063 ( .A(n_339), .Y(n_1063) );
INVx1_ASAP7_75t_L g1300 ( .A(n_340), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_341), .Y(n_1236) );
INVx1_ASAP7_75t_L g1252 ( .A(n_342), .Y(n_1252) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_366), .B(n_1557), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
AND2x4_ASAP7_75t_L g1870 ( .A(n_348), .B(n_354), .Y(n_1870) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_SL g1874 ( .A(n_349), .Y(n_1874) );
NAND2xp5_ASAP7_75t_L g1930 ( .A(n_349), .B(n_351), .Y(n_1930) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g1873 ( .A(n_351), .B(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_356), .B(n_471), .Y(n_1847) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g630 ( .A(n_357), .B(n_365), .Y(n_630) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g519 ( .A(n_358), .B(n_520), .Y(n_519) );
INVx8_ASAP7_75t_L g1835 ( .A(n_359), .Y(n_1835) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
OR2x2_ASAP7_75t_L g466 ( .A(n_360), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g523 ( .A(n_360), .Y(n_523) );
INVx2_ASAP7_75t_SL g548 ( .A(n_360), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_360), .A2(n_527), .B1(n_583), .B2(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_360), .Y(n_889) );
INVx2_ASAP7_75t_SL g931 ( .A(n_360), .Y(n_931) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_360), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_360), .A2(n_527), .B1(n_1336), .B2(n_1367), .Y(n_1366) );
OR2x6_ASAP7_75t_L g1842 ( .A(n_360), .B(n_1838), .Y(n_1842) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x4_ASAP7_75t_L g480 ( .A(n_362), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g490 ( .A(n_362), .Y(n_490) );
AND2x2_ASAP7_75t_L g496 ( .A(n_362), .B(n_363), .Y(n_496) );
INVx2_ASAP7_75t_L g500 ( .A(n_362), .Y(n_500) );
INVx1_ASAP7_75t_L g530 ( .A(n_362), .Y(n_530) );
INVx2_ASAP7_75t_L g481 ( .A(n_363), .Y(n_481) );
INVx1_ASAP7_75t_L g502 ( .A(n_363), .Y(n_502) );
INVx1_ASAP7_75t_L g509 ( .A(n_363), .Y(n_509) );
INVx1_ASAP7_75t_L g529 ( .A(n_363), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_363), .B(n_500), .Y(n_538) );
AND2x4_ASAP7_75t_L g1832 ( .A(n_364), .B(n_509), .Y(n_1832) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g1833 ( .A(n_365), .B(n_613), .Y(n_1833) );
XNOR2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_751), .Y(n_366) );
XNOR2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_643), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_557), .B1(n_558), .B2(n_642), .Y(n_369) );
INVx1_ASAP7_75t_SL g642 ( .A(n_370), .Y(n_642) );
XNOR2x1_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_473), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_379), .B1(n_463), .B2(n_464), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI31xp33_ASAP7_75t_SL g982 ( .A1(n_375), .A2(n_983), .A3(n_992), .B(n_998), .Y(n_982) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g559 ( .A1(n_376), .A2(n_560), .B(n_605), .C(n_621), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g810 ( .A(n_376), .B(n_714), .Y(n_810) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g629 ( .A(n_377), .B(n_630), .Y(n_629) );
OR2x6_ASAP7_75t_L g735 ( .A(n_377), .B(n_595), .Y(n_735) );
AOI31xp33_ASAP7_75t_L g947 ( .A1(n_377), .A2(n_948), .A3(n_961), .B(n_972), .Y(n_947) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_377), .Y(n_1158) );
AND2x4_ASAP7_75t_L g1200 ( .A(n_377), .B(n_630), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_377), .B(n_702), .Y(n_1380) );
OR2x2_ASAP7_75t_L g1859 ( .A(n_377), .B(n_1860), .Y(n_1859) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x6_ASAP7_75t_L g518 ( .A(n_378), .B(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g684 ( .A(n_378), .Y(n_684) );
NAND5xp2_ASAP7_75t_SL g379 ( .A(n_380), .B(n_424), .C(n_435), .D(n_445), .E(n_460), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_391), .B1(n_392), .B2(n_404), .C(n_416), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_383), .A2(n_416), .B1(n_864), .B2(n_867), .C(n_869), .Y(n_863) );
INVx1_ASAP7_75t_L g963 ( .A(n_383), .Y(n_963) );
BUFx6f_ASAP7_75t_L g1049 ( .A(n_383), .Y(n_1049) );
INVx1_ASAP7_75t_L g1181 ( .A(n_383), .Y(n_1181) );
INVx2_ASAP7_75t_SL g1240 ( .A(n_383), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_383), .A2(n_1334), .B1(n_1440), .B2(n_1450), .C(n_1453), .Y(n_1449) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
BUFx3_ASAP7_75t_L g393 ( .A(n_384), .Y(n_393) );
BUFx6f_ASAP7_75t_L g792 ( .A(n_384), .Y(n_792) );
BUFx4f_ASAP7_75t_L g854 ( .A(n_384), .Y(n_854) );
INVx2_ASAP7_75t_SL g995 ( .A(n_384), .Y(n_995) );
AND2x4_ASAP7_75t_L g1334 ( .A(n_384), .B(n_581), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x4_ASAP7_75t_L g397 ( .A(n_386), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g409 ( .A(n_386), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_387), .Y(n_410) );
AND2x4_ASAP7_75t_L g414 ( .A(n_387), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g462 ( .A(n_388), .B(n_448), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_388), .A2(n_562), .B(n_567), .Y(n_561) );
AOI222xp33_ASAP7_75t_L g983 ( .A1(n_388), .A2(n_437), .B1(n_442), .B2(n_984), .C1(n_990), .C2(n_991), .Y(n_983) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_388), .A2(n_1153), .B(n_1156), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_388), .B(n_566), .Y(n_1306) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_388), .A2(n_426), .B1(n_1336), .B2(n_1337), .C(n_1342), .Y(n_1335) );
A2O1A1Ixp33_ASAP7_75t_L g1404 ( .A1(n_388), .A2(n_854), .B(n_1405), .C(n_1406), .Y(n_1404) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g427 ( .A(n_389), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g433 ( .A(n_389), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g763 ( .A(n_389), .B(n_483), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_SL g1902 ( .A1(n_389), .A2(n_1903), .B(n_1906), .C(n_1910), .Y(n_1902) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_391), .A2(n_425), .B1(n_546), .B2(n_549), .Y(n_545) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g802 ( .A(n_396), .Y(n_802) );
INVx1_ASAP7_75t_L g1141 ( .A(n_396), .Y(n_1141) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_397), .Y(n_448) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_397), .Y(n_566) );
INVx2_ASAP7_75t_SL g592 ( .A(n_397), .Y(n_592) );
BUFx3_ASAP7_75t_L g601 ( .A(n_397), .Y(n_601) );
AND2x6_ASAP7_75t_L g681 ( .A(n_397), .B(n_652), .Y(n_681) );
BUFx2_ASAP7_75t_L g954 ( .A(n_397), .Y(n_954) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_397), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g1138 ( .A(n_397), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g1330 ( .A(n_397), .Y(n_1330) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g1173 ( .A(n_400), .Y(n_1173) );
OAI221xp5_ASAP7_75t_L g1917 ( .A1(n_400), .A2(n_958), .B1(n_1889), .B2(n_1893), .C(n_1918), .Y(n_1917) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g595 ( .A(n_401), .Y(n_595) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_401), .Y(n_1059) );
INVx1_ASAP7_75t_L g1452 ( .A(n_401), .Y(n_1452) );
INVx1_ASAP7_75t_L g1860 ( .A(n_401), .Y(n_1860) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AND2x4_ASAP7_75t_L g459 ( .A(n_402), .B(n_421), .Y(n_459) );
INVx1_ASAP7_75t_L g683 ( .A(n_402), .Y(n_683) );
INVx2_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
INVx1_ASAP7_75t_L g653 ( .A(n_403), .Y(n_653) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_403), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_403), .Y(n_662) );
BUFx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_407), .Y(n_576) );
INVx1_ASAP7_75t_L g587 ( .A(n_407), .Y(n_587) );
INVx2_ASAP7_75t_L g679 ( .A(n_407), .Y(n_679) );
INVx1_ASAP7_75t_L g795 ( .A(n_407), .Y(n_795) );
INVx2_ASAP7_75t_SL g1312 ( .A(n_407), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1333 ( .A(n_407), .Y(n_1333) );
INVx6_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g472 ( .A(n_408), .B(n_419), .Y(n_472) );
BUFx2_ASAP7_75t_L g603 ( .A(n_408), .Y(n_603) );
AND2x4_ASAP7_75t_L g656 ( .A(n_408), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g772 ( .A(n_408), .Y(n_772) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g444 ( .A(n_409), .Y(n_444) );
INVx1_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g742 ( .A(n_413), .Y(n_742) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_413), .Y(n_858) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
INVx1_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_414), .Y(n_569) );
INVx1_ASAP7_75t_L g767 ( .A(n_414), .Y(n_767) );
INVx1_ASAP7_75t_L g429 ( .A(n_415), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_416), .A2(n_942), .B1(n_962), .B2(n_964), .C(n_968), .Y(n_961) );
AOI21xp33_ASAP7_75t_L g992 ( .A1(n_416), .A2(n_993), .B(n_997), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_416), .A2(n_1049), .B1(n_1050), .B2(n_1051), .C(n_1060), .Y(n_1048) );
INVx1_ASAP7_75t_L g1187 ( .A(n_416), .Y(n_1187) );
AOI221xp5_ASAP7_75t_L g1238 ( .A1(n_416), .A2(n_1239), .B1(n_1241), .B2(n_1242), .C(n_1244), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_416), .A2(n_1239), .B1(n_1300), .B2(n_1308), .C(n_1309), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_416), .A2(n_962), .B1(n_1532), .B2(n_1546), .C(n_1550), .Y(n_1545) );
INVx1_ASAP7_75t_L g1910 ( .A(n_416), .Y(n_1910) );
AND2x4_ASAP7_75t_L g416 ( .A(n_417), .B(n_422), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g1913 ( .A(n_418), .B(n_787), .Y(n_1913) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g437 ( .A(n_419), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g442 ( .A(n_419), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g581 ( .A(n_419), .Y(n_581) );
NAND2x1p5_ASAP7_75t_L g783 ( .A(n_419), .B(n_553), .Y(n_783) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_419), .B(n_438), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_419), .B(n_443), .Y(n_1186) );
AND2x4_ASAP7_75t_L g1318 ( .A(n_419), .B(n_443), .Y(n_1318) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g866 ( .A(n_422), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_422), .A2(n_566), .B1(n_988), .B2(n_989), .Y(n_987) );
BUFx6f_ASAP7_75t_L g1148 ( .A(n_422), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g650 ( .A(n_423), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g668 ( .A(n_423), .Y(n_668) );
INVx1_ASAP7_75t_L g1056 ( .A(n_423), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g1451 ( .A(n_423), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_431), .B2(n_432), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_426), .A2(n_432), .B1(n_871), .B2(n_872), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_426), .A2(n_432), .B1(n_938), .B2(n_940), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_426), .A2(n_432), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_426), .A2(n_462), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_426), .A2(n_462), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1303 ( .A1(n_426), .A2(n_1296), .B1(n_1299), .B2(n_1304), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_426), .A2(n_432), .B1(n_1434), .B2(n_1439), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_426), .A2(n_1306), .B1(n_1462), .B2(n_1463), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_426), .A2(n_432), .B1(n_1528), .B2(n_1531), .Y(n_1551) );
INVx6_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g564 ( .A(n_428), .Y(n_564) );
INVx1_ASAP7_75t_L g1144 ( .A(n_428), .Y(n_1144) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AND2x2_ASAP7_75t_L g572 ( .A(n_429), .B(n_430), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_431), .A2(n_461), .B1(n_533), .B2(n_540), .Y(n_544) );
AOI211xp5_ASAP7_75t_L g1230 ( .A1(n_432), .A2(n_1231), .B(n_1232), .C(n_1234), .Y(n_1230) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_432), .A2(n_1297), .B1(n_1314), .B2(n_1315), .C(n_1316), .Y(n_1313) );
AOI221xp5_ASAP7_75t_L g1464 ( .A1(n_432), .A2(n_1465), .B1(n_1466), .B2(n_1469), .C(n_1470), .Y(n_1464) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g589 ( .A(n_434), .Y(n_589) );
INVx1_ASAP7_75t_L g1155 ( .A(n_434), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B1(n_441), .B2(n_442), .Y(n_435) );
INVx2_ASAP7_75t_SL g861 ( .A(n_437), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_437), .A2(n_442), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
AOI222xp33_ASAP7_75t_L g1182 ( .A1(n_437), .A2(n_1003), .B1(n_1183), .B2(n_1184), .C1(n_1185), .C2(n_1186), .Y(n_1182) );
INVx1_ASAP7_75t_L g1538 ( .A(n_437), .Y(n_1538) );
INVx2_ASAP7_75t_SL g1912 ( .A(n_437), .Y(n_1912) );
INVxp67_ASAP7_75t_L g578 ( .A(n_438), .Y(n_578) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g781 ( .A(n_439), .Y(n_781) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g673 ( .A(n_440), .Y(n_673) );
INVx3_ASAP7_75t_L g862 ( .A(n_442), .Y(n_862) );
INVx1_ASAP7_75t_L g579 ( .A(n_443), .Y(n_579) );
INVx2_ASAP7_75t_L g787 ( .A(n_443), .Y(n_787) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x6_ASAP7_75t_L g675 ( .A(n_444), .B(n_653), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B1(n_450), .B2(n_453), .C(n_454), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g1920 ( .A1(n_446), .A2(n_568), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
INVxp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g966 ( .A(n_448), .Y(n_966) );
INVx1_ASAP7_75t_L g1541 ( .A(n_448), .Y(n_1541) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_449), .A2(n_492), .B1(n_493), .B2(n_497), .Y(n_491) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g1002 ( .A(n_452), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_453), .A2(n_476), .B1(n_486), .B2(n_487), .Y(n_475) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g996 ( .A(n_457), .Y(n_996) );
INVx1_ASAP7_75t_L g1544 ( .A(n_458), .Y(n_1544) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g604 ( .A(n_459), .Y(n_604) );
AND2x4_ASAP7_75t_L g744 ( .A(n_459), .B(n_471), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_459), .Y(n_856) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_459), .Y(n_1145) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_459), .Y(n_1401) );
AND2x4_ASAP7_75t_L g1864 ( .A(n_459), .B(n_471), .Y(n_1864) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_462), .A2(n_853), .B1(n_857), .B2(n_859), .C(n_860), .Y(n_852) );
INVx1_ASAP7_75t_L g950 ( .A(n_462), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_462), .A2(n_1039), .B(n_1040), .Y(n_1038) );
AOI211xp5_ASAP7_75t_L g1536 ( .A1(n_462), .A2(n_1529), .B(n_1537), .C(n_1539), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_464), .A2(n_850), .B1(n_851), .B2(n_873), .Y(n_849) );
AOI21xp33_ASAP7_75t_SL g1035 ( .A1(n_464), .A2(n_1036), .B(n_1037), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_464), .A2(n_1066), .B1(n_1229), .B2(n_1249), .Y(n_1228) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g945 ( .A(n_465), .Y(n_945) );
INVx1_ASAP7_75t_L g1320 ( .A(n_465), .Y(n_1320) );
INVx2_ASAP7_75t_SL g1455 ( .A(n_465), .Y(n_1455) );
INVx2_ASAP7_75t_L g1478 ( .A(n_465), .Y(n_1478) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
INVx2_ASAP7_75t_L g609 ( .A(n_466), .Y(n_609) );
INVx3_ASAP7_75t_L g510 ( .A(n_467), .Y(n_510) );
INVx1_ASAP7_75t_L g692 ( .A(n_468), .Y(n_692) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x6_ASAP7_75t_L g809 ( .A(n_470), .B(n_810), .Y(n_809) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g1004 ( .A(n_472), .Y(n_1004) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_503), .C(n_517), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_491), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_476), .A2(n_487), .B1(n_914), .B2(n_915), .Y(n_913) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g878 ( .A(n_477), .Y(n_878) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_477), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1105 ( .A(n_477), .Y(n_1105) );
BUFx2_ASAP7_75t_L g1353 ( .A(n_477), .Y(n_1353) );
BUFx2_ASAP7_75t_L g1483 ( .A(n_477), .Y(n_1483) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
BUFx3_ASAP7_75t_L g901 ( .A(n_478), .Y(n_901) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_479), .Y(n_542) );
INVx3_ASAP7_75t_L g620 ( .A(n_479), .Y(n_620) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_480), .Y(n_632) );
INVx1_ASAP7_75t_L g729 ( .A(n_480), .Y(n_729) );
INVx1_ASAP7_75t_L g1845 ( .A(n_480), .Y(n_1845) );
AND2x4_ASAP7_75t_L g489 ( .A(n_481), .B(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_L g487 ( .A(n_482), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g493 ( .A(n_482), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g497 ( .A(n_482), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g607 ( .A(n_482), .B(n_498), .Y(n_607) );
AND2x2_ASAP7_75t_L g616 ( .A(n_482), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g619 ( .A(n_482), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g635 ( .A(n_482), .B(n_628), .Y(n_635) );
AND2x2_ASAP7_75t_L g919 ( .A(n_482), .B(n_498), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_482), .A2(n_551), .B1(n_1008), .B2(n_1016), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_482), .B(n_498), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_482), .B(n_498), .Y(n_1488) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g553 ( .A(n_483), .Y(n_553) );
INVx2_ASAP7_75t_L g719 ( .A(n_484), .Y(n_719) );
AND2x4_ASAP7_75t_L g722 ( .A(n_484), .B(n_627), .Y(n_722) );
AND2x2_ASAP7_75t_L g725 ( .A(n_484), .B(n_499), .Y(n_725) );
INVx1_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
INVx1_ASAP7_75t_L g555 ( .A(n_485), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_487), .A2(n_877), .B1(n_878), .B2(n_879), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_487), .A2(n_1044), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_487), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
INVx1_ASAP7_75t_SL g1191 ( .A(n_487), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_487), .A2(n_878), .B1(n_1236), .B2(n_1264), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_487), .A2(n_878), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
AOI22xp5_ASAP7_75t_L g1348 ( .A1(n_487), .A2(n_1268), .B1(n_1349), .B2(n_1350), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_487), .A2(n_607), .B1(n_1385), .B2(n_1386), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_487), .A2(n_1482), .B1(n_1483), .B2(n_1484), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_487), .A2(n_1353), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_488), .B(n_510), .Y(n_516) );
BUFx2_ASAP7_75t_L g1199 ( .A(n_488), .Y(n_1199) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_489), .Y(n_628) );
BUFx2_ASAP7_75t_L g641 ( .A(n_489), .Y(n_641) );
INVx1_ASAP7_75t_L g711 ( .A(n_489), .Y(n_711) );
BUFx3_ASAP7_75t_L g720 ( .A(n_489), .Y(n_720) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_489), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1827 ( .A(n_489), .B(n_1828), .Y(n_1827) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_493), .A2(n_497), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_493), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_493), .A2(n_497), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_493), .A2(n_1111), .B(n_1112), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_493), .A2(n_497), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_493), .A2(n_1266), .B1(n_1267), .B2(n_1268), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_493), .A2(n_1268), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_493), .B(n_1382), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_493), .A2(n_1486), .B1(n_1487), .B2(n_1488), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_493), .A2(n_919), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g617 ( .A(n_495), .Y(n_617) );
INVx2_ASAP7_75t_L g1198 ( .A(n_495), .Y(n_1198) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_496), .Y(n_627) );
INVx2_ASAP7_75t_SL g1213 ( .A(n_498), .Y(n_1213) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_499), .Y(n_624) );
INVx1_ASAP7_75t_L g1018 ( .A(n_499), .Y(n_1018) );
INVx1_ASAP7_75t_L g1027 ( .A(n_499), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_499), .Y(n_1194) );
BUFx6f_ASAP7_75t_L g1378 ( .A(n_499), .Y(n_1378) );
AND2x4_ASAP7_75t_L g1837 ( .A(n_499), .B(n_1838), .Y(n_1837) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g514 ( .A(n_500), .Y(n_514) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g921 ( .A(n_505), .Y(n_921) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g1490 ( .A(n_506), .Y(n_1490) );
NAND2x1_ASAP7_75t_SL g506 ( .A(n_507), .B(n_510), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g704 ( .A(n_507), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_507), .A2(n_513), .B1(n_1184), .B2(n_1185), .Y(n_1205) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_509), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_510), .B(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g611 ( .A(n_510), .B(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g637 ( .A(n_510), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g640 ( .A(n_510), .B(n_641), .Y(n_640) );
AOI32xp33_ASAP7_75t_L g1192 ( .A1(n_510), .A2(n_1193), .A3(n_1197), .B1(n_1200), .B2(n_1201), .Y(n_1192) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx4f_ASAP7_75t_L g922 ( .A(n_512), .Y(n_922) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x6_ASAP7_75t_L g706 ( .A(n_514), .B(n_691), .Y(n_706) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g884 ( .A(n_516), .Y(n_884) );
BUFx2_ASAP7_75t_L g1282 ( .A(n_516), .Y(n_1282) );
OAI33xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .A3(n_532), .B1(n_544), .B2(n_545), .B3(n_550), .Y(n_517) );
OAI33xp33_ASAP7_75t_L g885 ( .A1(n_518), .A2(n_886), .A3(n_892), .B1(n_899), .B2(n_902), .B3(n_905), .Y(n_885) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_518), .Y(n_924) );
OAI33xp33_ASAP7_75t_L g1076 ( .A1(n_518), .A2(n_905), .A3(n_1077), .B1(n_1081), .B2(n_1087), .B3(n_1090), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_518), .A2(n_905), .B1(n_1113), .B2(n_1123), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_518), .Y(n_1284) );
OAI33xp33_ASAP7_75t_L g1421 ( .A1(n_518), .A2(n_943), .A3(n_1422), .B1(n_1425), .B2(n_1431), .B3(n_1438), .Y(n_1421) );
OAI33xp33_ASAP7_75t_L g1491 ( .A1(n_518), .A2(n_905), .A3(n_1492), .B1(n_1496), .B2(n_1501), .B3(n_1502), .Y(n_1491) );
OAI33xp33_ASAP7_75t_L g1516 ( .A1(n_518), .A2(n_905), .A3(n_1517), .B1(n_1522), .B2(n_1527), .B3(n_1530), .Y(n_1516) );
INVx1_ASAP7_75t_L g1838 ( .A(n_520), .Y(n_1838) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B1(n_525), .B2(n_531), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g1891 ( .A1(n_522), .A2(n_828), .B1(n_1892), .B2(n_1893), .Y(n_1891) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g1078 ( .A(n_523), .Y(n_1078) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g928 ( .A(n_526), .Y(n_928) );
INVx2_ASAP7_75t_L g1216 ( .A(n_526), .Y(n_1216) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
BUFx3_ASAP7_75t_L g828 ( .A(n_527), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_527), .A2(n_1204), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_L g690 ( .A(n_529), .B(n_530), .Y(n_690) );
INVx1_ASAP7_75t_L g613 ( .A(n_530), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_539), .B1(n_540), .B2(n_543), .Y(n_532) );
OAI22xp33_ASAP7_75t_SL g929 ( .A1(n_533), .A2(n_930), .B1(n_932), .B2(n_933), .Y(n_929) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_535), .A2(n_1039), .B1(n_1064), .B2(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1888 ( .A1(n_535), .A2(n_1196), .B1(n_1889), .B2(n_1890), .Y(n_1888) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g815 ( .A(n_536), .Y(n_815) );
INVx2_ASAP7_75t_SL g936 ( .A(n_536), .Y(n_936) );
INVx2_ASAP7_75t_L g1433 ( .A(n_536), .Y(n_1433) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g896 ( .A(n_537), .Y(n_896) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g836 ( .A(n_538), .Y(n_836) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_538), .Y(n_1116) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g694 ( .A(n_542), .Y(n_694) );
INVx2_ASAP7_75t_L g1119 ( .A(n_542), .Y(n_1119) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g826 ( .A1(n_547), .A2(n_827), .B1(n_829), .B2(n_830), .C(n_831), .Y(n_826) );
OAI22xp5_ASAP7_75t_SL g1438 ( .A1(n_547), .A2(n_928), .B1(n_1439), .B2(n_1440), .Y(n_1438) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_551), .A2(n_597), .A3(n_623), .B1(n_625), .B2(n_629), .C1(n_631), .C2(n_635), .Y(n_622) );
INVx1_ASAP7_75t_L g943 ( .A(n_551), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_551), .A2(n_878), .B1(n_1211), .B2(n_1217), .Y(n_1210) );
AOI33xp33_ASAP7_75t_L g1254 ( .A1(n_551), .A2(n_629), .A3(n_1255), .B1(n_1257), .B2(n_1258), .B3(n_1261), .Y(n_1254) );
AOI222xp33_ASAP7_75t_L g1355 ( .A1(n_551), .A2(n_616), .B1(n_629), .B2(n_1356), .C1(n_1357), .C2(n_1362), .Y(n_1355) );
INVx6_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx5_ASAP7_75t_L g906 ( .A(n_552), .Y(n_906) );
OR2x6_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g702 ( .A(n_554), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g1829 ( .A(n_555), .Y(n_1829) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_573), .C(n_582), .D(n_596), .Y(n_560) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g737 ( .A(n_564), .Y(n_737) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_564), .Y(n_747) );
INVx2_ASAP7_75t_L g985 ( .A(n_564), .Y(n_985) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g1053 ( .A(n_566), .Y(n_1053) );
INVx1_ASAP7_75t_L g1245 ( .A(n_568), .Y(n_1245) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x6_ASAP7_75t_L g660 ( .A(n_569), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g797 ( .A(n_569), .Y(n_797) );
INVx1_ASAP7_75t_L g971 ( .A(n_569), .Y(n_971) );
BUFx6f_ASAP7_75t_L g1061 ( .A(n_569), .Y(n_1061) );
BUFx6f_ASAP7_75t_L g1130 ( .A(n_569), .Y(n_1130) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g1045 ( .A(n_571), .Y(n_1045) );
INVx1_ASAP7_75t_L g1395 ( .A(n_571), .Y(n_1395) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g585 ( .A(n_572), .Y(n_585) );
INVx1_ASAP7_75t_L g959 ( .A(n_572), .Y(n_959) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_572), .Y(n_1135) );
INVx1_ASAP7_75t_L g1339 ( .A(n_572), .Y(n_1339) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_577), .C(n_580), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_574), .A2(n_609), .B1(n_610), .B2(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g800 ( .A(n_576), .Y(n_800) );
INVx4_ASAP7_75t_L g855 ( .A(n_576), .Y(n_855) );
A2O1A1Ixp33_ASAP7_75t_L g1147 ( .A1(n_580), .A2(n_603), .B(n_1109), .C(n_1148), .Y(n_1147) );
BUFx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_586), .C(n_590), .Y(n_582) );
OAI211xp5_ASAP7_75t_L g1398 ( .A1(n_584), .A2(n_1386), .B(n_1399), .C(n_1400), .Y(n_1398) );
BUFx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g599 ( .A(n_585), .Y(n_599) );
OR2x6_ASAP7_75t_L g775 ( .A(n_585), .B(n_763), .Y(n_775) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_587), .Y(n_969) );
INVx1_ASAP7_75t_L g1132 ( .A(n_587), .Y(n_1132) );
INVx1_ASAP7_75t_L g986 ( .A(n_588), .Y(n_986) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g750 ( .A(n_589), .Y(n_750) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g761 ( .A(n_592), .Y(n_761) );
INVx1_ASAP7_75t_L g1473 ( .A(n_592), .Y(n_1473) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .C(n_602), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_598), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_598), .A2(n_716), .B1(n_721), .B2(n_746), .C(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g741 ( .A(n_601), .Y(n_741) );
INVx2_ASAP7_75t_SL g1908 ( .A(n_601), .Y(n_1908) );
INVx1_ASAP7_75t_L g1926 ( .A(n_604), .Y(n_1926) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g1417 ( .A1(n_607), .A2(n_616), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
INVx1_ASAP7_75t_L g1882 ( .A(n_607), .Y(n_1882) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_609), .A2(n_629), .B1(n_1005), .B2(n_1025), .Y(n_1024) );
AOI22xp33_ASAP7_75t_SL g1107 ( .A1(n_609), .A2(n_919), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_609), .A2(n_1352), .B1(n_1353), .B2(n_1354), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_609), .A2(n_619), .B1(n_1388), .B2(n_1389), .Y(n_1387) );
AOI221xp5_ASAP7_75t_L g1032 ( .A1(n_611), .A2(n_637), .B1(n_640), .B2(n_990), .C(n_991), .Y(n_1032) );
INVx1_ASAP7_75t_L g1161 ( .A(n_611), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_611), .A2(n_637), .B1(n_640), .B2(n_1252), .C(n_1253), .Y(n_1251) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_611), .A2(n_637), .B1(n_640), .B2(n_1346), .C(n_1347), .Y(n_1345) );
AOI221xp5_ASAP7_75t_L g1371 ( .A1(n_611), .A2(n_637), .B1(n_640), .B2(n_1372), .C(n_1373), .Y(n_1371) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_618), .B2(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g1900 ( .A(n_616), .Y(n_1900) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_617), .B(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g1414 ( .A1(n_619), .A2(n_635), .B1(n_1415), .B2(n_1416), .Y(n_1414) );
INVx2_ASAP7_75t_L g1884 ( .A(n_619), .Y(n_1884) );
INVx1_ASAP7_75t_L g1020 ( .A(n_620), .Y(n_1020) );
INVx2_ASAP7_75t_L g1089 ( .A(n_620), .Y(n_1089) );
INVx2_ASAP7_75t_L g1260 ( .A(n_620), .Y(n_1260) );
INVx2_ASAP7_75t_L g1365 ( .A(n_620), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_636), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g1010 ( .A1(n_626), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g700 ( .A(n_627), .Y(n_700) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_628), .Y(n_818) );
AOI33xp33_ASAP7_75t_L g1374 ( .A1(n_629), .A2(n_1375), .A3(n_1376), .B1(n_1377), .B2(n_1379), .B3(n_1380), .Y(n_1374) );
INVx1_ASAP7_75t_L g832 ( .A(n_630), .Y(n_832) );
INVx2_ASAP7_75t_SL g816 ( .A(n_632), .Y(n_816) );
INVx2_ASAP7_75t_SL g898 ( .A(n_632), .Y(n_898) );
INVx2_ASAP7_75t_SL g1009 ( .A(n_632), .Y(n_1009) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_632), .Y(n_1085) );
INVx4_ASAP7_75t_L g1196 ( .A(n_632), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_640), .Y(n_636) );
INVx1_ASAP7_75t_L g1163 ( .A(n_637), .Y(n_1163) );
AND2x2_ASAP7_75t_L g822 ( .A(n_638), .B(n_715), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g1159 ( .A1(n_640), .A2(n_1150), .B1(n_1151), .B2(n_1160), .C(n_1162), .Y(n_1159) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI221x1_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_682), .B1(n_685), .B2(n_730), .C(n_732), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .C(n_663), .D(n_676), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g1807 ( .A(n_649), .B(n_1808), .C(n_1812), .D(n_1815), .Y(n_1807) );
INVx5_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_652), .B(n_1451), .Y(n_1816) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_659), .B2(n_660), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_655), .A2(n_713), .B1(n_716), .B2(n_717), .C1(n_721), .C2(n_722), .Y(n_712) );
AOI22xp5_ASAP7_75t_SL g1808 ( .A1(n_656), .A2(n_1809), .B1(n_1810), .B2(n_1811), .Y(n_1808) );
AND2x4_ASAP7_75t_L g671 ( .A(n_657), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g1812 ( .A1(n_660), .A2(n_681), .B1(n_1813), .B2(n_1814), .Y(n_1812) );
AND2x4_ASAP7_75t_L g678 ( .A(n_661), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g1810 ( .A(n_661), .B(n_679), .Y(n_1810) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_662), .B(n_1821), .Y(n_1820) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_669), .B2(n_670), .C1(n_674), .C2(n_675), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_664), .A2(n_696), .B(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g1549 ( .A(n_668), .Y(n_1549) );
BUFx4f_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g1821 ( .A(n_673), .Y(n_1821) );
INVx3_ASAP7_75t_L g1822 ( .A(n_675), .Y(n_1822) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_681), .Y(n_676) );
AND2x4_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x4_ASAP7_75t_L g1823 ( .A(n_683), .B(n_684), .Y(n_1823) );
INVx2_ASAP7_75t_L g731 ( .A(n_684), .Y(n_731) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_684), .Y(n_1066) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_712), .C(n_723), .Y(n_685) );
NOR3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_693), .C(n_703), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x6_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g697 ( .A(n_689), .Y(n_697) );
OR2x2_ASAP7_75t_L g842 ( .A(n_689), .B(n_691), .Y(n_842) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_689), .Y(n_941) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g891 ( .A(n_690), .Y(n_891) );
BUFx2_ASAP7_75t_L g904 ( .A(n_690), .Y(n_904) );
INVx3_ASAP7_75t_L g1023 ( .A(n_690), .Y(n_1023) );
INVx1_ASAP7_75t_L g705 ( .A(n_691), .Y(n_705) );
INVx1_ASAP7_75t_L g715 ( .A(n_691), .Y(n_715) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g819 ( .A(n_700), .Y(n_819) );
INVx2_ASAP7_75t_L g1122 ( .A(n_700), .Y(n_1122) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
CKINVDCx11_ASAP7_75t_R g823 ( .A(n_706), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx8_ASAP7_75t_L g813 ( .A(n_717), .Y(n_813) );
AND2x4_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
AND2x4_ASAP7_75t_L g727 ( .A(n_718), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx6f_ASAP7_75t_L g1127 ( .A(n_720), .Y(n_1127) );
CKINVDCx6p67_ASAP7_75t_R g825 ( .A(n_722), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_723) );
INVx3_ASAP7_75t_L g844 ( .A(n_725), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_727), .Y(n_845) );
INVx1_ASAP7_75t_L g840 ( .A(n_728), .Y(n_840) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g1437 ( .A(n_729), .Y(n_1437) );
OAI31xp33_ASAP7_75t_L g811 ( .A1(n_730), .A2(n_812), .A3(n_824), .B(n_843), .Y(n_811) );
INVx5_ASAP7_75t_L g1188 ( .A(n_730), .Y(n_1188) );
BUFx8_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g850 ( .A(n_731), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B1(n_743), .B2(n_745), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_735), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g1923 ( .A1(n_737), .A2(n_958), .B1(n_1924), .B2(n_1925), .C(n_1926), .Y(n_1923) );
INVx4_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI33xp33_ASAP7_75t_L g788 ( .A1(n_744), .A2(n_789), .A3(n_790), .B1(n_793), .B2(n_798), .B3(n_801), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g1915 ( .A1(n_746), .A2(n_1890), .B1(n_1892), .B2(n_1916), .Y(n_1915) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_1221), .B1(n_1222), .B2(n_1556), .Y(n_751) );
INVx1_ASAP7_75t_L g1556 ( .A(n_752), .Y(n_1556) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_975), .Y(n_752) );
XNOR2x1_ASAP7_75t_L g753 ( .A(n_754), .B(n_846), .Y(n_753) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_807), .C(n_811), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_776), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_768), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_764), .B2(n_765), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g814 ( .A1(n_759), .A2(n_764), .B1(n_815), .B2(n_816), .C(n_817), .Y(n_814) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AND2x2_ASAP7_75t_L g770 ( .A(n_762), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OR2x6_ASAP7_75t_L g766 ( .A(n_763), .B(n_767), .Y(n_766) );
CKINVDCx6p67_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g1905 ( .A(n_767), .Y(n_1905) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_773), .B2(n_774), .Y(n_768) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g868 ( .A(n_772), .Y(n_868) );
INVx1_ASAP7_75t_L g1467 ( .A(n_772), .Y(n_1467) );
CKINVDCx6p67_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
NAND3xp33_ASAP7_75t_SL g776 ( .A(n_777), .B(n_788), .C(n_803), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_784), .B2(n_785), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_778), .A2(n_784), .B1(n_821), .B2(n_823), .Y(n_820) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
OR2x6_ASAP7_75t_L g786 ( .A(n_783), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g806 ( .A(n_783), .Y(n_806) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_792), .B(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_SL g1909 ( .A(n_792), .Y(n_1909) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_816), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
INVxp67_ASAP7_75t_L g1028 ( .A(n_816), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
BUFx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_837), .B1(n_838), .B2(n_841), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g1082 ( .A(n_836), .Y(n_1082) );
INVx1_ASAP7_75t_L g1428 ( .A(n_836), .Y(n_1428) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AO22x2_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_908), .B1(n_973), .B2(n_974), .Y(n_846) );
INVx1_ASAP7_75t_L g974 ( .A(n_847), .Y(n_974) );
XOR2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_907), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_874), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_850), .A2(n_1460), .B1(n_1477), .B2(n_1478), .Y(n_1459) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_863), .C(n_870), .Y(n_851) );
BUFx2_ASAP7_75t_L g967 ( .A(n_854), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1903 ( .A1(n_855), .A2(n_1896), .B1(n_1898), .B2(n_1904), .Y(n_1903) );
INVx1_ASAP7_75t_L g1916 ( .A(n_858), .Y(n_1916) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_859), .A2(n_872), .B1(n_894), .B2(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g1243 ( .A(n_866), .Y(n_1243) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_869), .A2(n_871), .B1(n_888), .B2(n_903), .Y(n_902) );
NOR3xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_883), .C(n_885), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_880), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_890), .B2(n_891), .Y(n_886) );
BUFx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_889), .A2(n_940), .B1(n_941), .B2(n_942), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g1021 ( .A1(n_889), .A2(n_989), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_889), .A2(n_1023), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
INVx1_ASAP7_75t_L g1092 ( .A(n_889), .Y(n_1092) );
INVx1_ASAP7_75t_L g1287 ( .A(n_889), .Y(n_1287) );
OAI22xp33_ASAP7_75t_L g1527 ( .A1(n_889), .A2(n_1295), .B1(n_1528), .B2(n_1529), .Y(n_1527) );
OAI22xp5_ASAP7_75t_SL g1897 ( .A1(n_889), .A2(n_928), .B1(n_1898), .B2(n_1899), .Y(n_1897) );
OAI22xp33_ASAP7_75t_L g1422 ( .A1(n_891), .A2(n_1202), .B1(n_1423), .B2(n_1424), .Y(n_1422) );
OAI22xp5_ASAP7_75t_SL g892 ( .A1(n_893), .A2(n_894), .B1(n_897), .B2(n_898), .Y(n_892) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g1498 ( .A(n_895), .Y(n_1498) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_896), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_898), .A2(n_935), .B1(n_937), .B2(n_938), .Y(n_934) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_898), .A2(n_936), .B1(n_1124), .B2(n_1125), .C(n_1126), .Y(n_1123) );
OAI22xp33_ASAP7_75t_L g1530 ( .A1(n_900), .A2(n_1519), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_901), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1077 ( .A1(n_903), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
OAI22xp33_ASAP7_75t_L g1492 ( .A1(n_903), .A2(n_1493), .B1(n_1494), .B2(n_1495), .Y(n_1492) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI33xp33_ASAP7_75t_L g1283 ( .A1(n_905), .A2(n_1284), .A3(n_1285), .B1(n_1290), .B2(n_1294), .B3(n_1298), .Y(n_1283) );
CKINVDCx8_ASAP7_75t_R g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g973 ( .A(n_908), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_944), .Y(n_910) );
NOR3xp33_ASAP7_75t_SL g911 ( .A(n_912), .B(n_920), .C(n_923), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_916), .Y(n_912) );
OAI33xp33_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_925), .A3(n_929), .B1(n_934), .B2(n_939), .B3(n_943), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g1298 ( .A1(n_928), .A2(n_1286), .B1(n_1299), .B2(n_1300), .Y(n_1298) );
OAI22xp33_ASAP7_75t_L g1502 ( .A1(n_928), .A2(n_1462), .B1(n_1476), .B2(n_1493), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1517 ( .A1(n_930), .A2(n_1518), .B1(n_1519), .B2(n_1521), .Y(n_1517) );
INVx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_937), .A2(n_949), .B(n_951), .Y(n_948) );
AOI21xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B(n_947), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g1533 ( .A1(n_945), .A2(n_1534), .B(n_1535), .Y(n_1533) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
AOI31xp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .A3(n_956), .B(n_960), .Y(n_952) );
INVx1_ASAP7_75t_L g1340 ( .A(n_954), .Y(n_1340) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
BUFx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_1096), .B1(n_1097), .B2(n_1220), .Y(n_975) );
INVx1_ASAP7_75t_L g1220 ( .A(n_976), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_1033), .B2(n_1095), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
XNOR2x1_ASAP7_75t_L g979 ( .A(n_980), .B(n_981), .Y(n_979) );
OR2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_1006), .Y(n_981) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g1176 ( .A(n_995), .Y(n_1176) );
INVx1_ASAP7_75t_L g1468 ( .A(n_995), .Y(n_1468) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1001), .B1(n_1003), .B2(n_1005), .Y(n_998) );
INVx2_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND3xp33_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1024), .C(n_1032), .Y(n_1006) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1014), .Y(n_1256) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1020), .Y(n_1525) );
BUFx2_ASAP7_75t_L g1093 ( .A(n_1023), .Y(n_1093) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1023), .Y(n_1520) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1027), .Y(n_1363) );
INVx1_ASAP7_75t_SL g1095 ( .A(n_1033), .Y(n_1095) );
XNOR2x1_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1094), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1067), .Y(n_1034) );
AOI31xp33_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1048), .A3(n_1062), .B(n_1065), .Y(n_1037) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_SL g1343 ( .A(n_1042), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_1042), .A2(n_1318), .B1(n_1372), .B2(n_1373), .Y(n_1407) );
INVx4_ASAP7_75t_L g1447 ( .A(n_1042), .Y(n_1447) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B(n_1046), .C(n_1047), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1142 ( .A1(n_1045), .A2(n_1106), .B1(n_1111), .B2(n_1143), .C(n_1145), .Y(n_1142) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_1050), .A2(n_1063), .B1(n_1091), .B2(n_1093), .Y(n_1090) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1058), .A2(n_1117), .B1(n_1134), .B2(n_1136), .C(n_1137), .Y(n_1133) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1341 ( .A(n_1061), .Y(n_1341) );
AOI21xp5_ASAP7_75t_L g1325 ( .A1(n_1065), .A2(n_1326), .B(n_1335), .Y(n_1325) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI31xp33_ASAP7_75t_L g1390 ( .A1(n_1066), .A2(n_1391), .A3(n_1392), .B(n_1403), .Y(n_1390) );
NOR3xp33_ASAP7_75t_SL g1067 ( .A(n_1068), .B(n_1075), .C(n_1076), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1072), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1214 ( .A1(n_1078), .A2(n_1178), .B1(n_1215), .B2(n_1216), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1084), .B2(n_1086), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_1082), .Y(n_1291) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1089), .Y(n_1358) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OAI22xp33_ASAP7_75t_L g1285 ( .A1(n_1093), .A2(n_1286), .B1(n_1288), .B2(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B1(n_1164), .B2(n_1165), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
NAND4xp25_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1110), .C(n_1128), .D(n_1159), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1107), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1117), .B1(n_1118), .B2(n_1120), .C(n_1121), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1522 ( .A1(n_1114), .A2(n_1523), .B1(n_1524), .B2(n_1526), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1894 ( .A1(n_1114), .A2(n_1365), .B1(n_1895), .B2(n_1896), .Y(n_1894) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
OAI31xp33_ASAP7_75t_SL g1128 ( .A1(n_1129), .A2(n_1139), .A3(n_1146), .B(n_1157), .Y(n_1128) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
OAI21xp5_ASAP7_75t_SL g1235 ( .A1(n_1134), .A2(n_1236), .B(n_1237), .Y(n_1235) );
INVx2_ASAP7_75t_SL g1134 ( .A(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1135), .Y(n_1543) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1137), .Y(n_1172) );
INVx2_ASAP7_75t_SL g1137 ( .A(n_1138), .Y(n_1137) );
BUFx3_ASAP7_75t_L g1919 ( .A(n_1138), .Y(n_1919) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g1542 ( .A1(n_1143), .A2(n_1511), .B1(n_1513), .B2(n_1543), .C(n_1544), .Y(n_1542) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1149), .C(n_1152), .Y(n_1146) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_1157), .A2(n_1442), .B1(n_1455), .B2(n_1456), .Y(n_1441) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1157), .Y(n_1552) );
OAI31xp33_ASAP7_75t_L g1901 ( .A1(n_1157), .A2(n_1902), .A3(n_1911), .B(n_1914), .Y(n_1901) );
CKINVDCx8_ASAP7_75t_R g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1219 ( .A(n_1166), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1189), .Y(n_1166) );
OAI21xp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1180), .B(n_1188), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B1(n_1174), .B2(n_1175), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1233 ( .A(n_1186), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1301 ( .A1(n_1188), .A2(n_1302), .B1(n_1319), .B2(n_1320), .Y(n_1301) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1206), .Y(n_1189) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_1196), .A2(n_1291), .B1(n_1292), .B2(n_1293), .Y(n_1290) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_1196), .A2(n_1295), .B1(n_1296), .B2(n_1297), .Y(n_1294) );
BUFx3_ASAP7_75t_L g1262 ( .A(n_1198), .Y(n_1262) );
NAND3xp33_ASAP7_75t_L g1849 ( .A(n_1200), .B(n_1850), .C(n_1851), .Y(n_1849) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx2_ASAP7_75t_SL g1493 ( .A(n_1203), .Y(n_1493) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1204), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1210), .Y(n_1206) );
INVx3_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
OAI21x1_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1503), .B(n_1555), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1555 ( .A(n_1224), .B(n_1504), .Y(n_1555) );
XNOR2xp5_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1321), .Y(n_1224) );
XOR2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1270), .Y(n_1225) );
XNOR2xp5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1269), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1250), .Y(n_1227) );
NAND3xp33_ASAP7_75t_SL g1229 ( .A(n_1230), .B(n_1238), .C(n_1246), .Y(n_1229) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1240), .Y(n_1475) );
AND4x1_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1254), .C(n_1263), .D(n_1265), .Y(n_1250) );
AOI211xp5_ASAP7_75t_L g1825 ( .A1(n_1256), .A2(n_1826), .B(n_1827), .C(n_1830), .Y(n_1825) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_1260), .A2(n_1463), .B1(n_1465), .B2(n_1498), .Y(n_1501) );
XNOR2x1_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1272), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1301), .Y(n_1272) );
NOR3xp33_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1281), .C(n_1283), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1307), .C(n_1313), .Y(n_1302) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_1306), .A2(n_1432), .B1(n_1444), .B2(n_1445), .C(n_1446), .Y(n_1443) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx2_ASAP7_75t_SL g1448 ( .A(n_1318), .Y(n_1448) );
XOR2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1408), .Y(n_1321) );
XNOR2x1_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1368), .Y(n_1322) );
NOR2x1_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1344), .Y(n_1324) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B1(n_1329), .B2(n_1331), .C(n_1334), .Y(n_1326) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1334), .Y(n_1402) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_1334), .A2(n_1472), .B1(n_1474), .B2(n_1475), .C(n_1476), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NAND4xp25_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1348), .C(n_1351), .D(n_1355), .Y(n_1344) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1358), .Y(n_1500) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1364), .Y(n_1430) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NAND3xp33_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1383), .C(n_1390), .Y(n_1369) );
AND3x1_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1374), .C(n_1381), .Y(n_1370) );
NAND3xp33_ASAP7_75t_L g1852 ( .A(n_1380), .B(n_1853), .C(n_1854), .Y(n_1852) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1387), .Y(n_1383) );
NAND3xp33_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1398), .C(n_1402), .Y(n_1392) );
OAI211xp5_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1395), .B(n_1396), .C(n_1397), .Y(n_1393) );
XNOR2xp5_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1457), .Y(n_1408) );
XNOR2x1_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1411), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1441), .Y(n_1411) );
NOR3xp33_ASAP7_75t_L g1412 ( .A(n_1413), .B(n_1420), .C(n_1421), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1417), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_1426), .A2(n_1427), .B1(n_1429), .B2(n_1430), .Y(n_1425) );
BUFx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OAI22xp5_ASAP7_75t_SL g1431 ( .A1(n_1432), .A2(n_1433), .B1(n_1434), .B2(n_1435), .Y(n_1431) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
NAND3xp33_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1449), .C(n_1454), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1479), .Y(n_1458) );
NAND3xp33_ASAP7_75t_SL g1460 ( .A(n_1461), .B(n_1464), .C(n_1471), .Y(n_1460) );
NOR3xp33_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1489), .C(n_1491), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1485), .Y(n_1480) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_1497), .A2(n_1498), .B1(n_1499), .B2(n_1500), .Y(n_1496) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
HB1xp67_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1506), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1507), .B(n_1533), .Y(n_1506) );
NOR3xp33_ASAP7_75t_L g1507 ( .A(n_1508), .B(n_1515), .C(n_1516), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1512), .Y(n_1508) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx2_ASAP7_75t_SL g1524 ( .A(n_1525), .Y(n_1524) );
AOI31xp33_ASAP7_75t_L g1535 ( .A1(n_1536), .A2(n_1545), .A3(n_1551), .B(n_1552), .Y(n_1535) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
OAI221xp5_ASAP7_75t_SL g1557 ( .A1(n_1558), .A2(n_1800), .B1(n_1802), .B2(n_1865), .C(n_1871), .Y(n_1557) );
AND5x1_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1719), .C(n_1766), .D(n_1779), .E(n_1793), .Y(n_1558) );
OAI31xp33_ASAP7_75t_SL g1559 ( .A1(n_1560), .A2(n_1645), .A3(n_1680), .B(n_1709), .Y(n_1559) );
OAI322xp33_ASAP7_75t_L g1560 ( .A1(n_1561), .A2(n_1591), .A3(n_1609), .B1(n_1613), .B2(n_1619), .C1(n_1632), .C2(n_1634), .Y(n_1560) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
A2O1A1Ixp33_ASAP7_75t_L g1740 ( .A1(n_1562), .A2(n_1621), .B(n_1677), .C(n_1741), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1583), .Y(n_1562) );
NOR2xp33_ASAP7_75t_L g1672 ( .A(n_1563), .B(n_1657), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1563), .B(n_1609), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1563), .B(n_1652), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1563), .B(n_1630), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1563), .B(n_1584), .Y(n_1792) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1563), .Y(n_1798) );
INVx4_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx3_ASAP7_75t_L g1615 ( .A(n_1564), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1564), .B(n_1654), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1564), .B(n_1652), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1564), .B(n_1660), .Y(n_1746) );
NOR3xp33_ASAP7_75t_L g1752 ( .A(n_1564), .B(n_1618), .C(n_1709), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_1564), .B(n_1630), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1783 ( .A(n_1564), .B(n_1584), .Y(n_1783) );
NOR2xp33_ASAP7_75t_L g1794 ( .A(n_1564), .B(n_1607), .Y(n_1794) );
AND2x4_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1577), .Y(n_1564) );
AND2x4_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1572), .Y(n_1566) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
OR2x2_ASAP7_75t_L g1599 ( .A(n_1568), .B(n_1573), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1569), .B(n_1571), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1571), .Y(n_1580) );
AND2x4_ASAP7_75t_L g1574 ( .A(n_1572), .B(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
OR2x2_ASAP7_75t_L g1601 ( .A(n_1573), .B(n_1576), .Y(n_1601) );
HB1xp67_ASAP7_75t_L g1929 ( .A(n_1575), .Y(n_1929) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1578), .Y(n_1712) );
AND2x4_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1581), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1579), .B(n_1581), .Y(n_1589) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AND2x4_ASAP7_75t_L g1582 ( .A(n_1580), .B(n_1581), .Y(n_1582) );
INVx2_ASAP7_75t_L g1625 ( .A(n_1582), .Y(n_1625) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1583), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_1583), .A2(n_1734), .B1(n_1736), .B2(n_1739), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1753 ( .A(n_1583), .B(n_1622), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1587), .Y(n_1583) );
INVx1_ASAP7_75t_SL g1631 ( .A(n_1584), .Y(n_1631) );
CKINVDCx5p33_ASAP7_75t_R g1639 ( .A(n_1584), .Y(n_1639) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1584), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1584), .B(n_1640), .Y(n_1676) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1584), .Y(n_1703) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1584), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1585), .B(n_1586), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1587), .B(n_1631), .Y(n_1630) );
CKINVDCx6p67_ASAP7_75t_R g1640 ( .A(n_1587), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1587), .B(n_1657), .Y(n_1662) );
CKINVDCx5p33_ASAP7_75t_R g1698 ( .A(n_1587), .Y(n_1698) );
AOI221xp5_ASAP7_75t_L g1766 ( .A1(n_1587), .A2(n_1723), .B1(n_1767), .B2(n_1769), .C(n_1771), .Y(n_1766) );
OR2x6_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1590), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1607), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1593), .B(n_1610), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1593), .B(n_1609), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1593), .B(n_1682), .Y(n_1681) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1593), .B(n_1675), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1602), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1594), .B(n_1603), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1669 ( .A(n_1594), .B(n_1609), .Y(n_1669) );
INVx2_ASAP7_75t_L g1759 ( .A(n_1594), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1773 ( .A(n_1594), .B(n_1654), .Y(n_1773) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_1594), .B(n_1654), .Y(n_1799) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1595), .B(n_1603), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1595), .B(n_1602), .Y(n_1652) );
OAI22xp5_ASAP7_75t_L g1596 ( .A1(n_1597), .A2(n_1598), .B1(n_1600), .B2(n_1601), .Y(n_1596) );
OAI22xp33_ASAP7_75t_L g1604 ( .A1(n_1598), .A2(n_1601), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
OAI22xp33_ASAP7_75t_L g1626 ( .A1(n_1598), .A2(n_1627), .B1(n_1628), .B2(n_1629), .Y(n_1626) );
BUFx3_ASAP7_75t_L g1715 ( .A(n_1598), .Y(n_1715) );
BUFx6f_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
HB1xp67_ASAP7_75t_L g1629 ( .A(n_1601), .Y(n_1629) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1601), .Y(n_1718) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1603), .Y(n_1618) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1608), .B(n_1610), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1608), .B(n_1653), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1608), .B(n_1609), .Y(n_1724) );
NOR2x1_ASAP7_75t_L g1617 ( .A(n_1609), .B(n_1618), .Y(n_1617) );
OR2x2_ASAP7_75t_L g1658 ( .A(n_1609), .B(n_1659), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1609), .B(n_1688), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1609), .B(n_1618), .Y(n_1742) );
INVx2_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
BUFx3_ASAP7_75t_L g1654 ( .A(n_1610), .Y(n_1654) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_1610), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1610), .B(n_1618), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1610), .B(n_1652), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1612), .Y(n_1610) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
NOR2xp33_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
INVx2_ASAP7_75t_L g1637 ( .A(n_1615), .Y(n_1637) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_1615), .B(n_1660), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1668 ( .A(n_1615), .B(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1615), .B(n_1633), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1615), .B(n_1697), .Y(n_1696) );
OAI21xp5_ASAP7_75t_SL g1732 ( .A1(n_1615), .A2(n_1733), .B(n_1740), .Y(n_1732) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
OAI21xp33_ASAP7_75t_L g1670 ( .A1(n_1618), .A2(n_1671), .B(n_1673), .Y(n_1670) );
OR2x2_ASAP7_75t_L g1749 ( .A(n_1618), .B(n_1654), .Y(n_1749) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1630), .Y(n_1620) );
INVx2_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx2_ASAP7_75t_L g1644 ( .A(n_1622), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1622), .B(n_1710), .Y(n_1765) );
INVx2_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
INVx2_ASAP7_75t_SL g1657 ( .A(n_1623), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1623), .B(n_1640), .Y(n_1666) );
OR2x2_ASAP7_75t_L g1708 ( .A(n_1623), .B(n_1643), .Y(n_1708) );
INVx2_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1665 ( .A(n_1631), .B(n_1666), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1632), .B(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
NOR2xp33_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1641), .Y(n_1634) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1637), .B(n_1724), .Y(n_1723) );
OR2x2_ASAP7_75t_L g1748 ( .A(n_1637), .B(n_1749), .Y(n_1748) );
A2O1A1Ixp33_ASAP7_75t_L g1780 ( .A1(n_1637), .A2(n_1735), .B(n_1756), .C(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1638), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1640), .Y(n_1638) );
INVx3_ASAP7_75t_L g1643 ( .A(n_1639), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1639), .B(n_1656), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1639), .B(n_1723), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1726 ( .A(n_1639), .B(n_1727), .Y(n_1726) );
OAI32xp33_ASAP7_75t_L g1775 ( .A1(n_1639), .A2(n_1707), .A3(n_1724), .B1(n_1730), .B2(n_1776), .Y(n_1775) );
AND2x4_ASAP7_75t_SL g1656 ( .A(n_1640), .B(n_1657), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1692 ( .A(n_1640), .B(n_1657), .Y(n_1692) );
NOR2xp33_ASAP7_75t_L g1736 ( .A(n_1640), .B(n_1737), .Y(n_1736) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1640), .B(n_1738), .Y(n_1757) );
NAND3xp33_ASAP7_75t_L g1781 ( .A(n_1640), .B(n_1741), .C(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
OAI322xp33_ASAP7_75t_L g1786 ( .A1(n_1642), .A2(n_1655), .A3(n_1705), .B1(n_1708), .B2(n_1737), .C1(n_1787), .C2(n_1789), .Y(n_1786) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1685 ( .A(n_1643), .B(n_1686), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1768 ( .A(n_1643), .B(n_1657), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1643), .B(n_1651), .Y(n_1770) );
AOI21xp5_ASAP7_75t_L g1796 ( .A1(n_1643), .A2(n_1790), .B(n_1797), .Y(n_1796) );
NAND2xp5_ASAP7_75t_L g1778 ( .A(n_1644), .B(n_1710), .Y(n_1778) );
OAI221xp5_ASAP7_75t_SL g1645 ( .A1(n_1646), .A2(n_1655), .B1(n_1658), .B2(n_1661), .C(n_1663), .Y(n_1645) );
INVxp67_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1650), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1653), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1652), .B(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1652), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1653), .B(n_1660), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1654), .B(n_1730), .Y(n_1729) );
OR2x2_ASAP7_75t_L g1750 ( .A(n_1654), .B(n_1746), .Y(n_1750) );
NOR2xp33_ASAP7_75t_L g1747 ( .A(n_1655), .B(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
INVx2_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1662), .B(n_1703), .Y(n_1702) );
AOI21xp5_ASAP7_75t_L g1744 ( .A1(n_1662), .A2(n_1745), .B(n_1747), .Y(n_1744) );
AOI221xp5_ASAP7_75t_L g1663 ( .A1(n_1664), .A2(n_1667), .B1(n_1670), .B2(n_1676), .C(n_1677), .Y(n_1663) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1666), .Y(n_1731) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1676), .Y(n_1785) );
NOR2xp33_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1679), .Y(n_1677) );
NOR2xp33_ASAP7_75t_L g1784 ( .A(n_1679), .B(n_1785), .Y(n_1784) );
NAND4xp25_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1684), .C(n_1690), .D(n_1695), .Y(n_1680) );
O2A1O1Ixp33_ASAP7_75t_L g1793 ( .A1(n_1682), .A2(n_1687), .B(n_1794), .C(n_1795), .Y(n_1793) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1693), .Y(n_1690) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
AOI221xp5_ASAP7_75t_L g1695 ( .A1(n_1696), .A2(n_1698), .B1(n_1699), .B2(n_1702), .C(n_1704), .Y(n_1695) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1697), .Y(n_1727) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
AOI21xp33_ASAP7_75t_L g1704 ( .A1(n_1705), .A2(n_1706), .B(n_1708), .Y(n_1704) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
OAI221xp5_ASAP7_75t_SL g1743 ( .A1(n_1708), .A2(n_1737), .B1(n_1744), .B2(n_1750), .C(n_1751), .Y(n_1743) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
BUFx3_ASAP7_75t_L g1738 ( .A(n_1710), .Y(n_1738) );
O2A1O1Ixp33_ASAP7_75t_L g1779 ( .A1(n_1710), .A2(n_1780), .B(n_1784), .C(n_1786), .Y(n_1779) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
OAI22xp33_ASAP7_75t_L g1713 ( .A1(n_1714), .A2(n_1715), .B1(n_1716), .B2(n_1717), .Y(n_1713) );
HB1xp67_ASAP7_75t_L g1801 ( .A(n_1717), .Y(n_1801) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
NOR5xp2_ASAP7_75t_L g1719 ( .A(n_1720), .B(n_1732), .C(n_1743), .D(n_1754), .E(n_1758), .Y(n_1719) );
AOI31xp33_ASAP7_75t_L g1720 ( .A1(n_1721), .A2(n_1725), .A3(n_1728), .B(n_1731), .Y(n_1720) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1724), .Y(n_1735) );
OAI21xp33_ASAP7_75t_L g1751 ( .A1(n_1724), .A2(n_1752), .B(n_1753), .Y(n_1751) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
AOI31xp33_ASAP7_75t_L g1754 ( .A1(n_1728), .A2(n_1755), .A3(n_1756), .B(n_1757), .Y(n_1754) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
INVx2_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1753), .Y(n_1755) );
O2A1O1Ixp33_ASAP7_75t_L g1758 ( .A1(n_1759), .A2(n_1760), .B(n_1762), .C(n_1764), .Y(n_1758) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
OAI22xp5_ASAP7_75t_L g1795 ( .A1(n_1762), .A2(n_1764), .B1(n_1785), .B2(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
O2A1O1Ixp33_ASAP7_75t_SL g1771 ( .A1(n_1772), .A2(n_1774), .B(n_1775), .C(n_1778), .Y(n_1771) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
NOR2xp33_ASAP7_75t_L g1790 ( .A(n_1773), .B(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
INVxp67_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1798), .B(n_1799), .Y(n_1797) );
BUFx2_ASAP7_75t_SL g1800 ( .A(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
HB1xp67_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
AOI211xp5_ASAP7_75t_L g1806 ( .A1(n_1807), .A2(n_1823), .B(n_1824), .C(n_1848), .Y(n_1806) );
AOI22xp33_ASAP7_75t_L g1840 ( .A1(n_1811), .A2(n_1841), .B1(n_1843), .B2(n_1846), .Y(n_1840) );
AOI21xp5_ASAP7_75t_L g1815 ( .A1(n_1816), .A2(n_1817), .B(n_1818), .Y(n_1815) );
INVx1_ASAP7_75t_L g1819 ( .A(n_1820), .Y(n_1819) );
AOI31xp33_ASAP7_75t_L g1824 ( .A1(n_1825), .A2(n_1834), .A3(n_1840), .B(n_1847), .Y(n_1824) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
INVx2_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
AOI22xp33_ASAP7_75t_L g1834 ( .A1(n_1835), .A2(n_1836), .B1(n_1837), .B2(n_1839), .Y(n_1834) );
AND2x4_ASAP7_75t_L g1843 ( .A(n_1838), .B(n_1844), .Y(n_1843) );
INVx5_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
NAND4xp25_ASAP7_75t_L g1848 ( .A(n_1849), .B(n_1852), .C(n_1855), .D(n_1861), .Y(n_1848) );
NAND3xp33_ASAP7_75t_L g1855 ( .A(n_1856), .B(n_1857), .C(n_1858), .Y(n_1855) );
INVx3_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
NAND3xp33_ASAP7_75t_L g1861 ( .A(n_1862), .B(n_1863), .C(n_1864), .Y(n_1861) );
INVx1_ASAP7_75t_SL g1865 ( .A(n_1866), .Y(n_1865) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
BUFx2_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
OAI21xp5_ASAP7_75t_L g1928 ( .A1(n_1874), .A2(n_1929), .B(n_1930), .Y(n_1928) );
INVxp33_ASAP7_75t_SL g1875 ( .A(n_1876), .Y(n_1875) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1878), .Y(n_1877) );
HB1xp67_ASAP7_75t_L g1878 ( .A(n_1879), .Y(n_1878) );
NAND3xp33_ASAP7_75t_L g1879 ( .A(n_1880), .B(n_1885), .C(n_1901), .Y(n_1879) );
NOR2xp33_ASAP7_75t_L g1880 ( .A(n_1881), .B(n_1883), .Y(n_1880) );
NOR2xp33_ASAP7_75t_L g1885 ( .A(n_1886), .B(n_1887), .Y(n_1885) );
AOI22xp33_ASAP7_75t_L g1906 ( .A1(n_1895), .A2(n_1899), .B1(n_1907), .B2(n_1909), .Y(n_1906) );
BUFx2_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
OAI22xp5_ASAP7_75t_L g1914 ( .A1(n_1915), .A2(n_1917), .B1(n_1920), .B2(n_1923), .Y(n_1914) );
INVx1_ASAP7_75t_L g1918 ( .A(n_1919), .Y(n_1918) );
BUFx2_ASAP7_75t_L g1927 ( .A(n_1928), .Y(n_1927) );
endmodule