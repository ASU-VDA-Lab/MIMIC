module fake_jpeg_2807_n_510 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_22),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_63),
.Y(n_152)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_16),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_82),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_0),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g122 ( 
.A(n_87),
.Y(n_122)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_26),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_99),
.Y(n_146)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_26),
.C(n_34),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_27),
.C(n_45),
.Y(n_173)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_59),
.B1(n_69),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_117),
.A2(n_135),
.B1(n_31),
.B2(n_35),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_36),
.B(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_24),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_52),
.B(n_22),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_132),
.B(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_53),
.A2(n_21),
.B1(n_40),
.B2(n_24),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_40),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_101),
.A2(n_27),
.B1(n_21),
.B2(n_34),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_76),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_158),
.B(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_61),
.B(n_70),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_163),
.B(n_207),
.Y(n_234)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_169),
.B(n_173),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_120),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_170),
.Y(n_237)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_102),
.A2(n_70),
.B1(n_65),
.B2(n_99),
.Y(n_177)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_107),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_185),
.B(n_187),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_65),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_188),
.B(n_191),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_56),
.B1(n_84),
.B2(n_37),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_201),
.B(n_20),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_118),
.A2(n_35),
.B1(n_31),
.B2(n_20),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_210),
.B1(n_211),
.B2(n_37),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_63),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_95),
.B1(n_83),
.B2(n_90),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_205),
.B1(n_36),
.B2(n_50),
.Y(n_228)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_247)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_108),
.A2(n_41),
.B1(n_25),
.B2(n_39),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_206),
.Y(n_216)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_107),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_108),
.B(n_99),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_129),
.C(n_123),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_140),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_177),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_128),
.A2(n_20),
.B1(n_35),
.B2(n_36),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_150),
.A2(n_43),
.B1(n_71),
.B2(n_100),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_109),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_219),
.B(n_186),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_129),
.B(n_122),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_238),
.B(n_242),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_228),
.A2(n_235),
.B1(n_238),
.B2(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_153),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_251),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_162),
.A2(n_151),
.B1(n_155),
.B2(n_170),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_191),
.A2(n_37),
.B(n_23),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_239),
.A2(n_50),
.B1(n_45),
.B2(n_41),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_188),
.A2(n_122),
.B1(n_141),
.B2(n_136),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_189),
.A2(n_80),
.B1(n_81),
.B2(n_93),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_192),
.B1(n_172),
.B2(n_204),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_173),
.B(n_152),
.C(n_156),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_259),
.C(n_177),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_194),
.A2(n_121),
.B(n_98),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_121),
.B(n_39),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_153),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_257),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_182),
.B(n_41),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_168),
.B(n_121),
.C(n_96),
.Y(n_259)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_279),
.B1(n_288),
.B2(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_261),
.B1(n_255),
.B2(n_244),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_265),
.A2(n_286),
.B1(n_294),
.B2(n_302),
.Y(n_333)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_304),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_260),
.B1(n_220),
.B2(n_230),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_269),
.A2(n_276),
.B1(n_298),
.B2(n_8),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_227),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_285),
.C(n_23),
.Y(n_330)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_277),
.Y(n_325)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_228),
.A2(n_211),
.B1(n_164),
.B2(n_167),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_280),
.B(n_281),
.Y(n_334)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_291),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_232),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_174),
.B1(n_215),
.B2(n_180),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_175),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_289),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_222),
.A2(n_196),
.B1(n_203),
.B2(n_176),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_199),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_241),
.B(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_226),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_300),
.B(n_232),
.C(n_258),
.D(n_262),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_181),
.B1(n_195),
.B2(n_213),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_219),
.A2(n_144),
.B1(n_197),
.B2(n_200),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_299),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_45),
.B1(n_25),
.B2(n_38),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_257),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_242),
.A2(n_144),
.B1(n_160),
.B2(n_161),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_256),
.B1(n_218),
.B2(n_262),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_165),
.B1(n_39),
.B2(n_50),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_267),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_217),
.B(n_166),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_305),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_338)
);

AO22x1_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_258),
.B1(n_240),
.B2(n_229),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_312),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_248),
.C(n_251),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_337),
.C(n_340),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_236),
.B1(n_233),
.B2(n_232),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g373 ( 
.A1(n_309),
.A2(n_317),
.B(n_318),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_313),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_247),
.B(n_243),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_314),
.A2(n_294),
.B(n_275),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_272),
.A2(n_233),
.B1(n_241),
.B2(n_218),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_252),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_319),
.B(n_336),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_328),
.B1(n_335),
.B2(n_344),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_322),
.B(n_331),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_273),
.A2(n_254),
.B1(n_245),
.B2(n_38),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_324),
.A2(n_332),
.B(n_341),
.Y(n_351)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_265),
.A2(n_254),
.B1(n_38),
.B2(n_25),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_8),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_286),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_299),
.A2(n_283),
.B1(n_266),
.B2(n_281),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_283),
.A2(n_23),
.B1(n_33),
.B2(n_2),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_0),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_268),
.B(n_1),
.C(n_3),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_263),
.B1(n_301),
.B2(n_303),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_266),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_288),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_3),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_278),
.A2(n_4),
.B(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_332),
.A2(n_280),
.B1(n_264),
.B2(n_279),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_348),
.A2(n_350),
.B1(n_333),
.B2(n_316),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_360),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_352),
.B(n_366),
.Y(n_388)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_284),
.C(n_291),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_336),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_358),
.A2(n_324),
.B1(n_309),
.B2(n_320),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_302),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_297),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_328),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_365),
.Y(n_389)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_311),
.B(n_295),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_343),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_318),
.A2(n_314),
.B(n_312),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_340),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_339),
.A2(n_292),
.B(n_9),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_369),
.A2(n_341),
.B(n_306),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_8),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_8),
.Y(n_374)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_375),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_379),
.B(n_396),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_380),
.A2(n_384),
.B1(n_390),
.B2(n_401),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_382),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_348),
.A2(n_333),
.B1(n_316),
.B2(n_306),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_386),
.B(n_349),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_308),
.C(n_337),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_356),
.C(n_345),
.Y(n_424)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_356),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_345),
.A2(n_335),
.B1(n_313),
.B2(n_325),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_364),
.A2(n_325),
.B1(n_321),
.B2(n_338),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_403),
.A2(n_404),
.B1(n_406),
.B2(n_362),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_364),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_357),
.B(n_10),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_349),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_354),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_388),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_407),
.B(n_422),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_418),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_411),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_361),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_391),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_419),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_387),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_421),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_389),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_392),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_395),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_377),
.C(n_368),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_427),
.C(n_428),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_351),
.C(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_351),
.C(n_359),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_429),
.B(n_374),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_380),
.B(n_365),
.C(n_370),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_404),
.C(n_403),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_384),
.A2(n_346),
.B1(n_358),
.B2(n_373),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_373),
.B(n_389),
.Y(n_433)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_381),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_405),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_408),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_418),
.C(n_424),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_441),
.B(n_443),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_395),
.C(n_398),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_427),
.C(n_412),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_423),
.C(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_409),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_450),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_393),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_452),
.B(n_460),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_454),
.B(n_449),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_459),
.Y(n_469)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_435),
.Y(n_457)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_457),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_426),
.C(n_398),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_438),
.B(n_355),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_419),
.C(n_381),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_450),
.C(n_434),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_465),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_442),
.A2(n_406),
.B1(n_385),
.B2(n_392),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_375),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_385),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_467),
.Y(n_474)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_437),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_445),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_473),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_463),
.A2(n_442),
.B1(n_432),
.B2(n_436),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_472),
.A2(n_477),
.B1(n_478),
.B2(n_458),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_453),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_479),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_454),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_456),
.A2(n_440),
.B1(n_434),
.B2(n_446),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_455),
.A2(n_444),
.B1(n_439),
.B2(n_375),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_375),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_481),
.A2(n_464),
.B(n_461),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_469),
.B(n_462),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_487),
.B(n_488),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_483),
.B(n_490),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_492),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_486),
.A2(n_476),
.B(n_14),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_458),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_480),
.A2(n_468),
.B(n_474),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_477),
.B(n_11),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_473),
.B(n_12),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_12),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_12),
.Y(n_492)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_489),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_496),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_471),
.C(n_481),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_483),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_499),
.B(n_484),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_501),
.A2(n_503),
.B(n_497),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_497),
.C(n_494),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_505),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_502),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_15),
.C(n_13),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_14),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_509),
.B(n_15),
.Y(n_510)
);


endmodule