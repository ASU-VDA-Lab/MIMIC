module fake_netlist_6_4014_n_186 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_186);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_186;

wire n_52;
wire n_91;
wire n_146;
wire n_46;
wire n_119;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_5),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_29),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_1),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_32),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_49),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_47),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_45),
.B1(n_52),
.B2(n_36),
.C(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_54),
.Y(n_79)
);

OAI221xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_52),
.B1(n_36),
.B2(n_40),
.C(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_44),
.B1(n_14),
.B2(n_19),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_8),
.C(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_24),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_56),
.Y(n_90)
);

OAI221xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_72),
.B1(n_71),
.B2(n_74),
.C(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_67),
.B(n_74),
.Y(n_93)
);

NAND2x1p5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_76),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_76),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_59),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_66),
.B(n_68),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_66),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_66),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_92),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_80),
.B(n_84),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_83),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_83),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

OR2x6_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_98),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_101),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_77),
.Y(n_118)
);

NAND4xp25_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_58),
.C(n_91),
.D(n_97),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_114),
.Y(n_120)
);

O2A1O1Ixp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_106),
.B(n_98),
.C(n_115),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_111),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_118),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_107),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_125),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_135),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_148),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_133),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_130),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_128),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_147),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_155),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_99),
.C(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

HAxp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_99),
.CON(n_168),
.SN(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_159),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_162),
.B1(n_158),
.B2(n_68),
.C(n_58),
.Y(n_171)
);

AND4x1_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_105),
.C(n_102),
.D(n_68),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_119),
.C(n_58),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_68),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_112),
.C(n_107),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_166),
.B(n_107),
.C(n_93),
.Y(n_177)
);

AND3x1_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_112),
.C(n_107),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_169),
.B1(n_112),
.B2(n_100),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_171),
.A2(n_112),
.B(n_100),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_112),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.C(n_177),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_182),
.B(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_172),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_100),
.B1(n_183),
.B2(n_184),
.Y(n_186)
);


endmodule