module fake_jpeg_21863_n_305 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_8),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_25),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_28),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_65),
.Y(n_84)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_34),
.B2(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_22),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_17),
.Y(n_63)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_25),
.B1(n_34),
.B2(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_68),
.B1(n_42),
.B2(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_33),
.B1(n_22),
.B2(n_26),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_33),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_82),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_68),
.B1(n_86),
.B2(n_65),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_28),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_42),
.B1(n_32),
.B2(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_29),
.B1(n_18),
.B2(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_61),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_45),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_85),
.C(n_53),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_114),
.B1(n_88),
.B2(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_110),
.B1(n_29),
.B2(n_20),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_119),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_61),
.B1(n_35),
.B2(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_120),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_64),
.B1(n_35),
.B2(n_36),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_64),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_41),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_79),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_140),
.B1(n_98),
.B2(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_75),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_119),
.C(n_100),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_108),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_148),
.B(n_38),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_64),
.B1(n_51),
.B2(n_54),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_70),
.B1(n_90),
.B2(n_78),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_91),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_19),
.B(n_23),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_79),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_27),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_27),
.B1(n_26),
.B2(n_16),
.C(n_9),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_186)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_159),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_158),
.C(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_120),
.C(n_95),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_118),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_176),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_95),
.B1(n_97),
.B2(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_160),
.B1(n_156),
.B2(n_180),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_97),
.B(n_98),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_142),
.B(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_171),
.B1(n_179),
.B2(n_140),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_102),
.C(n_46),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_102),
.B(n_30),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_167),
.B(n_168),
.C(n_149),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_143),
.B1(n_137),
.B2(n_131),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_70),
.B1(n_92),
.B2(n_47),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_26),
.B(n_92),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_38),
.C(n_41),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_144),
.C(n_124),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_0),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_175),
.B(n_38),
.Y(n_202)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_145),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_70),
.B1(n_44),
.B2(n_56),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_184),
.Y(n_211)
);

INVxp33_ASAP7_75t_SL g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_136),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_195),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_194),
.B1(n_201),
.B2(n_190),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_123),
.B1(n_150),
.B2(n_141),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_175),
.B1(n_151),
.B2(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

OA21x2_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_202),
.B(n_167),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_134),
.B1(n_150),
.B2(n_124),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_136),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_204),
.C(n_205),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_135),
.B1(n_23),
.B2(n_19),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_38),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_41),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_41),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_178),
.C(n_163),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_173),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_210),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_216),
.B1(n_219),
.B2(n_8),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_162),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_223),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_227),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_162),
.B1(n_152),
.B2(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_226),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

AOI321xp33_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_152),
.A3(n_174),
.B1(n_161),
.B2(n_12),
.C(n_4),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_174),
.C(n_59),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_229),
.C(n_23),
.Y(n_242)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_59),
.C(n_56),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_191),
.B1(n_201),
.B2(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_235),
.B1(n_237),
.B2(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_191),
.B1(n_204),
.B2(n_90),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_78),
.B1(n_56),
.B2(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_240),
.B(n_245),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_23),
.B(n_44),
.C(n_78),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_207),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_0),
.B(n_1),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_233),
.A2(n_222),
.B1(n_210),
.B2(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_251),
.A2(n_257),
.B1(n_10),
.B2(n_5),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_212),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_259),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_208),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_220),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_11),
.C(n_6),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_225),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_241),
.C(n_231),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_220),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_244),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_234),
.B(n_233),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_272),
.B(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_259),
.B(n_11),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_SL g269 ( 
.A(n_264),
.B(n_251),
.C(n_246),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_260),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_237),
.B(n_3),
.C(n_2),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_275),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_14),
.B1(n_7),
.B2(n_10),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_280),
.B(n_286),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_272),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_14),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_14),
.B(n_15),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_271),
.C(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_271),
.C(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_3),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_298),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_15),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_16),
.B(n_288),
.C(n_287),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_292),
.B(n_16),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_295),
.C(n_302),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_301),
.Y(n_305)
);


endmodule