module fake_jpeg_2643_n_222 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_59),
.Y(n_88)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_58),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_69),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_66),
.B1(n_54),
.B2(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_67),
.B1(n_66),
.B2(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_68),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_109),
.Y(n_120)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_67),
.B1(n_85),
.B2(n_60),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_85),
.B1(n_81),
.B2(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_71),
.B1(n_60),
.B2(n_57),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2x1_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_131),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_65),
.B(n_77),
.C(n_61),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_130),
.B(n_70),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_71),
.B1(n_63),
.B2(n_86),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_134),
.B1(n_135),
.B2(n_121),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_138),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_65),
.B(n_53),
.C(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_99),
.B1(n_83),
.B2(n_84),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_86),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_57),
.CI(n_70),
.CON(n_136),
.SN(n_136)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_6),
.B(n_7),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_86),
.B1(n_57),
.B2(n_70),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_75),
.B1(n_26),
.B2(n_28),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_106),
.B1(n_103),
.B2(n_116),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_36),
.B(n_46),
.C(n_45),
.Y(n_179)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_141),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_146),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_75),
.B1(n_3),
.B2(n_4),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_154),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_29),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g155 ( 
.A1(n_136),
.A2(n_2),
.B(n_5),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_8),
.B(n_9),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_10),
.C(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_33),
.B1(n_51),
.B2(n_50),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_8),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_176),
.Y(n_185)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_180),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_133),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_172),
.B(n_179),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_10),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_32),
.C(n_48),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_168),
.C(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_151),
.B(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_187),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_153),
.B(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_183),
.B(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_174),
.B(n_167),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_25),
.B(n_43),
.C(n_41),
.D(n_40),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_21),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_166),
.C(n_172),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_166),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_173),
.B1(n_168),
.B2(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_52),
.B1(n_38),
.B2(n_37),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_179),
.B1(n_189),
.B2(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_179),
.C(n_23),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_208),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.C(n_194),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_206),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_195),
.Y(n_216)
);

AOI31xp67_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_214),
.A3(n_210),
.B(n_207),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_30),
.B1(n_13),
.B2(n_16),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_12),
.C(n_16),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_17),
.B(n_18),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_17),
.B(n_18),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);


endmodule