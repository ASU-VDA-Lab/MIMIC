module fake_jpeg_28614_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_16),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_66),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_42),
.Y(n_83)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_26),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_39),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_6),
.B(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_30),
.B1(n_38),
.B2(n_35),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_94),
.B1(n_113),
.B2(n_65),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_30),
.B1(n_38),
.B2(n_35),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_125),
.B1(n_58),
.B2(n_46),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_60),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_32),
.B(n_27),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_6),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_47),
.A2(n_37),
.B1(n_38),
.B2(n_35),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_38),
.B1(n_35),
.B2(n_23),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_123),
.B1(n_127),
.B2(n_92),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_57),
.B(n_41),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_14),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_63),
.A2(n_23),
.B1(n_33),
.B2(n_31),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_79),
.A2(n_33),
.B1(n_31),
.B2(n_23),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_59),
.B1(n_78),
.B2(n_72),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_129),
.A2(n_133),
.B1(n_142),
.B2(n_150),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_146),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_132),
.B(n_135),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_71),
.B1(n_77),
.B2(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_70),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_102),
.B1(n_108),
.B2(n_153),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_88),
.A2(n_68),
.B1(n_64),
.B2(n_52),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_116),
.B1(n_120),
.B2(n_118),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_51),
.B1(n_48),
.B2(n_53),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_70),
.B(n_73),
.C(n_75),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_145),
.A2(n_147),
.B(n_154),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_81),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_34),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_101),
.B(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_85),
.A2(n_34),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_110),
.B1(n_106),
.B2(n_121),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_102),
.B1(n_108),
.B2(n_170),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_34),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_159),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_6),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_84),
.B(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_161),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_89),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_89),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_12),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_12),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_13),
.C(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_13),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_14),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_141),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_128),
.B1(n_116),
.B2(n_100),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_171),
.B1(n_108),
.B2(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_127),
.B1(n_120),
.B2(n_112),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_111),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_145),
.B1(n_158),
.B2(n_167),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_124),
.C(n_118),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_180),
.B(n_184),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_124),
.C(n_108),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_193),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_208),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_201),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_130),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_204),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_156),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_165),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_214),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_187),
.A2(n_154),
.B1(n_143),
.B2(n_142),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_216),
.B(n_203),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_176),
.B1(n_209),
.B2(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_132),
.B1(n_139),
.B2(n_154),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_235),
.B1(n_239),
.B2(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_164),
.B1(n_142),
.B2(n_167),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_142),
.B1(n_167),
.B2(n_166),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_223),
.B(n_238),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_157),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_161),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_170),
.B1(n_140),
.B2(n_168),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_229),
.B(n_212),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_191),
.A2(n_201),
.B1(n_192),
.B2(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_162),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_167),
.B1(n_169),
.B2(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_144),
.B1(n_205),
.B2(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_144),
.Y(n_240)
);

AO21x2_ASAP7_75t_SL g241 ( 
.A1(n_192),
.A2(n_200),
.B(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_173),
.B(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_173),
.B(n_184),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_200),
.A2(n_193),
.B1(n_174),
.B2(n_183),
.Y(n_246)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_174),
.C(n_185),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_255),
.C(n_261),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_183),
.B1(n_185),
.B2(n_189),
.C(n_198),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_275),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_181),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_257),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_189),
.C(n_182),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_222),
.A2(n_197),
.B(n_182),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_260),
.B(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_181),
.C(n_199),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_276),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_231),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_203),
.C(n_207),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_228),
.B(n_207),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_248),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_212),
.B1(n_196),
.B2(n_190),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_234),
.B1(n_236),
.B2(n_231),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_196),
.C(n_226),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_246),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_228),
.A2(n_215),
.B(n_218),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_219),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_235),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_247),
.B(n_217),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_236),
.C(n_218),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_214),
.B1(n_221),
.B2(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_285),
.B(n_305),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_277),
.B1(n_267),
.B2(n_253),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_241),
.B1(n_238),
.B2(n_233),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_276),
.B(n_278),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_233),
.C(n_232),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_296),
.Y(n_329)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_280),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_213),
.Y(n_298)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_243),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_302),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_237),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_271),
.B(n_242),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_273),
.C(n_261),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_310),
.C(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_273),
.C(n_255),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_312),
.B(n_259),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_324),
.B1(n_283),
.B2(n_252),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_272),
.C(n_267),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_291),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_325),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_251),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_293),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_241),
.B1(n_274),
.B2(n_278),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_256),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_268),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_293),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_335),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_298),
.C(n_281),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_316),
.C(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_304),
.CI(n_290),
.CON(n_338),
.SN(n_338)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_287),
.B1(n_282),
.B2(n_301),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_340),
.B1(n_348),
.B2(n_349),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_329),
.A2(n_286),
.B1(n_282),
.B2(n_262),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_346),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_342),
.A2(n_350),
.B1(n_283),
.B2(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_344),
.Y(n_353)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_259),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_SL g349 ( 
.A(n_314),
.B(n_257),
.C(n_283),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_309),
.A2(n_284),
.B1(n_295),
.B2(n_289),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_345),
.A2(n_319),
.B(n_313),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_351),
.A2(n_337),
.B(n_258),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_354),
.B(n_362),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_322),
.C(n_258),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_356),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_342),
.A2(n_309),
.B(n_324),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_SL g359 ( 
.A(n_334),
.B(n_311),
.C(n_308),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_365),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_311),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_332),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_310),
.C(n_325),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_327),
.B1(n_321),
.B2(n_331),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_366),
.B(n_341),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_376),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_369),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_335),
.Y(n_369)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_336),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_371),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_361),
.B(n_346),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_375),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_327),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_372),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_387),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_377),
.A2(n_363),
.B1(n_365),
.B2(n_358),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_374),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_377),
.A2(n_352),
.B1(n_357),
.B2(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_299),
.B1(n_284),
.B2(n_288),
.Y(n_396)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_352),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_388),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_367),
.A2(n_353),
.B1(n_366),
.B2(n_318),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_389),
.A2(n_355),
.B1(n_338),
.B2(n_300),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_392),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_384),
.A2(n_369),
.B1(n_354),
.B2(n_338),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_395),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_394),
.A2(n_396),
.B1(n_385),
.B2(n_383),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_379),
.B(n_383),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_399),
.B(n_397),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_400),
.B(n_402),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_266),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_405),
.B(n_401),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_407),
.C(n_382),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_403),
.A2(n_399),
.B(n_394),
.Y(n_407)
);

NAND4xp25_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_382),
.C(n_380),
.D(n_279),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_380),
.B(n_242),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_410),
.B(n_248),
.Y(n_411)
);


endmodule