module fake_jpeg_804_n_48 (n_3, n_2, n_1, n_0, n_4, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_14),
.Y(n_21)
);

AO22x2_ASAP7_75t_L g13 ( 
.A1(n_7),
.A2(n_8),
.B1(n_10),
.B2(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_20),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_13),
.B(n_16),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.C(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_12),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_13),
.B(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_21),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_24),
.C(n_13),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_32),
.C(n_20),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_13),
.B(n_20),
.Y(n_36)
);

OAI21x1_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_4),
.C(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_9),
.B1(n_8),
.B2(n_4),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_42),
.B2(n_1),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_8),
.C(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_46),
.B(n_42),
.Y(n_47)
);

NOR2xp67_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_2),
.Y(n_48)
);


endmodule