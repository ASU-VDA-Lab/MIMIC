module fake_jpeg_28916_n_429 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_53),
.Y(n_94)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_86),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_24),
.B(n_15),
.CON(n_58),
.SN(n_58)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_58),
.B(n_3),
.Y(n_119)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_70),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_79),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_43),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_25),
.B(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_27),
.B1(n_43),
.B2(n_30),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_87),
.A2(n_100),
.B1(n_122),
.B2(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_103),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_58),
.B1(n_27),
.B2(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_132),
.B1(n_67),
.B2(n_37),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_28),
.B1(n_41),
.B2(n_39),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_28),
.B1(n_41),
.B2(n_39),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_119),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_47),
.B1(n_51),
.B2(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_38),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_31),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_74),
.A2(n_40),
.B1(n_35),
.B2(n_32),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

NAND2x1_ASAP7_75t_SL g193 ( 
.A(n_136),
.B(n_163),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_76),
.B1(n_75),
.B2(n_65),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_91),
.A2(n_59),
.B1(n_35),
.B2(n_32),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_173),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_63),
.B1(n_62),
.B2(n_60),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_145),
.B(n_166),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_95),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_45),
.B1(n_52),
.B2(n_30),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_108),
.Y(n_151)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_133),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_162),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_56),
.A3(n_57),
.B1(n_70),
.B2(n_40),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_172),
.Y(n_186)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_100),
.B(n_40),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_56),
.C(n_35),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_105),
.B(n_35),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_32),
.C(n_4),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_87),
.C(n_8),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_32),
.B(n_4),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_94),
.B(n_4),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_95),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_118),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_194),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_176),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_207),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_129),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_96),
.B1(n_98),
.B2(n_92),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_155),
.B(n_141),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_104),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_104),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_117),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_215),
.B(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_146),
.B1(n_140),
.B2(n_147),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_230),
.B1(n_206),
.B2(n_93),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_158),
.B1(n_154),
.B2(n_166),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_238),
.B1(n_248),
.B2(n_105),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_200),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_225),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_173),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_228),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_205),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_206),
.B1(n_186),
.B2(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_196),
.B(n_146),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_236),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_188),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_146),
.B(n_163),
.C(n_151),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_247),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_235),
.Y(n_268)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_164),
.B1(n_169),
.B2(n_174),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_192),
.A2(n_162),
.B1(n_165),
.B2(n_96),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_243),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_241),
.B(n_242),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_152),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

AO21x2_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_206),
.B(n_122),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_210),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_207),
.C(n_190),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_263),
.C(n_242),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_193),
.B(n_198),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_250),
.A2(n_277),
.B(n_209),
.Y(n_305)
);

AO22x1_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_246),
.B1(n_233),
.B2(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_253),
.B(n_217),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_266),
.B1(n_272),
.B2(n_243),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_177),
.B1(n_120),
.B2(n_116),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_262),
.B1(n_267),
.B2(n_273),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_120),
.B1(n_116),
.B2(n_208),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_182),
.C(n_139),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_218),
.A2(n_137),
.B1(n_138),
.B2(n_208),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_93),
.B1(n_111),
.B2(n_98),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_230),
.A2(n_111),
.B1(n_106),
.B2(n_113),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_113),
.B1(n_197),
.B2(n_201),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_199),
.B(n_195),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_280),
.A2(n_281),
.B1(n_292),
.B2(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_265),
.C(n_182),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_285),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_239),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_286),
.Y(n_323)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_291),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_258),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_306),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_239),
.B1(n_231),
.B2(n_234),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_294),
.B1(n_295),
.B2(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_257),
.A2(n_242),
.B1(n_216),
.B2(n_219),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_216),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_259),
.A2(n_227),
.B1(n_219),
.B2(n_229),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_222),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_249),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_266),
.A2(n_220),
.B1(n_224),
.B2(n_232),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_252),
.B(n_235),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_298),
.B(n_300),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_273),
.A2(n_221),
.B1(n_228),
.B2(n_245),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_304),
.B1(n_274),
.B2(n_268),
.Y(n_316)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_213),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_301),
.B(n_302),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_228),
.B1(n_221),
.B2(n_195),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_201),
.B1(n_209),
.B2(n_236),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_277),
.B(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

NAND2x1_ASAP7_75t_SL g333 ( 
.A(n_307),
.B(n_308),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_269),
.B(n_260),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_264),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_309),
.B(n_312),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_264),
.B(n_271),
.C(n_263),
.D(n_251),
.Y(n_313)
);

AOI211xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_161),
.B(n_168),
.C(n_171),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_316),
.A2(n_317),
.B1(n_325),
.B2(n_281),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_251),
.B1(n_276),
.B2(n_260),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_264),
.C(n_267),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_324),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_251),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_251),
.B1(n_276),
.B2(n_262),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_292),
.C(n_285),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_270),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_282),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_280),
.B(n_274),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_331),
.A2(n_286),
.B1(n_291),
.B2(n_287),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_302),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_337),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_321),
.A2(n_280),
.B1(n_288),
.B2(n_300),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_340),
.B1(n_352),
.B2(n_311),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_350),
.C(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_330),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_339),
.B(n_348),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_321),
.A2(n_306),
.B1(n_294),
.B2(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_347),
.Y(n_354)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_351),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_318),
.B(n_270),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_310),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_315),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_303),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_106),
.B1(n_112),
.B2(n_157),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_356),
.C(n_357),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_308),
.C(n_320),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_313),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_323),
.B1(n_307),
.B2(n_346),
.Y(n_378)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_350),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_320),
.C(n_331),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_370),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_371),
.B(n_378),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_368),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_383),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_356),
.A2(n_333),
.B(n_351),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_376),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_332),
.B1(n_333),
.B2(n_324),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_316),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_380),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_363),
.A2(n_340),
.B1(n_311),
.B2(n_325),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_360),
.B1(n_355),
.B2(n_354),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_352),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_364),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_369),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_317),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_353),
.C(n_385),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_389),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_359),
.B1(n_355),
.B2(n_354),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_391),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_375),
.Y(n_392)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_392),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_365),
.C(n_357),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_396),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_345),
.B(n_309),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_112),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_398),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_387),
.B(n_381),
.Y(n_400)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_400),
.Y(n_415)
);

AOI31xp33_ASAP7_75t_L g403 ( 
.A1(n_393),
.A2(n_383),
.A3(n_161),
.B(n_10),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g412 ( 
.A1(n_403),
.A2(n_11),
.B(n_13),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_393),
.A2(n_5),
.B(n_9),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_11),
.B(n_13),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_388),
.A2(n_99),
.B1(n_10),
.B2(n_11),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_9),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_99),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_11),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_412),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_398),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_414),
.B(n_399),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_413),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_416),
.A2(n_406),
.B(n_407),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_399),
.Y(n_417)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_405),
.C(n_408),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_419),
.A2(n_422),
.B(n_415),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_420),
.B(n_411),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_424),
.B(n_421),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_418),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_394),
.C(n_396),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_14),
.B(n_15),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_14),
.Y(n_429)
);


endmodule