module real_aes_2475_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_637;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_0), .A2(n_189), .B1(n_429), .B2(n_430), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_1), .A2(n_155), .B1(n_382), .B2(n_383), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_2), .A2(n_195), .B1(n_314), .B2(n_393), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_3), .A2(n_125), .B1(n_493), .B2(n_622), .Y(n_621) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_4), .A2(n_143), .B1(n_238), .B2(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g633 ( .A(n_4), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_5), .A2(n_90), .B1(n_315), .B2(n_453), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_6), .A2(n_191), .B1(n_382), .B2(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_7), .A2(n_144), .B1(n_383), .B2(n_534), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_8), .A2(n_62), .B1(n_494), .B2(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_9), .A2(n_162), .B1(n_299), .B2(n_305), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_10), .B(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_11), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_12), .Y(n_561) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_13), .A2(n_52), .B1(n_238), .B2(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_13), .B(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_14), .A2(n_171), .B1(n_305), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_15), .A2(n_71), .B1(n_422), .B2(n_423), .Y(n_421) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_16), .A2(n_138), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_17), .A2(n_168), .B1(n_401), .B2(n_571), .Y(n_570) );
AO222x2_ASAP7_75t_SL g531 ( .A1(n_18), .A2(n_37), .B1(n_119), .B2(n_415), .C1(n_418), .C2(n_419), .Y(n_531) );
AO22x2_ASAP7_75t_L g467 ( .A1(n_19), .A2(n_468), .B1(n_495), .B2(n_496), .Y(n_467) );
INVx1_ASAP7_75t_L g496 ( .A(n_19), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_20), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_21), .A2(n_70), .B1(n_432), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_22), .A2(n_205), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_23), .A2(n_98), .B1(n_476), .B2(n_490), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_24), .A2(n_115), .B1(n_425), .B2(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_25), .B(n_330), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_26), .A2(n_156), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_27), .A2(n_157), .B1(n_333), .B2(n_386), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_28), .A2(n_123), .B1(n_436), .B2(n_437), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_29), .A2(n_188), .B1(n_332), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_30), .A2(n_116), .B1(n_393), .B2(n_432), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_31), .A2(n_97), .B1(n_380), .B2(n_486), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_32), .A2(n_164), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_33), .A2(n_124), .B1(n_476), .B2(n_477), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_34), .A2(n_159), .B1(n_382), .B2(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_35), .A2(n_103), .B1(n_379), .B2(n_380), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_36), .A2(n_93), .B1(n_264), .B2(n_365), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_38), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_39), .A2(n_192), .B1(n_289), .B2(n_294), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_40), .A2(n_63), .B1(n_430), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_41), .A2(n_194), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_42), .A2(n_91), .B1(n_320), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_43), .A2(n_74), .B1(n_422), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_44), .A2(n_88), .B1(n_383), .B2(n_534), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_45), .A2(n_193), .B1(n_321), .B2(n_453), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_46), .A2(n_183), .B1(n_398), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_47), .A2(n_137), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_48), .A2(n_100), .B1(n_422), .B2(n_536), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_49), .A2(n_128), .B1(n_400), .B2(n_401), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_50), .A2(n_113), .B1(n_418), .B2(n_419), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_51), .A2(n_199), .B1(n_403), .B2(n_404), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_53), .A2(n_151), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_54), .A2(n_196), .B1(n_360), .B2(n_521), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_55), .A2(n_637), .B1(n_638), .B2(n_655), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_55), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_56), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_57), .A2(n_170), .B1(n_493), .B2(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g230 ( .A(n_58), .B(n_231), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_59), .A2(n_95), .B1(n_397), .B2(n_398), .Y(n_396) );
OA22x2_ASAP7_75t_L g548 ( .A1(n_60), .A2(n_549), .B1(n_550), .B2(n_573), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_60), .Y(n_549) );
INVx3_ASAP7_75t_L g238 ( .A(n_61), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_64), .A2(n_111), .B1(n_400), .B2(n_401), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_65), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_66), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_67), .A2(n_163), .B1(n_343), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_68), .A2(n_175), .B1(n_418), .B2(n_419), .Y(n_586) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_69), .A2(n_78), .B1(n_145), .B2(n_445), .C1(n_555), .C2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_72), .A2(n_185), .B1(n_429), .B2(n_430), .Y(n_572) );
INVx1_ASAP7_75t_SL g239 ( .A(n_73), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_73), .B(n_101), .Y(n_634) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_75), .A2(n_122), .B1(n_251), .B2(n_257), .Y(n_250) );
AOI22xp5_ASAP7_75t_SL g613 ( .A1(n_76), .A2(n_160), .B1(n_614), .B2(n_615), .Y(n_613) );
INVx2_ASAP7_75t_L g214 ( .A(n_77), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_79), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_80), .A2(n_105), .B1(n_418), .B2(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_81), .A2(n_112), .B1(n_400), .B2(n_401), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_82), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_83), .A2(n_110), .B1(n_310), .B2(n_313), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_84), .A2(n_96), .B1(n_317), .B2(n_320), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_85), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_86), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_87), .A2(n_139), .B1(n_429), .B2(n_430), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_89), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_92), .A2(n_187), .B1(n_264), .B2(n_606), .Y(n_651) );
INVx1_ASAP7_75t_L g225 ( .A(n_94), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_99), .A2(n_134), .B1(n_429), .B2(n_430), .Y(n_451) );
AO22x2_ASAP7_75t_L g241 ( .A1(n_101), .A2(n_152), .B1(n_238), .B2(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_102), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_104), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_106), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_107), .A2(n_181), .B1(n_380), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_108), .A2(n_204), .B1(n_391), .B2(n_394), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_109), .A2(n_167), .B1(n_393), .B2(n_432), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_114), .A2(n_206), .B1(n_291), .B2(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g240 ( .A(n_117), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_118), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_120), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_121), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_126), .A2(n_140), .B1(n_333), .B2(n_386), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_127), .A2(n_169), .B1(n_394), .B2(n_476), .Y(n_647) );
INVx1_ASAP7_75t_L g599 ( .A(n_129), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_130), .A2(n_133), .B1(n_400), .B2(n_401), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_131), .B(n_443), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_132), .A2(n_142), .B1(n_610), .B2(n_611), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_135), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_136), .A2(n_147), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_141), .A2(n_184), .B1(n_436), .B2(n_437), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_146), .A2(n_179), .B1(n_393), .B2(n_432), .Y(n_431) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_148), .A2(n_208), .B(n_217), .C(n_635), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_149), .Y(n_262) );
OA22x2_ASAP7_75t_L g375 ( .A1(n_150), .A2(n_376), .B1(n_405), .B2(n_406), .Y(n_375) );
INVx1_ASAP7_75t_L g405 ( .A(n_150), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_153), .A2(n_154), .B1(n_422), .B2(n_423), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_158), .A2(n_176), .B1(n_368), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_161), .A2(n_202), .B1(n_432), .B2(n_453), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_165), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g629 ( .A(n_165), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_166), .Y(n_416) );
INVx1_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
AND2x2_ASAP7_75t_R g657 ( .A(n_172), .B(n_629), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_173), .B(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_174), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_177), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_178), .B(n_336), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_180), .A2(n_203), .B1(n_393), .B2(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g216 ( .A(n_182), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_186), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_190), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_197), .B(n_443), .Y(n_442) );
XOR2x2_ASAP7_75t_L g499 ( .A(n_198), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g659 ( .A1(n_200), .A2(n_640), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_200), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g410 ( .A(n_201), .B(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2x1_ASAP7_75t_R g209 ( .A(n_210), .B(n_212), .Y(n_209) );
OR2x2_ASAP7_75t_L g666 ( .A(n_210), .B(n_213), .Y(n_666) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_211), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_461), .B1(n_624), .B2(n_625), .C(n_626), .Y(n_217) );
INVx1_ASAP7_75t_L g624 ( .A(n_218), .Y(n_624) );
AOI22xp5_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_438), .B1(n_459), .B2(n_460), .Y(n_218) );
INVx1_ASAP7_75t_L g459 ( .A(n_219), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B1(n_408), .B2(n_409), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OAI22xp5_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_223), .B1(n_371), .B2(n_407), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
XNOR2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_323), .Y(n_223) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_322), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_225), .B(n_228), .Y(n_322) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_286), .Y(n_228) );
NOR4xp75_ASAP7_75t_L g229 ( .A(n_230), .B(n_250), .C(n_261), .D(n_275), .Y(n_229) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_SL g330 ( .A(n_233), .Y(n_330) );
INVx4_ASAP7_75t_SL g443 ( .A(n_233), .Y(n_443) );
INVx4_ASAP7_75t_SL g504 ( .A(n_233), .Y(n_504) );
INVx3_ASAP7_75t_L g603 ( .A(n_233), .Y(n_603) );
INVx6_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_243), .Y(n_234) );
AND2x4_ASAP7_75t_L g272 ( .A(n_235), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g284 ( .A(n_235), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g383 ( .A(n_235), .B(n_285), .Y(n_383) );
AND2x4_ASAP7_75t_L g415 ( .A(n_235), .B(n_243), .Y(n_415) );
AND2x2_ASAP7_75t_L g423 ( .A(n_235), .B(n_273), .Y(n_423) );
AND2x2_ASAP7_75t_L g425 ( .A(n_235), .B(n_285), .Y(n_425) );
AND2x2_ASAP7_75t_L g536 ( .A(n_235), .B(n_273), .Y(n_536) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_241), .Y(n_235) );
AND2x2_ASAP7_75t_L g255 ( .A(n_236), .B(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx2_ASAP7_75t_L g281 ( .A(n_236), .Y(n_281) );
OAI22x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_239), .B2(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g242 ( .A(n_238), .Y(n_242) );
INVx2_ASAP7_75t_L g246 ( .A(n_238), .Y(n_246) );
INVx1_ASAP7_75t_L g249 ( .A(n_238), .Y(n_249) );
INVx2_ASAP7_75t_L g256 ( .A(n_241), .Y(n_256) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
AND2x4_ASAP7_75t_L g303 ( .A(n_243), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g312 ( .A(n_243), .B(n_280), .Y(n_312) );
AND2x4_ASAP7_75t_L g319 ( .A(n_243), .B(n_255), .Y(n_319) );
AND2x6_ASAP7_75t_L g393 ( .A(n_243), .B(n_280), .Y(n_393) );
AND2x2_ASAP7_75t_L g400 ( .A(n_243), .B(n_255), .Y(n_400) );
AND2x2_ASAP7_75t_L g436 ( .A(n_243), .B(n_304), .Y(n_436) );
AND2x2_ASAP7_75t_L g571 ( .A(n_243), .B(n_255), .Y(n_571) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g254 ( .A(n_245), .B(n_247), .Y(n_254) );
AND2x2_ASAP7_75t_L g259 ( .A(n_245), .B(n_248), .Y(n_259) );
INVx1_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
INVxp67_ASAP7_75t_L g285 ( .A(n_247), .Y(n_285) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g267 ( .A(n_248), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx3_ASAP7_75t_L g333 ( .A(n_253), .Y(n_333) );
BUFx3_ASAP7_75t_L g385 ( .A(n_253), .Y(n_385) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x4_ASAP7_75t_L g279 ( .A(n_254), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g315 ( .A(n_254), .B(n_304), .Y(n_315) );
AND2x2_ASAP7_75t_L g382 ( .A(n_254), .B(n_280), .Y(n_382) );
AND2x4_ASAP7_75t_L g418 ( .A(n_254), .B(n_255), .Y(n_418) );
AND2x2_ASAP7_75t_L g437 ( .A(n_254), .B(n_304), .Y(n_437) );
AND2x2_ASAP7_75t_L g534 ( .A(n_254), .B(n_280), .Y(n_534) );
AND2x2_ASAP7_75t_L g266 ( .A(n_255), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g422 ( .A(n_255), .B(n_267), .Y(n_422) );
AND2x4_ASAP7_75t_L g304 ( .A(n_256), .B(n_281), .Y(n_304) );
INVx2_ASAP7_75t_L g337 ( .A(n_257), .Y(n_337) );
BUFx3_ASAP7_75t_L g620 ( .A(n_257), .Y(n_620) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g387 ( .A(n_258), .Y(n_387) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x4_ASAP7_75t_L g296 ( .A(n_259), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g321 ( .A(n_259), .B(n_304), .Y(n_321) );
AND2x4_ASAP7_75t_L g401 ( .A(n_259), .B(n_304), .Y(n_401) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_259), .B(n_260), .Y(n_419) );
AND2x4_ASAP7_75t_L g430 ( .A(n_259), .B(n_297), .Y(n_430) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_259), .B(n_260), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B1(n_269), .B2(n_270), .Y(n_261) );
INVx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g486 ( .A(n_265), .Y(n_486) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_266), .Y(n_379) );
AND2x2_ASAP7_75t_L g293 ( .A(n_267), .B(n_280), .Y(n_293) );
AND2x4_ASAP7_75t_L g307 ( .A(n_267), .B(n_304), .Y(n_307) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_267), .B(n_280), .Y(n_429) );
AND2x6_ASAP7_75t_L g432 ( .A(n_267), .B(n_304), .Y(n_432) );
AND2x2_ASAP7_75t_L g591 ( .A(n_267), .B(n_280), .Y(n_591) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_268), .Y(n_274) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g366 ( .A(n_272), .Y(n_366) );
BUFx6f_ASAP7_75t_SL g380 ( .A(n_272), .Y(n_380) );
BUFx3_ASAP7_75t_L g606 ( .A(n_272), .Y(n_606) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B1(n_282), .B2(n_283), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g368 ( .A(n_278), .Y(n_368) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
BUFx3_ASAP7_75t_L g483 ( .A(n_279), .Y(n_483) );
BUFx2_ASAP7_75t_L g510 ( .A(n_279), .Y(n_510) );
INVx2_ASAP7_75t_L g369 ( .A(n_283), .Y(n_369) );
INVx2_ASAP7_75t_SL g484 ( .A(n_283), .Y(n_484) );
INVx2_ASAP7_75t_L g511 ( .A(n_283), .Y(n_511) );
INVx2_ASAP7_75t_L g618 ( .A(n_283), .Y(n_618) );
INVx6_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_308), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_298), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g610 ( .A(n_290), .Y(n_610) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g397 ( .A(n_292), .Y(n_397) );
INVx1_ASAP7_75t_L g515 ( .A(n_292), .Y(n_515) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_293), .Y(n_343) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_340), .B1(n_341), .B2(n_344), .Y(n_339) );
INVx2_ASAP7_75t_L g643 ( .A(n_295), .Y(n_643) );
INVx5_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g398 ( .A(n_296), .Y(n_398) );
BUFx2_ASAP7_75t_L g479 ( .A(n_296), .Y(n_479) );
BUFx3_ASAP7_75t_L g611 ( .A(n_296), .Y(n_611) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_SL g360 ( .A(n_302), .Y(n_360) );
INVx3_ASAP7_75t_SL g403 ( .A(n_302), .Y(n_403) );
INVx3_ASAP7_75t_L g453 ( .A(n_302), .Y(n_453) );
INVx2_ASAP7_75t_SL g489 ( .A(n_302), .Y(n_489) );
INVx2_ASAP7_75t_L g615 ( .A(n_302), .Y(n_615) );
INVx8_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_306), .A2(n_346), .B1(n_347), .B2(n_350), .Y(n_345) );
INVx2_ASAP7_75t_SL g404 ( .A(n_306), .Y(n_404) );
INVx2_ASAP7_75t_L g494 ( .A(n_306), .Y(n_494) );
INVx2_ASAP7_75t_L g614 ( .A(n_306), .Y(n_614) );
INVx8_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_316), .Y(n_308) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
INVx2_ASAP7_75t_L g517 ( .A(n_311), .Y(n_517) );
INVx3_ASAP7_75t_L g645 ( .A(n_311), .Y(n_645) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g493 ( .A(n_312), .Y(n_493) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g362 ( .A(n_314), .Y(n_362) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g395 ( .A(n_315), .Y(n_395) );
BUFx3_ASAP7_75t_L g477 ( .A(n_315), .Y(n_477) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_315), .Y(n_521) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_318), .A2(n_353), .B1(n_354), .B2(n_355), .Y(n_352) );
INVx2_ASAP7_75t_L g608 ( .A(n_318), .Y(n_608) );
INVx6_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx3_ASAP7_75t_L g476 ( .A(n_319), .Y(n_476) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
BUFx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g491 ( .A(n_321), .Y(n_491) );
XNOR2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_370), .Y(n_323) );
NAND4xp75_ASAP7_75t_L g324 ( .A(n_325), .B(n_338), .C(n_351), .D(n_363), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_331), .B2(n_334), .C(n_335), .Y(n_326) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g471 ( .A(n_330), .Y(n_471) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_L g338 ( .A(n_339), .B(n_345), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2x1_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_361), .B2(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx2_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_366), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_556) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_389), .Y(n_376) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .C(n_384), .D(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g558 ( .A(n_379), .Y(n_558) );
BUFx6f_ASAP7_75t_SL g617 ( .A(n_379), .Y(n_617) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_390), .B(n_396), .C(n_399), .D(n_402), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_394), .Y(n_622) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g457 ( .A(n_395), .Y(n_457) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_426), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_420), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_416), .B(n_417), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g555 ( .A(n_415), .Y(n_555) );
INVx1_ASAP7_75t_SL g654 ( .A(n_418), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVxp67_ASAP7_75t_L g564 ( .A(n_425), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_433), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g460 ( .A(n_438), .Y(n_460) );
XOR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_458), .Y(n_438) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_449), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_446), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g625 ( .A(n_461), .Y(n_625) );
XOR2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_579), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_524), .B1(n_576), .B2(n_578), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g577 ( .A(n_464), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_497), .B(n_522), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_465), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g495 ( .A(n_468), .Y(n_495) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_480), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
OAI21xp33_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_472), .B(n_473), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_478), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_487), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .Y(n_487) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g523 ( .A(n_498), .Y(n_523) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
OAI21xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_505), .B(n_506), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_545), .B2(n_574), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_544), .Y(n_528) );
NAND2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_537), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVxp67_ASAP7_75t_L g562 ( .A(n_534), .Y(n_562) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g575 ( .A(n_548), .Y(n_575) );
INVx1_ASAP7_75t_L g573 ( .A(n_550), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_565), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .C(n_560), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_596), .B2(n_623), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
XNOR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_595), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .C(n_587), .D(n_588), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .C(n_593), .D(n_594), .Y(n_589) );
INVx1_ASAP7_75t_L g623 ( .A(n_596), .Y(n_623) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
XNOR2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_612), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .C(n_607), .D(n_609), .Y(n_601) );
BUFx6f_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .C(n_619), .D(n_621), .Y(n_612) );
INVx3_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_628), .B(n_631), .Y(n_665) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OAI222xp33_ASAP7_75t_R g635 ( .A1(n_636), .A2(n_656), .B1(n_658), .B2(n_662), .C1(n_663), .C2(n_666), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2x1_ASAP7_75t_SL g660 ( .A(n_640), .B(n_661), .Y(n_660) );
NAND4xp75_ASAP7_75t_L g640 ( .A(n_641), .B(n_646), .C(n_649), .D(n_652), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
CKINVDCx6p67_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
endmodule