module real_jpeg_23833_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_288;
wire n_292;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_295;
wire n_202;
wire n_133;
wire n_167;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_4),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_131),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_131),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_8),
.A2(n_29),
.B1(n_31),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_34),
.B1(n_51),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_20),
.B1(n_62),
.B2(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_20),
.B1(n_29),
.B2(n_31),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_27),
.B(n_186),
.C(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_28),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_10),
.A2(n_31),
.B(n_43),
.C(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_10),
.B(n_60),
.C(n_62),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_10),
.B(n_71),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_10),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_10),
.B(n_61),
.Y(n_256)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_11),
.B(n_239),
.Y(n_244)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_93),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.C(n_78),
.Y(n_15)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_16),
.B(n_69),
.CI(n_78),
.CON(n_300),
.SN(n_300)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_37),
.B1(n_67),
.B2(n_68),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_17),
.A2(n_67),
.B1(n_95),
.B2(n_108),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_39),
.C(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_32),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_18),
.B(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_19),
.B(n_28),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_20),
.A2(n_26),
.B(n_31),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_20),
.A2(n_45),
.B(n_47),
.Y(n_210)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_23),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_23),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_28),
.A2(n_103),
.B(n_106),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_28),
.B(n_130),
.Y(n_151)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_31),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_32),
.B(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_50),
.B(n_52),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_40),
.B(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_53),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_41),
.A2(n_46),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_41),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_46),
.B(n_100),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_48),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_52),
.B(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_55),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_54),
.B(n_168),
.C(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_54),
.A2(n_55),
.B1(n_170),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_65),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_57),
.B(n_66),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_57),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_61),
.B(n_214),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_62),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_64),
.A2(n_76),
.B(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_69),
.A2(n_70),
.B(n_73),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_71),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_72),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_74),
.B(n_212),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_76),
.B(n_224),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B(n_88),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_85),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_79),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_79),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_79),
.A2(n_138),
.B1(n_209),
.B2(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_80),
.B(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_80),
.B(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_87),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_87),
.B(n_213),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_99),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_297),
.B(n_301),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_160),
.B(n_296),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_152),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_115),
.B(n_152),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_136),
.C(n_139),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_116),
.B(n_136),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_126),
.C(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_118),
.B(n_124),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_119),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_143),
.B(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_122),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_135),
.B(n_172),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_139),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_150),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_140),
.A2(n_141),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_145),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_145),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_148),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_149),
.A2(n_150),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_149),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_299)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_291),
.B(n_295),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_202),
.B(n_277),
.C(n_290),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_190),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_163),
.B(n_190),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_176),
.B2(n_189),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_174),
.B2(n_175),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_166),
.B(n_175),
.C(n_189),
.Y(n_278)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_169),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_178),
.B(n_183),
.C(n_184),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_192),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_276),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_218),
.B(n_275),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_205),
.B(n_215),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_211),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_270),
.B(n_274),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_261),
.B(n_269),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_241),
.B(n_260),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_240),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_234),
.C(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_235),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_247),
.B(n_259),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_245),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_258),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_287),
.B2(n_288),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_288),
.C(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_300),
.Y(n_303)
);


endmodule