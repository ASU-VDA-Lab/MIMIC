module fake_jpeg_11912_n_388 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_45),
.B(n_51),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_50),
.Y(n_97)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_25),
.B(n_0),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_61),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_62),
.B(n_70),
.Y(n_126)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_63),
.Y(n_107)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_9),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_73),
.Y(n_102)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_43),
.B1(n_19),
.B2(n_24),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_79),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_1),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_33),
.B1(n_21),
.B2(n_36),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_84),
.A2(n_103),
.B1(n_56),
.B2(n_61),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_21),
.B1(n_33),
.B2(n_17),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_101),
.B1(n_113),
.B2(n_122),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_21),
.B1(n_33),
.B2(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_89),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_91),
.B(n_4),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_28),
.B1(n_20),
.B2(n_36),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_115),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_28),
.B1(n_36),
.B2(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_28),
.B1(n_54),
.B2(n_80),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_35),
.B1(n_42),
.B2(n_18),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_42),
.B1(n_43),
.B2(n_35),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_60),
.B1(n_78),
.B2(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_41),
.B1(n_22),
.B2(n_17),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_41),
.B1(n_22),
.B2(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_124),
.B1(n_125),
.B2(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_119),
.B(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_51),
.B(n_10),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_66),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OR2x2_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_45),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g205 ( 
.A(n_130),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

OR2x4_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_45),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_57),
.C(n_16),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_164),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_89),
.A2(n_76),
.B1(n_46),
.B2(n_50),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_75),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_147),
.C(n_159),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_69),
.B1(n_64),
.B2(n_65),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_149),
.B(n_150),
.Y(n_201)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_163),
.B1(n_106),
.B2(n_108),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_1),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_63),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_151),
.B(n_160),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_105),
.A2(n_61),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_120),
.B1(n_106),
.B2(n_95),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_90),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_82),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_161),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_6),
.B(n_7),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_99),
.A2(n_7),
.B(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_13),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_169),
.Y(n_206)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_116),
.Y(n_182)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_14),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_104),
.B(n_16),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_129),
.B(n_98),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_118),
.B1(n_111),
.B2(n_85),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_191),
.B1(n_203),
.B2(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_98),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_114),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_168),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_118),
.B1(n_85),
.B2(n_111),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_81),
.Y(n_188)
);

CKINVDCx11_ASAP7_75t_R g197 ( 
.A(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_156),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_147),
.B(n_109),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_211),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_141),
.B(n_123),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_207),
.C(n_165),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_100),
.B1(n_108),
.B2(n_123),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_81),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_131),
.A2(n_100),
.B1(n_88),
.B2(n_116),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_210),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_140),
.B(n_88),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_147),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_140),
.B1(n_131),
.B2(n_148),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_212),
.A2(n_229),
.B1(n_240),
.B2(n_185),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_205),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_223),
.Y(n_257)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_230),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_160),
.B(n_148),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_136),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_233),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_207),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_134),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_238),
.C(n_199),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_184),
.A2(n_128),
.B1(n_139),
.B2(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_153),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_174),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_244),
.B(n_239),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_152),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_161),
.A3(n_155),
.B1(n_158),
.B2(n_162),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_144),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_146),
.B1(n_167),
.B2(n_178),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_172),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_202),
.B(n_185),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_197),
.B(n_182),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_172),
.B(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_185),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_254),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_198),
.B(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_262),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_261),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_234),
.C(n_225),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_230),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_227),
.A2(n_208),
.B1(n_186),
.B2(n_181),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_224),
.B1(n_275),
.B2(n_270),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_180),
.B(n_190),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_187),
.C(n_185),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_274),
.B1(n_277),
.B2(n_241),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_187),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_214),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_271),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_212),
.A2(n_194),
.B1(n_206),
.B2(n_187),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_227),
.A2(n_194),
.B1(n_192),
.B2(n_204),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_246),
.B1(n_229),
.B2(n_213),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_297),
.B1(n_299),
.B2(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_282),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_213),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_294),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_252),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_269),
.B1(n_253),
.B2(n_254),
.Y(n_307)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_302),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_270),
.B1(n_259),
.B2(n_275),
.Y(n_299)
);

BUFx12f_ASAP7_75t_SL g300 ( 
.A(n_264),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.C(n_258),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_242),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_320),
.B1(n_289),
.B2(n_288),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_261),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_309),
.C(n_317),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_247),
.B1(n_274),
.B2(n_251),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_249),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_246),
.B1(n_217),
.B2(n_221),
.Y(n_312)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_248),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_280),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_256),
.B(n_262),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_314),
.A2(n_302),
.B(n_218),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_248),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_217),
.B1(n_273),
.B2(n_223),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_285),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_237),
.B(n_252),
.C(n_190),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_319),
.A2(n_272),
.B(n_278),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_287),
.A2(n_265),
.B1(n_245),
.B2(n_272),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_230),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_279),
.C(n_291),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_283),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_326),
.B(n_334),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_330),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_331),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_306),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_286),
.C(n_296),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_335),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_319),
.B(n_303),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_177),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_268),
.C(n_281),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_336),
.A2(n_321),
.B1(n_315),
.B2(n_303),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_337),
.A2(n_314),
.B(n_319),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_268),
.C(n_298),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_340),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_260),
.C(n_216),
.Y(n_340)
);

AO22x1_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_347),
.B1(n_319),
.B2(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_349),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_320),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_354),
.B(n_325),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_321),
.B(n_311),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_336),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_340),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_260),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_L g355 ( 
.A1(n_346),
.A2(n_339),
.B(n_330),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_359),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_338),
.C(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_356),
.B(n_361),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_358),
.B(n_192),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_190),
.B(n_204),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_328),
.C(n_322),
.Y(n_361)
);

OAI221xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_313),
.B1(n_236),
.B2(n_215),
.C(n_231),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_362),
.B(n_364),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_363),
.A2(n_349),
.B1(n_347),
.B2(n_343),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_232),
.C(n_290),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_367),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_358),
.A2(n_352),
.B1(n_219),
.B2(n_353),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_357),
.A2(n_228),
.B1(n_290),
.B2(n_180),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_363),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_361),
.B(n_228),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_364),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_173),
.C(n_193),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_373),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_366),
.Y(n_374)
);

AOI322xp5_ASAP7_75t_L g383 ( 
.A1(n_374),
.A2(n_355),
.A3(n_368),
.B1(n_376),
.B2(n_366),
.C1(n_378),
.C2(n_365),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_375),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_377),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_379),
.A2(n_370),
.B(n_367),
.Y(n_381)
);

AOI21x1_ASAP7_75t_L g385 ( 
.A1(n_381),
.A2(n_383),
.B(n_173),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_376),
.C(n_173),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_384),
.A2(n_385),
.B(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_193),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_193),
.Y(n_388)
);


endmodule