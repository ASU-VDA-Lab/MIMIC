module real_jpeg_12379_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_249, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_249;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_65;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_5),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_67),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_6),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_8),
.A2(n_62),
.B1(n_68),
.B2(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_62),
.Y(n_150)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_71),
.B(n_74),
.C(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_10),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_68),
.B1(n_71),
.B2(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_10),
.B(n_79),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_10),
.A2(n_24),
.B1(n_35),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_10),
.B(n_107),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_68),
.B1(n_71),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_11),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_112),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_112),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_14),
.A2(n_68),
.B1(n_71),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_78),
.Y(n_213)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_140),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_20),
.B(n_114),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_92),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_21),
.B(n_80),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_52),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_22),
.B(n_53),
.C(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_23),
.B(n_38),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_24),
.A2(n_35),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_24),
.A2(n_35),
.B1(n_211),
.B2(n_219),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_24),
.A2(n_83),
.B(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_25),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_25),
.A2(n_34),
.B(n_84),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_25),
.A2(n_29),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_26),
.B(n_40),
.C(n_101),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_217),
.Y(n_216)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_35),
.A2(n_85),
.B(n_98),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_35),
.B(n_101),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_47),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_39),
.B(n_49),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_39),
.B(n_101),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_51)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

OA22x2_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_43),
.A2(n_56),
.B(n_180),
.C(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_43),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_44),
.B(n_57),
.C(n_59),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_90),
.B(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_50),
.A2(n_122),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_50),
.A2(n_89),
.B1(n_187),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_50),
.A2(n_89),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_50),
.A2(n_89),
.B1(n_196),
.B2(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_61),
.B(n_63),
.Y(n_53)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_54),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_54),
.A2(n_104),
.B1(n_107),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_54),
.A2(n_107),
.B1(n_168),
.B2(n_181),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_55),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_55),
.A2(n_105),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_75),
.B(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_60),
.B(n_101),
.CON(n_181),
.SN(n_181)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_72),
.B1(n_77),
.B2(n_79),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_72),
.A2(n_79),
.B1(n_111),
.B2(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_77),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_91),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_91),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_108),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_94),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B(n_106),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_138),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_123),
.B1(n_136),
.B2(n_137),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

AOI221xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_156),
.B1(n_172),
.B2(n_247),
.C(n_249),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_142),
.B(n_144),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_155),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_151),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_157),
.B(n_170),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_158),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_162),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.C(n_166),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_246),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_241),
.B(n_245),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_197),
.B(n_240),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_192),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_178),
.B(n_184),
.C(n_189),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B(n_188),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_195),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_235),
.B(n_239),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_225),
.B(n_234),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_214),
.B(n_224),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_207),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_220),
.B(n_223),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_230),
.C(n_233),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_238),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_244),
.Y(n_245)
);


endmodule