module fake_aes_6967_n_692 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_692);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_692;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g77 ( .A(n_33), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_22), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_17), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_74), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_76), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_57), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
CKINVDCx14_ASAP7_75t_R g85 ( .A(n_49), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_43), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_14), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_63), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_65), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_13), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_56), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_48), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_64), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_47), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_26), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_34), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_62), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_17), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_31), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_54), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_6), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_3), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_24), .Y(n_109) );
INVxp33_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_28), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_30), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_60), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_5), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_75), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_40), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_39), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_23), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_19), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_1), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_124), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_100), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_100), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_118), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_80), .A2(n_32), .B(n_70), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
INVx5_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_121), .B(n_0), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_121), .B(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
NOR2xp67_ASAP7_75t_L g144 ( .A(n_79), .B(n_1), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_79), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_118), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
NOR2xp33_ASAP7_75t_R g148 ( .A(n_85), .B(n_35), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_95), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_107), .B(n_2), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_106), .Y(n_153) );
NOR2xp33_ASAP7_75t_R g154 ( .A(n_120), .B(n_29), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_101), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_117), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_89), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_89), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_87), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_91), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_87), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_130), .B(n_84), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_139), .B(n_88), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_155), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_139), .B(n_97), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_130), .B(n_96), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_139), .B(n_94), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_139), .B(n_112), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_139), .B(n_116), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_145), .B(n_122), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx8_ASAP7_75t_L g188 ( .A(n_139), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_157), .A2(n_114), .B1(n_107), .B2(n_108), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_125), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_126), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_134), .A2(n_122), .B1(n_108), .B2(n_115), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_166), .B(n_119), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_125), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_166), .B(n_119), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_146), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_129), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_125), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_125), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_126), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
NAND3xp33_ASAP7_75t_L g203 ( .A(n_164), .B(n_115), .C(n_113), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_128), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx4_ASAP7_75t_SL g207 ( .A(n_158), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_167), .B(n_113), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_127), .Y(n_212) );
AND3x4_ASAP7_75t_L g213 ( .A(n_144), .B(n_2), .C(n_4), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_128), .B(n_111), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_131), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_136), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_131), .B(n_111), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_137), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_160), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_137), .B(n_109), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_165), .B(n_163), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_165), .B(n_163), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_162), .B(n_109), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_140), .B(n_105), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
BUFx4f_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_173), .B(n_133), .Y(n_230) );
AND3x1_ASAP7_75t_SL g231 ( .A(n_213), .B(n_197), .C(n_104), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_223), .B(n_162), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_159), .B1(n_143), .B2(n_147), .Y(n_235) );
BUFx4f_ASAP7_75t_SL g236 ( .A(n_184), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_211), .A2(n_159), .B1(n_143), .B2(n_147), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_208), .Y(n_238) );
AOI22xp5_ASAP7_75t_SL g239 ( .A1(n_197), .A2(n_149), .B1(n_153), .B2(n_98), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g240 ( .A(n_169), .B(n_132), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_177), .B(n_171), .Y(n_241) );
NOR2xp33_ASAP7_75t_R g242 ( .A(n_184), .B(n_141), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_223), .B(n_142), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_188), .Y(n_244) );
NOR3xp33_ASAP7_75t_SL g245 ( .A(n_203), .B(n_92), .C(n_98), .Y(n_245) );
NOR2xp33_ASAP7_75t_R g246 ( .A(n_183), .B(n_138), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_223), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_211), .B(n_150), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_183), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
BUFx12f_ASAP7_75t_L g251 ( .A(n_171), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_224), .B(n_154), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_210), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_224), .B(n_138), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_225), .B(n_138), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_187), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_225), .B(n_138), .Y(n_261) );
INVx5_ASAP7_75t_L g262 ( .A(n_188), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_188), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_217), .B(n_150), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
NOR3xp33_ASAP7_75t_SL g266 ( .A(n_222), .B(n_99), .C(n_103), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
NAND2xp33_ASAP7_75t_R g268 ( .A(n_185), .B(n_148), .Y(n_268) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_225), .B(n_105), .Y(n_269) );
INVx5_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_185), .B(n_150), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_218), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_170), .A2(n_161), .B1(n_160), .B2(n_132), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_192), .B(n_83), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_228), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_196), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_220), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_217), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_200), .B(n_150), .Y(n_282) );
INVx4_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_204), .B(n_104), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_215), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_213), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_212), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_219), .B(n_103), .Y(n_288) );
BUFx10_ASAP7_75t_L g289 ( .A(n_178), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_179), .B(n_99), .Y(n_290) );
INVx5_ASAP7_75t_L g291 ( .A(n_175), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_193), .Y(n_292) );
NOR3xp33_ASAP7_75t_SL g293 ( .A(n_227), .B(n_4), .C(n_5), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_241), .B(n_189), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_249), .B(n_195), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_262), .B(n_209), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_247), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_269), .A2(n_209), .B1(n_214), .B2(n_206), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_235), .A2(n_182), .B1(n_181), .B2(n_172), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
CKINVDCx6p67_ASAP7_75t_R g304 ( .A(n_251), .Y(n_304) );
AOI22xp5_ASAP7_75t_SL g305 ( .A1(n_286), .A2(n_209), .B1(n_180), .B2(n_174), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_266), .A2(n_199), .B(n_168), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_262), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_236), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_267), .A2(n_216), .B(n_206), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_276), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_281), .B(n_160), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
AND2x6_ASAP7_75t_L g313 ( .A(n_244), .B(n_216), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_250), .B(n_226), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_292), .B(n_206), .Y(n_315) );
NOR2x1_ASAP7_75t_L g316 ( .A(n_250), .B(n_221), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_230), .A2(n_216), .B1(n_206), .B2(n_205), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_269), .A2(n_216), .B1(n_205), .B2(n_206), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_251), .B(n_226), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_262), .Y(n_321) );
BUFx12f_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_244), .B(n_216), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_277), .B(n_226), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_283), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_235), .B(n_161), .Y(n_330) );
INVx4_ASAP7_75t_SL g331 ( .A(n_263), .Y(n_331) );
INVx3_ASAP7_75t_SL g332 ( .A(n_239), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_287), .B(n_7), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_248), .B(n_205), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_289), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_289), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_271), .A2(n_160), .B1(n_161), .B2(n_205), .C(n_221), .Y(n_337) );
INVx6_ASAP7_75t_L g338 ( .A(n_283), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_289), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_264), .B(n_161), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_229), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_229), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_229), .B(n_221), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_301), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_309), .A2(n_275), .B(n_285), .Y(n_346) );
NAND3xp33_ASAP7_75t_SL g347 ( .A(n_326), .B(n_242), .C(n_293), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_294), .A2(n_237), .B(n_274), .C(n_252), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
BUFx4f_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_295), .B(n_264), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_333), .A2(n_264), .B1(n_248), .B2(n_257), .C(n_290), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g353 ( .A(n_308), .B(n_245), .C(n_259), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_322), .A2(n_290), .B1(n_257), .B2(n_243), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_290), .B1(n_267), .B2(n_285), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_315), .A2(n_275), .A3(n_288), .B(n_284), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_298), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_304), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_310), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_260), .B1(n_258), .B2(n_232), .Y(n_361) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_321), .B(n_283), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_303), .A2(n_240), .B(n_258), .C(n_260), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_330), .A2(n_231), .B1(n_268), .B2(n_240), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_301), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_333), .A2(n_261), .B1(n_265), .B2(n_280), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_310), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_295), .A2(n_280), .B1(n_265), .B2(n_278), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_308), .A2(n_282), .B1(n_276), .B2(n_161), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_304), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_335), .B(n_272), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_314), .A2(n_332), .B1(n_316), .B2(n_330), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_332), .A2(n_278), .B1(n_272), .B2(n_220), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_335), .B(n_272), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_347), .A2(n_306), .B1(n_340), .B2(n_311), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_352), .A2(n_306), .B1(n_340), .B2(n_300), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_366), .A2(n_339), .B1(n_336), .B2(n_321), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_351), .B(n_327), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_364), .A2(n_317), .B(n_296), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_368), .A2(n_318), .B1(n_334), .B2(n_336), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g383 ( .A1(n_349), .A2(n_305), .B1(n_313), .B2(n_339), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_348), .A2(n_320), .B(n_337), .C(n_296), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_334), .B1(n_329), .B2(n_338), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_346), .A2(n_334), .B(n_312), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_306), .B1(n_302), .B2(n_328), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_334), .B(n_344), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_329), .B1(n_338), .B2(n_325), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_360), .A2(n_344), .B(n_312), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_374), .A2(n_338), .B1(n_325), .B2(n_341), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_354), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_321), .B1(n_324), .B2(n_341), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_351), .A2(n_328), .B1(n_324), .B2(n_325), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_365), .B(n_328), .Y(n_396) );
OR2x6_ASAP7_75t_L g397 ( .A(n_345), .B(n_367), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_360), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_355), .A2(n_324), .B1(n_342), .B2(n_307), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_360), .A2(n_168), .B(n_194), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_369), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_301), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_345), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_398), .B(n_357), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_391), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_398), .B(n_357), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_403), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_397), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_380), .B(n_359), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_401), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_402), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_401), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_380), .A2(n_365), .B1(n_358), .B2(n_363), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_403), .Y(n_417) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_386), .A2(n_369), .B(n_363), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g419 ( .A1(n_393), .A2(n_350), .B(n_362), .C(n_370), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_393), .B(n_357), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_383), .A2(n_371), .B1(n_350), .B2(n_345), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_378), .A2(n_372), .B1(n_375), .B2(n_161), .C(n_373), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_369), .B(n_367), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_381), .A2(n_194), .B(n_199), .Y(n_428) );
NOR2x1_ASAP7_75t_SL g429 ( .A(n_397), .B(n_345), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_385), .A2(n_350), .B1(n_362), .B2(n_307), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_404), .B(n_357), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_396), .B(n_357), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_396), .A2(n_373), .B1(n_313), .B2(n_376), .Y(n_433) );
AOI21xp5_ASAP7_75t_SL g434 ( .A1(n_385), .A2(n_342), .B(n_307), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_379), .A2(n_373), .B(n_357), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_404), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_377), .B(n_373), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_382), .A2(n_313), .B1(n_307), .B2(n_276), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_382), .A2(n_343), .B(n_238), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_411), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_431), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_431), .B(n_404), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_409), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_410), .B(n_387), .C(n_384), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_409), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_410), .B(n_397), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
AOI33xp33_ASAP7_75t_L g450 ( .A1(n_416), .A2(n_395), .A3(n_394), .B1(n_273), .B2(n_10), .B3(n_11), .Y(n_450) );
AOI221xp5_ASAP7_75t_SL g451 ( .A1(n_412), .A2(n_392), .B1(n_399), .B2(n_389), .C(n_175), .Y(n_451) );
HB1xp67_ASAP7_75t_SL g452 ( .A(n_421), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_432), .B(n_389), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_431), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_405), .B(n_407), .Y(n_457) );
INVxp67_ASAP7_75t_SL g458 ( .A(n_405), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_416), .A2(n_392), .B1(n_399), .B2(n_175), .C(n_190), .Y(n_460) );
OAI31xp33_ASAP7_75t_L g461 ( .A1(n_421), .A2(n_343), .A3(n_202), .B(n_279), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g462 ( .A(n_425), .B(n_400), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_420), .B(n_400), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_432), .B(n_7), .Y(n_466) );
NOR2xp33_ASAP7_75t_R g467 ( .A(n_412), .B(n_8), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_420), .B(n_8), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_408), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
NAND3xp33_ASAP7_75t_SL g471 ( .A(n_426), .B(n_9), .C(n_10), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_405), .B(n_11), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_426), .A2(n_313), .B1(n_331), .B2(n_175), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_407), .B(n_12), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_407), .B(n_12), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_430), .A2(n_190), .B1(n_198), .B2(n_233), .C(n_234), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_408), .B(n_13), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_425), .B(n_14), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_413), .B(n_15), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_418), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_425), .B(n_15), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_424), .B(n_16), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_424), .B(n_16), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_430), .A2(n_313), .B1(n_331), .B2(n_279), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_436), .B(n_18), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_457), .B(n_439), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_458), .B(n_435), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_469), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_457), .B(n_439), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_442), .B(n_439), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_464), .B(n_435), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_440), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_442), .B(n_439), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_476), .B(n_429), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_476), .B(n_429), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_442), .B(n_439), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_464), .B(n_456), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_448), .B(n_18), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_443), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_455), .B(n_435), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_445), .B(n_19), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_455), .B(n_435), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_467), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_480), .Y(n_512) );
INVxp33_ASAP7_75t_SL g513 ( .A(n_477), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_449), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_454), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_470), .B(n_473), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_444), .B(n_435), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_477), .B(n_437), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_463), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_444), .B(n_418), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_480), .Y(n_522) );
NAND5xp2_ASAP7_75t_L g523 ( .A(n_451), .B(n_438), .C(n_419), .D(n_433), .E(n_437), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_449), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_466), .B(n_418), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_466), .B(n_418), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_453), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_468), .B(n_418), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_453), .B(n_418), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_454), .B(n_427), .Y(n_532) );
OAI33xp33_ASAP7_75t_L g533 ( .A1(n_481), .A2(n_20), .A3(n_423), .B1(n_422), .B2(n_419), .B3(n_434), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_446), .B(n_438), .C(n_433), .D(n_423), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_483), .Y(n_535) );
AOI32xp33_ASAP7_75t_L g536 ( .A1(n_484), .A2(n_20), .A3(n_423), .B1(n_422), .B2(n_427), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_441), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_482), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_465), .B(n_427), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_481), .A2(n_423), .B1(n_427), .B2(n_422), .C(n_414), .Y(n_541) );
OAI31xp33_ASAP7_75t_L g542 ( .A1(n_484), .A2(n_422), .A3(n_331), .B(n_427), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_445), .B(n_21), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_478), .B(n_414), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_474), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_472), .B(n_414), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
A2O1A1O1Ixp25_ASAP7_75t_L g549 ( .A1(n_505), .A2(n_452), .B(n_486), .C(n_485), .D(n_489), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_511), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_533), .B(n_471), .C(n_450), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_447), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_491), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_512), .B(n_447), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_522), .B(n_474), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_504), .B(n_513), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_531), .B(n_474), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_509), .A2(n_461), .B(n_475), .C(n_460), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_493), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_513), .B(n_414), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_511), .A2(n_462), .B(n_488), .C(n_479), .Y(n_566) );
INVx4_ASAP7_75t_L g567 ( .A(n_516), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_531), .B(n_414), .Y(n_568) );
INVx3_ASAP7_75t_SL g569 ( .A(n_538), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_506), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_514), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_500), .B(n_414), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_535), .B(n_414), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_541), .A2(n_462), .B(n_428), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_517), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_514), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_532), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_501), .B(n_414), .Y(n_578) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_532), .A2(n_331), .A3(n_41), .B1(n_42), .B2(n_44), .Y(n_579) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_536), .A2(n_428), .B(n_45), .Y(n_580) );
AOI21xp33_ASAP7_75t_SL g581 ( .A1(n_542), .A2(n_428), .B(n_46), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_524), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_518), .A2(n_190), .B(n_198), .Y(n_583) );
NOR4xp25_ASAP7_75t_L g584 ( .A(n_534), .B(n_428), .C(n_50), .D(n_51), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_518), .B(n_428), .Y(n_585) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_492), .A2(n_428), .B(n_53), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_524), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_507), .A2(n_198), .B(n_190), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_540), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_535), .B(n_198), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_521), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_528), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_519), .A2(n_313), .B1(n_207), .B2(n_291), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_521), .B(n_36), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_544), .A2(n_207), .B1(n_291), .B2(n_270), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_530), .B(n_55), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_256), .B(n_255), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_530), .B(n_59), .Y(n_599) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_567), .A2(n_507), .B1(n_510), .B2(n_492), .C1(n_497), .C2(n_526), .Y(n_600) );
AOI211xp5_ASAP7_75t_SL g601 ( .A1(n_580), .A2(n_510), .B(n_497), .C(n_529), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_592), .B(n_539), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_589), .B(n_575), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_551), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_590), .B(n_490), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_563), .B(n_494), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_577), .B(n_494), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_569), .B(n_523), .Y(n_610) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_567), .A2(n_539), .B(n_546), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_560), .B(n_543), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_556), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_559), .B(n_546), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_561), .B(n_543), .Y(n_615) );
O2A1O1Ixp33_ASAP7_75t_SL g616 ( .A1(n_566), .A2(n_528), .B(n_498), .C(n_547), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_561), .B(n_496), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_570), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_585), .B(n_496), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_550), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_576), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_554), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_582), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_587), .B(n_499), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_593), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_557), .B(n_499), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_579), .A2(n_502), .B(n_545), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_545), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_568), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_568), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_572), .B(n_502), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_573), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_552), .B(n_527), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_635), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_615), .Y(n_638) );
O2A1O1Ixp5_ASAP7_75t_L g639 ( .A1(n_610), .A2(n_574), .B(n_595), .C(n_580), .Y(n_639) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_610), .A2(n_553), .B(n_574), .C(n_562), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_611), .A2(n_581), .B(n_584), .C(n_595), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_630), .A2(n_578), .B(n_573), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_623), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_625), .A2(n_599), .B1(n_597), .B2(n_586), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_603), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_616), .B(n_599), .C(n_597), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_605), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_635), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_614), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_636), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_616), .B(n_591), .C(n_598), .Y(n_651) );
XOR2x2_ASAP7_75t_L g652 ( .A(n_604), .B(n_549), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_632), .B(n_495), .Y(n_653) );
OA22x2_ASAP7_75t_L g654 ( .A1(n_608), .A2(n_583), .B1(n_588), .B2(n_598), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_633), .Y(n_655) );
NOR2xp33_ASAP7_75t_SL g656 ( .A(n_600), .B(n_527), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_612), .B(n_591), .Y(n_657) );
OAI31xp33_ASAP7_75t_L g658 ( .A1(n_601), .A2(n_520), .A3(n_515), .B(n_508), .Y(n_658) );
AO22x2_ASAP7_75t_L g659 ( .A1(n_643), .A2(n_621), .B1(n_606), .B2(n_613), .Y(n_659) );
NAND4xp75_ASAP7_75t_L g660 ( .A(n_639), .B(n_636), .C(n_629), .D(n_607), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_640), .B(n_596), .C(n_609), .D(n_617), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_642), .A2(n_626), .B1(n_618), .B2(n_628), .C(n_619), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_645), .Y(n_663) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_656), .A2(n_614), .B(n_627), .C(n_624), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_657), .B(n_622), .Y(n_665) );
NOR2xp33_ASAP7_75t_R g666 ( .A(n_657), .B(n_620), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_655), .B(n_602), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_650), .A2(n_622), .B1(n_634), .B2(n_602), .C(n_631), .Y(n_668) );
INVxp33_ASAP7_75t_SL g669 ( .A(n_644), .Y(n_669) );
AOI32xp33_ASAP7_75t_L g670 ( .A1(n_641), .A2(n_634), .A3(n_495), .B1(n_594), .B2(n_68), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_638), .A2(n_233), .B1(n_255), .B2(n_253), .C(n_234), .Y(n_671) );
XNOR2x2_ASAP7_75t_L g672 ( .A(n_652), .B(n_61), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_207), .B1(n_291), .B2(n_270), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_658), .B(n_253), .C(n_66), .D(n_69), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_649), .B(n_270), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_654), .A2(n_270), .B1(n_291), .B2(n_651), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_655), .A2(n_291), .B(n_647), .C(n_649), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_653), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_653), .A2(n_637), .B1(n_648), .B2(n_654), .C(n_640), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_659), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_666), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_679), .B(n_660), .C(n_677), .Y(n_682) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_669), .A2(n_678), .B1(n_663), .B2(n_665), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_674), .A2(n_661), .B(n_664), .C(n_667), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_684), .B(n_676), .Y(n_685) );
OAI322xp33_ASAP7_75t_L g686 ( .A1(n_683), .A2(n_672), .A3(n_673), .B1(n_659), .B2(n_637), .C1(n_648), .C2(n_670), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_680), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_685), .A2(n_681), .B(n_682), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_686), .A2(n_662), .B(n_668), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_688), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_687), .B1(n_689), .B2(n_675), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_671), .B(n_653), .Y(n_692) );
endmodule