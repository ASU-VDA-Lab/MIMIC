module real_jpeg_26046_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.C(n_37),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_22),
.B1(n_33),
.B2(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_22),
.B1(n_35),
.B2(n_45),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_22),
.B1(n_54),
.B2(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_6),
.B(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_53),
.C(n_55),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_23),
.C(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_6),
.B(n_144),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_98),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_97),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.C(n_80),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_16),
.A2(n_17),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_38),
.B1(n_39),
.B2(n_62),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_18),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_19),
.A2(n_20),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_50),
.C(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_19),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_19),
.A2(n_20),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_19),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_19),
.A2(n_20),
.B1(n_110),
.B2(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_20),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_20),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_20),
.B(n_79),
.C(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_23),
.A2(n_25),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_23),
.B(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_27),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_27),
.A2(n_69),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_29),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_37),
.B1(n_44),
.B2(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_45),
.B1(n_53),
.B2(n_57),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_35),
.B(n_112),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_38),
.A2(n_39),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_50),
.B2(n_61),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_40),
.A2(n_41),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI211xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_71),
.B(n_81),
.C(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_50),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_49),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_61),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_50),
.A2(n_61),
.B1(n_71),
.B2(n_79),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_50),
.A2(n_71),
.B(n_81),
.C(n_152),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_55),
.B1(n_75),
.B2(n_76),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_79),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_63),
.B(n_80),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_71),
.B2(n_79),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_79),
.B1(n_89),
.B2(n_93),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_71),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_71),
.A2(n_79),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_71),
.A2(n_79),
.B1(n_127),
.B2(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_71),
.A2(n_79),
.B1(n_109),
.B2(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_103),
.C(n_109),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_86),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_166),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_161),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_122),
.B(n_160),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_102),
.B(n_113),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_118),
.C(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_116),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_154),
.B(n_159),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_148),
.B(n_153),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_136),
.B(n_147),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_130),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);


endmodule