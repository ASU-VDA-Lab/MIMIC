module fake_aes_6476_n_1347 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1347);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1347;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g297 ( .A(n_30), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_261), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_15), .Y(n_299) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_249), .B(n_47), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_247), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_164), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_221), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_144), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_132), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_157), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_229), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_281), .B(n_201), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_58), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_239), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_22), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_161), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_244), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_96), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_230), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_141), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_291), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_223), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_196), .B(n_83), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_18), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_9), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_18), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_246), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_31), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_75), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_5), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_101), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_195), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_70), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_216), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_84), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_280), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_176), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_260), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_56), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_243), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_70), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_33), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_168), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_16), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_215), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_288), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_17), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_139), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_55), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_178), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_180), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_4), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_208), .Y(n_352) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_295), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_173), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_273), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_166), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_134), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_26), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_140), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_123), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_160), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_29), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_6), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_5), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_279), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_171), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_90), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_203), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_220), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_19), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_50), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_97), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_84), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_152), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_209), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_117), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_78), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_213), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_185), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_262), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_294), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_293), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g383 ( .A(n_151), .B(n_206), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_197), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_181), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_126), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_31), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_200), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_258), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_292), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_179), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_68), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_90), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_225), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_240), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_250), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_182), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_175), .Y(n_398) );
INVxp33_ASAP7_75t_SL g399 ( .A(n_271), .Y(n_399) );
INVxp33_ASAP7_75t_SL g400 ( .A(n_219), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_46), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_259), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_138), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_282), .B(n_290), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_56), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_71), .Y(n_406) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_127), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_241), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_149), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_276), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_286), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_48), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_140), .B(n_129), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_198), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_8), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_121), .Y(n_416) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_202), .B(n_263), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_238), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_152), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_50), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_174), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_14), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_151), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_89), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_141), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_147), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_74), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_194), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_93), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_118), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_36), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_46), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_117), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_17), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_40), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_222), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_157), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_130), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_237), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_132), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_224), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_3), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_144), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_284), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_199), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_63), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_135), .Y(n_447) );
BUFx10_ASAP7_75t_L g448 ( .A(n_272), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_268), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_283), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_53), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_106), .B(n_275), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_51), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_81), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_110), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_234), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_19), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_211), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_76), .Y(n_459) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_21), .B(n_68), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_233), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_59), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_9), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_189), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_21), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_133), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_312), .B(n_0), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_387), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_334), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_312), .B(n_0), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
OAI21x1_ASAP7_75t_L g473 ( .A1(n_395), .A2(n_163), .B(n_162), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_387), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_387), .B(n_1), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_356), .B(n_1), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_298), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_421), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_334), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_421), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_298), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_433), .B(n_2), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_353), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_428), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_395), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_448), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_356), .B(n_6), .Y(n_493) );
INVx5_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
INVx5_ASAP7_75t_L g495 ( .A(n_345), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_299), .B(n_7), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_344), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_398), .B(n_7), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_345), .Y(n_499) );
OAI22x1_ASAP7_75t_R g500 ( .A1(n_314), .A2(n_11), .B1(n_8), .B2(n_10), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_322), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_355), .Y(n_502) );
OAI21x1_ASAP7_75t_L g503 ( .A1(n_355), .A2(n_167), .B(n_165), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_302), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_439), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_447), .B(n_12), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_302), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_439), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_375), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_470), .B(n_401), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_469), .Y(n_511) );
INVx6_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_492), .B(n_335), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_492), .B(n_448), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_420), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_507), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_507), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_507), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_304), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_469), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_478), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_469), .B(n_307), .Y(n_524) );
BUFx8_ASAP7_75t_SL g525 ( .A(n_487), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_484), .A2(n_304), .B1(n_357), .B2(n_305), .Y(n_526) );
NOR2xp33_ASAP7_75t_SL g527 ( .A(n_479), .B(n_301), .Y(n_527) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_475), .B(n_452), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_507), .Y(n_529) );
BUFx8_ASAP7_75t_SL g530 ( .A(n_487), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_489), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_492), .B(n_368), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_492), .B(n_448), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_507), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_485), .B(n_305), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_489), .B(n_310), .Y(n_537) );
NAND2xp33_ASAP7_75t_L g538 ( .A(n_492), .B(n_301), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_492), .B(n_384), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_489), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_479), .B(n_317), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_507), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_475), .Y(n_544) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_475), .B(n_405), .Y(n_546) );
INVx4_ASAP7_75t_SL g547 ( .A(n_475), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_484), .A2(n_346), .B1(n_348), .B2(n_297), .Y(n_548) );
AND2x6_ASAP7_75t_L g549 ( .A(n_496), .B(n_344), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_479), .B(n_303), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_484), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_468), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_483), .B(n_319), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_509), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_468), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_509), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_483), .B(n_320), .Y(n_557) );
BUFx5_ASAP7_75t_L g558 ( .A(n_549), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_528), .A2(n_467), .B1(n_506), .B2(n_476), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_515), .B(n_471), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_528), .A2(n_497), .B1(n_483), .B2(n_496), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_551), .B(n_471), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_551), .B(n_549), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_549), .B(n_476), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_552), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_545), .B(n_496), .Y(n_566) );
OAI22xp5_ASAP7_75t_SL g567 ( .A1(n_554), .A2(n_454), .B1(n_362), .B2(n_501), .Y(n_567) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_526), .B(n_467), .C(n_506), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_545), .A2(n_497), .B(n_496), .C(n_468), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_534), .B(n_493), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_522), .B(n_493), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_545), .B(n_496), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_522), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_520), .B(n_474), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_545), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_536), .B(n_498), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_511), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_527), .B(n_496), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_512), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_513), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_549), .A2(n_499), .B1(n_505), .B2(n_502), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_544), .A2(n_473), .B(n_503), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_550), .B(n_303), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_512), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_357), .Y(n_588) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_544), .A2(n_473), .B(n_503), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_550), .B(n_313), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_547), .B(n_495), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_547), .B(n_495), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_536), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_512), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_514), .B(n_504), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_547), .B(n_313), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
OR2x6_ASAP7_75t_L g599 ( .A(n_556), .B(n_501), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_533), .B(n_399), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_510), .A2(n_501), .B1(n_359), .B2(n_363), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_542), .A2(n_481), .B(n_474), .C(n_374), .Y(n_602) );
OAI22xp5_ASAP7_75t_SL g603 ( .A1(n_526), .A2(n_481), .B1(n_500), .B2(n_360), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_546), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_539), .B(n_474), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_546), .B(n_315), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_556), .A2(n_456), .B1(n_464), .B2(n_352), .Y(n_607) );
BUFx3_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_510), .A2(n_359), .B1(n_363), .B2(n_360), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_516), .B(n_452), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_521), .B(n_495), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_538), .B(n_399), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_516), .B(n_315), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_524), .B(n_318), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_531), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_525), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_542), .A2(n_502), .B1(n_505), .B2(n_499), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_553), .A2(n_502), .B1(n_505), .B2(n_499), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_553), .A2(n_502), .B1(n_505), .B2(n_499), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_537), .B(n_318), .Y(n_622) );
NAND2xp33_ASAP7_75t_L g623 ( .A(n_531), .B(n_507), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_548), .B(n_326), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_530), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_532), .A2(n_508), .B1(n_466), .B2(n_351), .Y(n_627) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_541), .B(n_351), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_541), .A2(n_376), .B1(n_386), .B2(n_367), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_517), .B(n_333), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_517), .B(n_333), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_517), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_518), .A2(n_376), .B1(n_416), .B2(n_386), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_518), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_519), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_519), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_519), .B(n_495), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_529), .B(n_337), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_575), .Y(n_639) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_568), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_568), .A2(n_400), .B1(n_419), .B2(n_416), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_602), .A2(n_430), .B(n_407), .C(n_371), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_585), .A2(n_473), .B(n_503), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_626), .B(n_419), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_617), .B(n_423), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_581), .A2(n_473), .B(n_503), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_561), .A2(n_425), .B1(n_426), .B2(n_423), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_593), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_614), .B(n_425), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_620), .B(n_561), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_572), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_576), .B(n_432), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_595), .A2(n_543), .B(n_535), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_562), .B(n_432), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_598), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_600), .A2(n_508), .B(n_405), .C(n_451), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_588), .B(n_435), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_625), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_603), .B(n_437), .C(n_435), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_569), .B(n_437), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_566), .A2(n_543), .B(n_308), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_594), .Y(n_662) );
NOR2xp67_ASAP7_75t_L g663 ( .A(n_601), .B(n_442), .Y(n_663) );
BUFx6f_ASAP7_75t_SL g664 ( .A(n_599), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_598), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_597), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_566), .A2(n_336), .B(n_331), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_610), .B(n_443), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_609), .A2(n_306), .B(n_311), .C(n_309), .Y(n_669) );
NOR2xp33_ASAP7_75t_SL g670 ( .A(n_558), .B(n_443), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_605), .A2(n_354), .B(n_349), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_577), .Y(n_672) );
INVx4_ASAP7_75t_L g673 ( .A(n_577), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_600), .A2(n_508), .B(n_451), .C(n_349), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_613), .B(n_457), .Y(n_675) );
BUFx2_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_564), .B(n_457), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_559), .A2(n_465), .B1(n_463), .B2(n_342), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_565), .A2(n_508), .B(n_316), .C(n_323), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_607), .B(n_466), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_628), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_629), .B(n_327), .Y(n_682) );
CKINVDCx8_ASAP7_75t_R g683 ( .A(n_577), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_574), .A2(n_329), .B(n_330), .C(n_328), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_573), .A2(n_342), .B1(n_350), .B2(n_339), .Y(n_685) );
INVxp33_ASAP7_75t_SL g686 ( .A(n_567), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_624), .B(n_332), .Y(n_687) );
BUFx8_ASAP7_75t_L g688 ( .A(n_558), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_560), .B(n_340), .C(n_338), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_SL g690 ( .A1(n_570), .A2(n_366), .B(n_385), .C(n_381), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_560), .A2(n_341), .B1(n_364), .B2(n_358), .C(n_343), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_633), .Y(n_692) );
BUFx2_ASAP7_75t_L g693 ( .A(n_573), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_589), .A2(n_391), .B(n_390), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_563), .A2(n_397), .B(n_396), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_628), .Y(n_696) );
OR2x6_ASAP7_75t_L g697 ( .A(n_577), .B(n_500), .Y(n_697) );
INVx8_ASAP7_75t_L g698 ( .A(n_558), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_604), .A2(n_372), .B(n_373), .C(n_370), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_615), .B(n_377), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_622), .B(n_350), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_606), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_571), .B(n_393), .Y(n_703) );
NOR3xp33_ASAP7_75t_SL g704 ( .A(n_571), .B(n_379), .C(n_365), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_612), .A2(n_409), .B(n_412), .C(n_403), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_584), .A2(n_388), .B1(n_389), .B2(n_382), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_618), .B(n_495), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_608), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_631), .A2(n_408), .B(n_402), .Y(n_709) );
AO21x1_ASAP7_75t_L g710 ( .A1(n_611), .A2(n_477), .B(n_472), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_586), .A2(n_422), .B(n_427), .C(n_415), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_618), .B(n_495), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_579), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_619), .B(n_495), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_612), .A2(n_389), .B1(n_410), .B2(n_388), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_619), .A2(n_436), .B1(n_449), .B2(n_410), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_590), .B(n_429), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_582), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_621), .A2(n_431), .B(n_438), .C(n_434), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_621), .A2(n_440), .B(n_453), .C(n_446), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_627), .B(n_455), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_638), .A2(n_418), .B(n_414), .Y(n_722) );
NAND2xp33_ASAP7_75t_SL g723 ( .A(n_591), .B(n_449), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_627), .B(n_459), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_579), .B(n_299), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_580), .B(n_324), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_580), .A2(n_413), .B(n_460), .C(n_321), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_583), .Y(n_728) );
BUFx8_ASAP7_75t_SL g729 ( .A(n_583), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_616), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_587), .Y(n_731) );
AOI21x1_ASAP7_75t_L g732 ( .A1(n_591), .A2(n_417), .B(n_404), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g733 ( .A1(n_616), .A2(n_383), .B(n_300), .C(n_347), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_592), .B(n_324), .Y(n_734) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_596), .A2(n_347), .B(n_406), .C(n_392), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_634), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_592), .B(n_392), .Y(n_737) );
O2A1O1Ixp33_ASAP7_75t_L g738 ( .A1(n_630), .A2(n_424), .B(n_462), .C(n_406), .Y(n_738) );
BUFx8_ASAP7_75t_L g739 ( .A(n_632), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_611), .B(n_424), .Y(n_740) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_637), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_635), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_636), .B(n_450), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_623), .A2(n_507), .B1(n_441), .B2(n_444), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_598), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_578), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_598), .Y(n_747) );
AND2x6_ASAP7_75t_L g748 ( .A(n_577), .B(n_325), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_598), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_594), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_568), .B(n_450), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_568), .A2(n_461), .B1(n_458), .B2(n_445), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_578), .B(n_458), .Y(n_753) );
INVx4_ASAP7_75t_L g754 ( .A(n_577), .Y(n_754) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_577), .Y(n_755) );
BUFx3_ASAP7_75t_L g756 ( .A(n_625), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_568), .B(n_461), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_626), .B(n_361), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_626), .B(n_380), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_626), .B(n_411), .Y(n_760) );
BUFx2_ASAP7_75t_L g761 ( .A(n_575), .Y(n_761) );
O2A1O1Ixp33_ASAP7_75t_L g762 ( .A1(n_705), .A2(n_369), .B(n_378), .C(n_325), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_694), .A2(n_480), .A3(n_488), .B(n_482), .Y(n_763) );
AO31x2_ASAP7_75t_L g764 ( .A1(n_643), .A2(n_488), .A3(n_486), .B(n_478), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_746), .B(n_13), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_719), .A2(n_378), .B(n_394), .C(n_369), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_683), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_739), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_659), .A2(n_394), .B1(n_500), .B2(n_488), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_697), .A2(n_494), .B1(n_16), .B2(n_14), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_651), .B(n_15), .Y(n_771) );
NOR2x1p5_ASAP7_75t_L g772 ( .A(n_658), .B(n_20), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_646), .A2(n_540), .B(n_523), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_739), .Y(n_774) );
O2A1O1Ixp5_ASAP7_75t_L g775 ( .A1(n_656), .A2(n_488), .B(n_494), .C(n_486), .Y(n_775) );
NOR2xp67_ASAP7_75t_SL g776 ( .A(n_696), .B(n_494), .Y(n_776) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_672), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_SL g778 ( .A1(n_674), .A2(n_170), .B(n_172), .C(n_169), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_736), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_650), .A2(n_494), .B1(n_486), .B2(n_490), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_737), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_713), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_697), .A2(n_494), .B1(n_23), .B2(n_20), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_728), .Y(n_784) );
BUFx3_ASAP7_75t_L g785 ( .A(n_729), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_730), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_648), .A2(n_494), .B1(n_486), .B2(n_490), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_734), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_653), .A2(n_540), .B(n_523), .Y(n_789) );
NOR2x1_ASAP7_75t_L g790 ( .A(n_697), .B(n_478), .Y(n_790) );
INVxp67_ASAP7_75t_L g791 ( .A(n_639), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_734), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_649), .B(n_23), .Y(n_793) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_707), .A2(n_494), .B(n_486), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_681), .B(n_24), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_756), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g797 ( .A1(n_720), .A2(n_26), .B(n_24), .C(n_25), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_644), .B(n_25), .Y(n_798) );
AND2x4_ASAP7_75t_SL g799 ( .A(n_668), .B(n_478), .Y(n_799) );
AO22x1_ASAP7_75t_L g800 ( .A1(n_686), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_661), .A2(n_540), .B(n_523), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_725), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_664), .A2(n_490), .B1(n_491), .B2(n_478), .Y(n_803) );
O2A1O1Ixp33_ASAP7_75t_L g804 ( .A1(n_684), .A2(n_30), .B(n_27), .C(n_28), .Y(n_804) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_645), .Y(n_805) );
OAI22x1_ASAP7_75t_SL g806 ( .A1(n_692), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_742), .Y(n_807) );
A2O1A1Ixp33_ASAP7_75t_L g808 ( .A1(n_703), .A2(n_711), .B(n_722), .C(n_709), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_712), .A2(n_491), .B(n_490), .Y(n_809) );
AO22x2_ASAP7_75t_L g810 ( .A1(n_678), .A2(n_35), .B1(n_32), .B2(n_34), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_650), .A2(n_491), .B1(n_490), .B2(n_37), .Y(n_811) );
INVxp67_ASAP7_75t_L g812 ( .A(n_761), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_665), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_673), .Y(n_814) );
AO32x2_ASAP7_75t_L g815 ( .A1(n_702), .A2(n_491), .A3(n_36), .B1(n_37), .B2(n_38), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_666), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_664), .A2(n_491), .B1(n_39), .B2(n_35), .Y(n_817) );
O2A1O1Ixp33_ASAP7_75t_L g818 ( .A1(n_642), .A2(n_40), .B(n_38), .C(n_39), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_753), .B(n_41), .Y(n_819) );
BUFx3_ASAP7_75t_L g820 ( .A(n_693), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g821 ( .A1(n_679), .A2(n_43), .B(n_41), .C(n_42), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_725), .Y(n_822) );
OAI21x1_ASAP7_75t_L g823 ( .A1(n_732), .A2(n_183), .B(n_177), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_714), .A2(n_42), .B(n_43), .Y(n_824) );
AO31x2_ASAP7_75t_L g825 ( .A1(n_727), .A2(n_47), .A3(n_44), .B(n_45), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_655), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_654), .B(n_44), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_677), .A2(n_186), .B(n_184), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_748), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_726), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_726), .A2(n_49), .B1(n_45), .B2(n_48), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_714), .A2(n_49), .B(n_51), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_673), .B(n_52), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_685), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_676), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_760), .A2(n_188), .B(n_187), .Y(n_836) );
INVx1_ASAP7_75t_SL g837 ( .A(n_748), .Y(n_837) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_641), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_745), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_647), .B(n_52), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_710), .A2(n_191), .B(n_190), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_747), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_657), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_654), .B(n_54), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_759), .A2(n_193), .B(n_192), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_754), .Y(n_846) );
AND2x6_ASAP7_75t_L g847 ( .A(n_672), .B(n_57), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_660), .A2(n_57), .B(n_58), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_740), .Y(n_849) );
A2O1A1Ixp33_ASAP7_75t_L g850 ( .A1(n_738), .A2(n_59), .B(n_60), .C(n_61), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_689), .B(n_60), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_748), .Y(n_852) );
AO32x2_ASAP7_75t_L g853 ( .A1(n_752), .A2(n_61), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_749), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_663), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_740), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_759), .Y(n_857) );
INVx4_ASAP7_75t_L g858 ( .A(n_672), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_704), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_760), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_718), .Y(n_861) );
AOI221xp5_ASAP7_75t_SL g862 ( .A1(n_733), .A2(n_65), .B1(n_66), .B2(n_67), .C(n_69), .Y(n_862) );
INVx2_ASAP7_75t_SL g863 ( .A(n_721), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_735), .A2(n_67), .B(n_69), .C(n_71), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_669), .A2(n_72), .B(n_73), .C(n_74), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_695), .A2(n_758), .B(n_701), .Y(n_866) );
INVx1_ASAP7_75t_SL g867 ( .A(n_748), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_724), .A2(n_72), .B1(n_73), .B2(n_75), .Y(n_868) );
O2A1O1Ixp33_ASAP7_75t_L g869 ( .A1(n_699), .A2(n_76), .B(n_77), .C(n_78), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_671), .A2(n_77), .B(n_79), .Y(n_870) );
O2A1O1Ixp33_ASAP7_75t_L g871 ( .A1(n_690), .A2(n_79), .B(n_80), .C(n_81), .Y(n_871) );
INVx3_ASAP7_75t_L g872 ( .A(n_754), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_675), .B(n_80), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_731), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_680), .A2(n_82), .B1(n_83), .B2(n_85), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_682), .A2(n_82), .B1(n_85), .B2(n_86), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_715), .B(n_86), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_700), .B(n_87), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_687), .B(n_87), .Y(n_879) );
O2A1O1Ixp5_ASAP7_75t_L g880 ( .A1(n_717), .A2(n_212), .B(n_289), .C(n_287), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_652), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_652), .B(n_88), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_716), .A2(n_88), .B1(n_89), .B2(n_91), .Y(n_883) );
INVx6_ASAP7_75t_L g884 ( .A(n_688), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_691), .B(n_92), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_724), .B(n_93), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_743), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_887) );
AO31x2_ASAP7_75t_L g888 ( .A1(n_667), .A2(n_98), .A3(n_99), .B(n_100), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_640), .B(n_98), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_688), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_706), .B(n_102), .Y(n_891) );
OAI21x1_ASAP7_75t_L g892 ( .A1(n_708), .A2(n_217), .B(n_285), .Y(n_892) );
AO31x2_ASAP7_75t_L g893 ( .A1(n_748), .A2(n_103), .A3(n_104), .B(n_105), .Y(n_893) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_670), .B(n_104), .C(n_105), .Y(n_894) );
BUFx10_ASAP7_75t_L g895 ( .A(n_741), .Y(n_895) );
OAI22x1_ASAP7_75t_L g896 ( .A1(n_751), .A2(n_106), .B1(n_107), .B2(n_108), .Y(n_896) );
BUFx6f_ASAP7_75t_L g897 ( .A(n_755), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_757), .B(n_107), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_662), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_750), .B(n_109), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_750), .Y(n_901) );
O2A1O1Ixp33_ASAP7_75t_L g902 ( .A1(n_744), .A2(n_111), .B(n_112), .C(n_113), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_723), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_755), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_741), .B(n_114), .Y(n_905) );
AOI211xp5_ASAP7_75t_L g906 ( .A1(n_770), .A2(n_783), .B(n_800), .C(n_878), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_863), .A2(n_698), .B1(n_116), .B2(n_118), .Y(n_907) );
OR2x2_ASAP7_75t_L g908 ( .A(n_791), .B(n_115), .Y(n_908) );
BUFx2_ASAP7_75t_L g909 ( .A(n_796), .Y(n_909) );
A2O1A1Ixp33_ASAP7_75t_L g910 ( .A1(n_808), .A2(n_698), .B(n_120), .C(n_121), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_805), .Y(n_911) );
A2O1A1Ixp33_ASAP7_75t_L g912 ( .A1(n_873), .A2(n_698), .B(n_120), .C(n_122), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g913 ( .A1(n_773), .A2(n_231), .B(n_277), .Y(n_913) );
A2O1A1Ixp33_ASAP7_75t_L g914 ( .A1(n_866), .A2(n_119), .B(n_122), .C(n_123), .Y(n_914) );
AO31x2_ASAP7_75t_L g915 ( .A1(n_780), .A2(n_119), .A3(n_124), .B(n_125), .Y(n_915) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_769), .A2(n_124), .B1(n_125), .B2(n_126), .C(n_127), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_857), .B(n_128), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_789), .A2(n_236), .B(n_274), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_812), .Y(n_919) );
BUFx2_ASAP7_75t_L g920 ( .A(n_795), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_816), .Y(n_921) );
NAND2x1p5_ASAP7_75t_L g922 ( .A(n_776), .B(n_128), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_838), .A2(n_129), .B1(n_130), .B2(n_131), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_860), .A2(n_131), .B1(n_133), .B2(n_134), .Y(n_924) );
AND2x4_ASAP7_75t_L g925 ( .A(n_820), .B(n_135), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_795), .B(n_136), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_807), .Y(n_927) );
AO21x2_ASAP7_75t_L g928 ( .A1(n_809), .A2(n_235), .B(n_270), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_765), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_795), .A2(n_136), .B1(n_137), .B2(n_138), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_877), .A2(n_137), .B1(n_139), .B2(n_142), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_785), .B(n_142), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_861), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_802), .B(n_143), .Y(n_934) );
AOI21x1_ASAP7_75t_L g935 ( .A1(n_780), .A2(n_242), .B(n_269), .Y(n_935) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_766), .A2(n_143), .B(n_145), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_782), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_771), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_810), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_822), .B(n_145), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_810), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_891), .A2(n_146), .B1(n_147), .B2(n_148), .Y(n_942) );
AOI21xp33_ASAP7_75t_L g943 ( .A1(n_811), .A2(n_146), .B(n_148), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_830), .B(n_149), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_881), .B(n_150), .Y(n_945) );
INVx4_ASAP7_75t_L g946 ( .A(n_774), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_819), .B(n_150), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_890), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_868), .Y(n_949) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_777), .Y(n_950) );
BUFx3_ASAP7_75t_L g951 ( .A(n_884), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_868), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_762), .A2(n_869), .B(n_848), .C(n_818), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_831), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_772), .B(n_153), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_835), .B(n_153), .Y(n_956) );
AO21x2_ASAP7_75t_L g957 ( .A1(n_811), .A2(n_248), .B(n_267), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_784), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_885), .A2(n_154), .B1(n_155), .B2(n_156), .C(n_158), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_831), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_843), .A2(n_154), .B(n_155), .C(n_156), .Y(n_961) );
AND2x4_ASAP7_75t_L g962 ( .A(n_781), .B(n_158), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_849), .B(n_159), .Y(n_963) );
BUFx3_ASAP7_75t_L g964 ( .A(n_767), .Y(n_964) );
AO22x1_ASAP7_75t_L g965 ( .A1(n_847), .A2(n_159), .B1(n_204), .B2(n_205), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_851), .A2(n_207), .B1(n_210), .B2(n_214), .C(n_218), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_855), .A2(n_226), .B1(n_227), .B2(n_228), .C(n_232), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_856), .B(n_251), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_788), .B(n_792), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_834), .B(n_252), .Y(n_970) );
AOI21xp5_ASAP7_75t_L g971 ( .A1(n_794), .A2(n_253), .B(n_254), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_840), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_896), .Y(n_973) );
BUFx12f_ASAP7_75t_L g974 ( .A(n_847), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_859), .A2(n_264), .B1(n_265), .B2(n_266), .Y(n_975) );
A2O1A1Ixp33_ASAP7_75t_L g976 ( .A1(n_848), .A2(n_865), .B(n_797), .C(n_804), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_882), .Y(n_977) );
OA21x2_ASAP7_75t_L g978 ( .A1(n_892), .A2(n_841), .B(n_823), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_793), .A2(n_798), .B1(n_827), .B2(n_844), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_786), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_900), .A2(n_790), .B1(n_879), .B2(n_898), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g982 ( .A1(n_794), .A2(n_778), .B(n_828), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_833), .A2(n_824), .B1(n_832), .B2(n_886), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_833), .Y(n_984) );
A2O1A1Ixp33_ASAP7_75t_L g985 ( .A1(n_821), .A2(n_871), .B(n_902), .C(n_832), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_870), .Y(n_986) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_775), .A2(n_862), .B(n_880), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_779), .Y(n_988) );
AO31x2_ASAP7_75t_L g989 ( .A1(n_864), .A2(n_850), .A3(n_836), .B(n_845), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_870), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_824), .A2(n_799), .B1(n_894), .B2(n_883), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g992 ( .A(n_806), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_767), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_876), .A2(n_904), .B1(n_852), .B2(n_867), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_875), .B(n_854), .Y(n_995) );
BUFx4f_ASAP7_75t_SL g996 ( .A(n_847), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_888), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g998 ( .A1(n_862), .A2(n_887), .B1(n_817), .B2(n_903), .C(n_899), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_904), .A2(n_829), .B1(n_867), .B2(n_852), .Y(n_999) );
OAI321xp33_ASAP7_75t_L g1000 ( .A1(n_889), .A2(n_787), .A3(n_905), .B1(n_803), .B2(n_842), .C(n_839), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_829), .A2(n_837), .B1(n_872), .B2(n_846), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_826), .A2(n_901), .B1(n_813), .B2(n_846), .C(n_872), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1003 ( .A1(n_847), .A2(n_814), .B1(n_837), .B2(n_858), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_853), .B(n_815), .Y(n_1004) );
AOI21xp5_ASAP7_75t_L g1005 ( .A1(n_777), .A2(n_897), .B(n_858), .Y(n_1005) );
BUFx8_ASAP7_75t_L g1006 ( .A(n_853), .Y(n_1006) );
A2O1A1Ixp33_ASAP7_75t_L g1007 ( .A1(n_853), .A2(n_825), .B(n_893), .C(n_763), .Y(n_1007) );
AOI21xp5_ASAP7_75t_L g1008 ( .A1(n_764), .A2(n_773), .B(n_789), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_874), .Y(n_1009) );
INVx4_ASAP7_75t_L g1010 ( .A(n_768), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_834), .B(n_686), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_773), .A2(n_789), .B(n_801), .Y(n_1012) );
INVx3_ASAP7_75t_L g1013 ( .A(n_895), .Y(n_1013) );
OAI21xp33_ASAP7_75t_L g1014 ( .A1(n_873), .A2(n_550), .B(n_527), .Y(n_1014) );
OAI21xp5_ASAP7_75t_SL g1015 ( .A1(n_769), .A2(n_607), .B(n_686), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_857), .B(n_650), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_838), .A2(n_599), .B1(n_697), .B2(n_659), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_857), .B(n_650), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_857), .B(n_746), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_874), .Y(n_1020) );
NOR2xp67_ASAP7_75t_L g1021 ( .A(n_890), .B(n_768), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_773), .A2(n_789), .B(n_801), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_857), .B(n_650), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_863), .A2(n_568), .B1(n_561), .B2(n_795), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_791), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_773), .A2(n_789), .B(n_801), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_857), .B(n_650), .Y(n_1027) );
OAI22xp33_ASAP7_75t_L g1028 ( .A1(n_795), .A2(n_697), .B1(n_599), .B2(n_568), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_874), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_773), .A2(n_789), .B(n_801), .Y(n_1030) );
INVx3_ASAP7_75t_L g1031 ( .A(n_895), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_857), .B(n_696), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_838), .A2(n_599), .B1(n_697), .B2(n_659), .Y(n_1033) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_796), .Y(n_1034) );
OA21x2_ASAP7_75t_L g1035 ( .A1(n_1008), .A2(n_1007), .B(n_1012), .Y(n_1035) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_909), .Y(n_1036) );
BUFx2_ASAP7_75t_SL g1037 ( .A(n_1021), .Y(n_1037) );
AOI33xp33_ASAP7_75t_L g1038 ( .A1(n_939), .A2(n_941), .A3(n_955), .B1(n_1017), .B2(n_1033), .B3(n_973), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_1025), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_919), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1041 ( .A1(n_1015), .A2(n_906), .B1(n_1024), .B2(n_953), .C(n_976), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_937), .B(n_958), .Y(n_1042) );
OA21x2_ASAP7_75t_L g1043 ( .A1(n_1022), .A2(n_1030), .B(n_1026), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_980), .B(n_988), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_997), .Y(n_1045) );
AND2x4_ASAP7_75t_L g1046 ( .A(n_984), .B(n_969), .Y(n_1046) );
NOR2xp33_ASAP7_75t_L g1047 ( .A(n_1011), .B(n_920), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1019), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1024), .B(n_949), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_969), .B(n_950), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_996), .A2(n_930), .B1(n_974), .B2(n_1006), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_952), .B(n_954), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1009), .Y(n_1053) );
AND2x4_ASAP7_75t_SL g1054 ( .A(n_946), .B(n_1010), .Y(n_1054) );
OR2x6_ASAP7_75t_L g1055 ( .A(n_922), .B(n_965), .Y(n_1055) );
AO21x2_ASAP7_75t_L g1056 ( .A1(n_983), .A2(n_982), .B(n_990), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1020), .Y(n_1057) );
AO21x2_ASAP7_75t_L g1058 ( .A1(n_983), .A2(n_986), .B(n_910), .Y(n_1058) );
OR2x6_ASAP7_75t_L g1059 ( .A(n_922), .B(n_999), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_1028), .B(n_1032), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1004), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_960), .A2(n_907), .B1(n_930), .B2(n_962), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_907), .A2(n_926), .B1(n_962), .B2(n_916), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1064 ( .A1(n_1006), .A2(n_925), .B1(n_970), .B2(n_991), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1016), .B(n_1018), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1029), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_921), .B(n_933), .Y(n_1067) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_911), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_1034), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_915), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_925), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_915), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_927), .B(n_1016), .Y(n_1073) );
AO21x2_ASAP7_75t_L g1074 ( .A1(n_985), .A2(n_936), .B(n_943), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1018), .B(n_1023), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1023), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1027), .B(n_934), .Y(n_1077) );
NAND2xp5_ASAP7_75t_SL g1078 ( .A(n_1003), .B(n_943), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_977), .B(n_1027), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_999), .B(n_991), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_995), .B(n_934), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_917), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_917), .Y(n_1083) );
OR2x6_ASAP7_75t_L g1084 ( .A(n_994), .B(n_1001), .Y(n_1084) );
OAI321xp33_ASAP7_75t_L g1085 ( .A1(n_916), .A2(n_998), .A3(n_961), .B1(n_931), .B2(n_967), .C(n_923), .Y(n_1085) );
OA21x2_ASAP7_75t_L g1086 ( .A1(n_979), .A2(n_914), .B(n_935), .Y(n_1086) );
OR2x6_ASAP7_75t_L g1087 ( .A(n_994), .B(n_1001), .Y(n_1087) );
AOI321xp33_ASAP7_75t_L g1088 ( .A1(n_942), .A2(n_959), .A3(n_998), .B1(n_924), .B2(n_938), .C(n_929), .Y(n_1088) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_951), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_940), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_940), .B(n_944), .Y(n_1091) );
OAI21xp5_ASAP7_75t_SL g1092 ( .A1(n_912), .A2(n_932), .B(n_975), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_944), .B(n_963), .Y(n_1093) );
OAI21xp5_ASAP7_75t_SL g1094 ( .A1(n_948), .A2(n_1014), .B(n_947), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_963), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_945), .B(n_956), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_945), .B(n_1031), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_908), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1013), .B(n_1031), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1013), .B(n_957), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1002), .B(n_968), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1102 ( .A(n_1005), .B(n_928), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_992), .A2(n_993), .B1(n_981), .B2(n_964), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_989), .B(n_987), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_946), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_989), .B(n_1010), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_989), .B(n_972), .Y(n_1107) );
INVx2_ASAP7_75t_L g1108 ( .A(n_978), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1109 ( .A(n_966), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_971), .B(n_918), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_913), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1000), .Y(n_1112) );
AO21x2_ASAP7_75t_L g1113 ( .A1(n_1007), .A2(n_1008), .B(n_1030), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_997), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_996), .Y(n_1115) );
OA21x2_ASAP7_75t_L g1116 ( .A1(n_1008), .A2(n_1007), .B(n_1012), .Y(n_1116) );
INVx2_ASAP7_75t_SL g1117 ( .A(n_996), .Y(n_1117) );
BUFx2_ASAP7_75t_SL g1118 ( .A(n_1021), .Y(n_1118) );
OR2x6_ASAP7_75t_L g1119 ( .A(n_974), .B(n_795), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_911), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_939), .B(n_941), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_919), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1024), .A2(n_996), .B1(n_795), .B2(n_1028), .Y(n_1123) );
OA21x2_ASAP7_75t_L g1124 ( .A1(n_1008), .A2(n_1007), .B(n_1012), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_919), .Y(n_1125) );
OA21x2_ASAP7_75t_L g1126 ( .A1(n_1008), .A2(n_1007), .B(n_1012), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1121), .B(n_1061), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_1036), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1061), .B(n_1080), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_1100), .B(n_1106), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1045), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1080), .B(n_1049), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1045), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1080), .B(n_1049), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1080), .B(n_1052), .Y(n_1135) );
BUFx3_ASAP7_75t_L g1136 ( .A(n_1036), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1052), .B(n_1075), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1108), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1114), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1073), .B(n_1075), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1073), .B(n_1067), .Y(n_1141) );
INVxp67_ASAP7_75t_L g1142 ( .A(n_1040), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1121), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1106), .B(n_1081), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1066), .B(n_1081), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1070), .B(n_1072), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1072), .B(n_1096), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1042), .B(n_1044), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_1122), .Y(n_1149) );
INVx3_ASAP7_75t_SL g1150 ( .A(n_1054), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1096), .B(n_1065), .Y(n_1151) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1100), .B(n_1059), .Y(n_1152) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_1059), .Y(n_1153) );
NAND2x1p5_ASAP7_75t_L g1154 ( .A(n_1046), .B(n_1050), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1077), .B(n_1084), .Y(n_1155) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_1059), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_1041), .A2(n_1123), .B1(n_1064), .B2(n_1063), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1079), .B(n_1048), .Y(n_1158) );
INVx1_ASAP7_75t_SL g1159 ( .A(n_1069), .Y(n_1159) );
HB1xp67_ASAP7_75t_L g1160 ( .A(n_1125), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1084), .B(n_1087), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1039), .Y(n_1162) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_1059), .B(n_1084), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1046), .B(n_1076), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1095), .B(n_1091), .Y(n_1165) );
AND2x4_ASAP7_75t_L g1166 ( .A(n_1084), .B(n_1087), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1087), .B(n_1058), .Y(n_1167) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_1069), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1058), .B(n_1050), .Y(n_1169) );
INVxp67_ASAP7_75t_SL g1170 ( .A(n_1050), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1053), .B(n_1057), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1071), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1082), .B(n_1083), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1091), .B(n_1093), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1043), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1038), .B(n_1093), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1090), .B(n_1098), .Y(n_1177) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_1097), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1179 ( .A(n_1099), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1104), .B(n_1062), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1043), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1043), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1043), .Y(n_1183) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_1099), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1107), .B(n_1113), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1107), .B(n_1113), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_1128), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1174), .B(n_1094), .Y(n_1188) );
INVx1_ASAP7_75t_SL g1189 ( .A(n_1150), .Y(n_1189) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1138), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1129), .B(n_1113), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1129), .B(n_1035), .Y(n_1192) );
AND2x4_ASAP7_75t_L g1193 ( .A(n_1169), .B(n_1102), .Y(n_1193) );
NAND3xp33_ASAP7_75t_L g1194 ( .A(n_1157), .B(n_1092), .C(n_1051), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1185), .B(n_1035), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1185), .B(n_1035), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1186), .B(n_1035), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1186), .B(n_1126), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1144), .B(n_1104), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1144), .B(n_1126), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1132), .B(n_1126), .Y(n_1201) );
AND2x4_ASAP7_75t_SL g1202 ( .A(n_1163), .B(n_1055), .Y(n_1202) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1128), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1204 ( .A(n_1150), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1132), .B(n_1126), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1137), .B(n_1060), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1134), .B(n_1124), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1145), .B(n_1101), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1134), .B(n_1124), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1131), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g1211 ( .A1(n_1150), .A2(n_1103), .B1(n_1119), .B2(n_1088), .C(n_1142), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1141), .B(n_1047), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1131), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1133), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_1162), .B(n_1078), .C(n_1055), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1135), .B(n_1130), .Y(n_1216) );
NAND2x1p5_ASAP7_75t_L g1217 ( .A(n_1128), .B(n_1115), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1135), .B(n_1124), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1133), .Y(n_1219) );
INVxp67_ASAP7_75t_L g1220 ( .A(n_1149), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_1136), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1139), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1139), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1148), .B(n_1074), .Y(n_1224) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1160), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1169), .B(n_1116), .Y(n_1226) );
NOR2x1_ASAP7_75t_SL g1227 ( .A(n_1136), .B(n_1055), .Y(n_1227) );
NAND2x1_ASAP7_75t_L g1228 ( .A(n_1153), .B(n_1055), .Y(n_1228) );
NAND2xp5_ASAP7_75t_SL g1229 ( .A(n_1159), .B(n_1115), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1180), .B(n_1056), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1189), .B(n_1105), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1201), .B(n_1167), .Y(n_1232) );
NAND2x1_ASAP7_75t_L g1233 ( .A(n_1215), .B(n_1187), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1202), .B(n_1163), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1210), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1225), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1210), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1208), .B(n_1171), .Y(n_1238) );
NAND2xp5_ASAP7_75t_SL g1239 ( .A(n_1215), .B(n_1159), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1221), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1213), .Y(n_1241) );
AND2x4_ASAP7_75t_L g1242 ( .A(n_1202), .B(n_1163), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1213), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1205), .B(n_1166), .Y(n_1244) );
INVx3_ASAP7_75t_SL g1245 ( .A(n_1204), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1246 ( .A1(n_1194), .A2(n_1176), .B1(n_1119), .B2(n_1166), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1224), .B(n_1147), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1214), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1207), .B(n_1166), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1207), .B(n_1166), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1214), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1219), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1209), .B(n_1152), .Y(n_1253) );
NAND2xp5_ASAP7_75t_SL g1254 ( .A(n_1203), .B(n_1136), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1209), .B(n_1152), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1199), .B(n_1155), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1194), .B(n_1089), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_L g1258 ( .A1(n_1228), .A2(n_1037), .B(n_1118), .C(n_1054), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1222), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1211), .A2(n_1119), .B1(n_1156), .B2(n_1178), .Y(n_1260) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1190), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1218), .B(n_1152), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1218), .B(n_1152), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1222), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1223), .Y(n_1265) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1199), .B(n_1155), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1195), .B(n_1163), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1200), .B(n_1127), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1195), .B(n_1146), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1196), .B(n_1146), .Y(n_1270) );
NOR2xp33_ASAP7_75t_L g1271 ( .A(n_1257), .B(n_1220), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1269), .B(n_1216), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_1260), .A2(n_1161), .B1(n_1156), .B2(n_1188), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1268), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1269), .B(n_1196), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1268), .Y(n_1276) );
OAI332xp33_ASAP7_75t_L g1277 ( .A1(n_1236), .A2(n_1177), .A3(n_1212), .B1(n_1151), .B2(n_1230), .B3(n_1158), .C1(n_1165), .C2(n_1206), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1245), .B(n_1229), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1270), .B(n_1197), .Y(n_1279) );
NOR2xp33_ASAP7_75t_SL g1280 ( .A(n_1245), .B(n_1037), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1270), .B(n_1216), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1235), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1235), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1247), .B(n_1200), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1237), .Y(n_1285) );
INVx3_ASAP7_75t_L g1286 ( .A(n_1234), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1234), .B(n_1193), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1237), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1289 ( .A(n_1240), .Y(n_1289) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_1258), .A2(n_1227), .B(n_1202), .Y(n_1290) );
AND2x2_ASAP7_75t_SL g1291 ( .A(n_1242), .B(n_1161), .Y(n_1291) );
AOI221xp5_ASAP7_75t_L g1292 ( .A1(n_1238), .A2(n_1143), .B1(n_1172), .B2(n_1165), .C(n_1198), .Y(n_1292) );
INVxp67_ASAP7_75t_SL g1293 ( .A(n_1239), .Y(n_1293) );
AOI21xp33_ASAP7_75t_SL g1294 ( .A1(n_1254), .A2(n_1217), .B(n_1227), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1241), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1232), .B(n_1198), .Y(n_1296) );
OAI22x1_ASAP7_75t_L g1297 ( .A1(n_1242), .A2(n_1217), .B1(n_1193), .B2(n_1120), .Y(n_1297) );
OAI22xp33_ASAP7_75t_L g1298 ( .A1(n_1280), .A2(n_1246), .B1(n_1233), .B2(n_1168), .Y(n_1298) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_1271), .A2(n_1267), .B1(n_1231), .B2(n_1244), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1274), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1277), .B(n_1232), .Y(n_1301) );
AOI322xp5_ASAP7_75t_L g1302 ( .A1(n_1271), .A2(n_1293), .A3(n_1292), .B1(n_1278), .B2(n_1276), .C1(n_1296), .C2(n_1273), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1284), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1282), .Y(n_1304) );
AOI211xp5_ASAP7_75t_SL g1305 ( .A1(n_1290), .A2(n_1242), .B(n_1085), .C(n_1179), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1283), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1285), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1288), .Y(n_1308) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1295), .Y(n_1309) );
OAI211xp5_ASAP7_75t_L g1310 ( .A1(n_1294), .A2(n_1168), .B(n_1256), .C(n_1266), .Y(n_1310) );
AOI21xp5_ASAP7_75t_SL g1311 ( .A1(n_1297), .A2(n_1117), .B(n_1151), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1304), .Y(n_1312) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_1302), .A2(n_1273), .B1(n_1278), .B2(n_1286), .C(n_1289), .Y(n_1313) );
AOI322xp5_ASAP7_75t_L g1314 ( .A1(n_1301), .A2(n_1275), .A3(n_1279), .B1(n_1291), .B2(n_1281), .C1(n_1272), .C2(n_1286), .Y(n_1314) );
AOI222xp33_ASAP7_75t_L g1315 ( .A1(n_1310), .A2(n_1191), .B1(n_1287), .B2(n_1267), .C1(n_1226), .C2(n_1244), .Y(n_1315) );
OAI22xp5_ASAP7_75t_SL g1316 ( .A1(n_1311), .A2(n_1068), .B1(n_1120), .B2(n_1118), .Y(n_1316) );
OAI21xp5_ASAP7_75t_L g1317 ( .A1(n_1305), .A2(n_1287), .B(n_1068), .Y(n_1317) );
OAI21xp5_ASAP7_75t_L g1318 ( .A1(n_1311), .A2(n_1287), .B(n_1109), .Y(n_1318) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1309), .Y(n_1319) );
OAI31xp33_ASAP7_75t_SL g1320 ( .A1(n_1298), .A2(n_1262), .A3(n_1253), .B(n_1255), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1306), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1299), .B(n_1249), .Y(n_1322) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_1303), .A2(n_1250), .B1(n_1263), .B2(n_1262), .Y(n_1323) );
AOI211xp5_ASAP7_75t_SL g1324 ( .A1(n_1316), .A2(n_1300), .B(n_1177), .C(n_1173), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1314), .B(n_1307), .Y(n_1325) );
AO31x2_ASAP7_75t_L g1326 ( .A1(n_1312), .A2(n_1321), .A3(n_1322), .B(n_1319), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1317), .B(n_1308), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_1313), .A2(n_1309), .B1(n_1251), .B2(n_1252), .C(n_1243), .Y(n_1328) );
NAND3xp33_ASAP7_75t_L g1329 ( .A(n_1315), .B(n_1265), .C(n_1264), .Y(n_1329) );
NAND3xp33_ASAP7_75t_L g1330 ( .A(n_1320), .B(n_1248), .C(n_1259), .Y(n_1330) );
A2O1A1Ixp33_ASAP7_75t_L g1331 ( .A1(n_1324), .A2(n_1318), .B(n_1322), .C(n_1323), .Y(n_1331) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1328), .B(n_1086), .C(n_1183), .Y(n_1332) );
INVx3_ASAP7_75t_L g1333 ( .A(n_1326), .Y(n_1333) );
OAI22x1_ASAP7_75t_L g1334 ( .A1(n_1327), .A2(n_1112), .B1(n_1154), .B2(n_1184), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1331), .B(n_1325), .C(n_1329), .Y(n_1335) );
NOR2xp67_ASAP7_75t_L g1336 ( .A(n_1333), .B(n_1330), .Y(n_1336) );
AND4x1_ASAP7_75t_L g1337 ( .A(n_1332), .B(n_1164), .C(n_1140), .D(n_1192), .Y(n_1337) );
AND2x4_ASAP7_75t_L g1338 ( .A(n_1335), .B(n_1193), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1336), .B(n_1334), .Y(n_1339) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_1337), .B(n_1223), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1338), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1340), .Y(n_1342) );
AOI21xp5_ASAP7_75t_L g1343 ( .A1(n_1341), .A2(n_1339), .B(n_1340), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1344 ( .A1(n_1343), .A2(n_1342), .B(n_1175), .Y(n_1344) );
OAI21xp5_ASAP7_75t_L g1345 ( .A1(n_1344), .A2(n_1111), .B(n_1110), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_1345), .A2(n_1181), .B1(n_1175), .B2(n_1182), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_1346), .A2(n_1192), .B1(n_1170), .B2(n_1261), .Y(n_1347) );
endmodule