module fake_jpeg_19450_n_311 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_56),
.Y(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_25),
.B1(n_34),
.B2(n_26),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_60),
.B1(n_36),
.B2(n_35),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_21),
.C(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_19),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_26),
.B1(n_29),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_57),
.B1(n_37),
.B2(n_54),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_59),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_44),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_77),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_52),
.B1(n_51),
.B2(n_55),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_90),
.B1(n_40),
.B2(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_21),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_31),
.B(n_11),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_73),
.B(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_93),
.Y(n_100)
);

AOI22x1_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_31),
.B1(n_40),
.B2(n_24),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_30),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_73),
.B(n_72),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_97),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_102),
.B(n_113),
.Y(n_130)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_107),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_71),
.B1(n_70),
.B2(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_116),
.B1(n_96),
.B2(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_69),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_73),
.B(n_67),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_118),
.B(n_66),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_117),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_78),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_120),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_71),
.B1(n_70),
.B2(n_62),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_90),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_78),
.B(n_71),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_78),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_90),
.A2(n_64),
.B1(n_62),
.B2(n_52),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_79),
.B1(n_86),
.B2(n_62),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_78),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_148),
.B(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_135),
.B1(n_110),
.B2(n_101),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_133),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_142),
.B1(n_117),
.B2(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_85),
.C(n_83),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_146),
.C(n_20),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_97),
.B1(n_78),
.B2(n_93),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_95),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_75),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_56),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_66),
.B1(n_64),
.B2(n_48),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_66),
.C(n_43),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_33),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_30),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_64),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_165),
.B1(n_150),
.B2(n_142),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_43),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_167),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_98),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_135),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_171),
.C(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_33),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_160),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_132),
.B(n_23),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_64),
.B1(n_21),
.B2(n_15),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_169),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_64),
.B1(n_13),
.B2(n_39),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_14),
.B(n_11),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_131),
.C(n_146),
.Y(n_171)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_149),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_130),
.B(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_14),
.B(n_11),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_64),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_151),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_193),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_164),
.C(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_189),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_145),
.B(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_191),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_195),
.B1(n_206),
.B2(n_163),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_40),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_13),
.B1(n_39),
.B2(n_44),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_205),
.B1(n_196),
.B2(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_40),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_203),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_13),
.B1(n_44),
.B2(n_22),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_223),
.C(n_18),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_160),
.C(n_164),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_191),
.B(n_189),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_166),
.C(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_216),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_179),
.C(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_32),
.C(n_28),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_222),
.B1(n_197),
.B2(n_199),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_155),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_167),
.B1(n_180),
.B2(n_16),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_167),
.C(n_43),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_195),
.B1(n_206),
.B2(n_14),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_40),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_231),
.B1(n_235),
.B2(n_247),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_220),
.B1(n_215),
.B2(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_189),
.B1(n_199),
.B2(n_194),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_244),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_210),
.B1(n_228),
.B2(n_226),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_23),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_246),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_245),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_23),
.C(n_9),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_17),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_24),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_13),
.B1(n_14),
.B2(n_22),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_221),
.C(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_253),
.C(n_255),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_218),
.B1(n_9),
.B2(n_10),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_254),
.B1(n_260),
.B2(n_0),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_27),
.C(n_20),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_22),
.B1(n_17),
.B2(n_7),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_20),
.C(n_18),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_20),
.C(n_18),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_232),
.C(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_8),
.B1(n_7),
.B2(n_22),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_234),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_257),
.B(n_258),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_269),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_8),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_271),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_12),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_8),
.B(n_1),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_0),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_275),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_18),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_2),
.C(n_3),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_18),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_0),
.B(n_2),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_254),
.C(n_1),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_280),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_4),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_3),
.C(n_4),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_3),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_4),
.B(n_5),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_295),
.B(n_297),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_287),
.A2(n_284),
.B(n_279),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_283),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_296),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_294),
.C(n_4),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_301),
.B(n_6),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_307),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_306),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_6),
.B(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_6),
.Y(n_311)
);


endmodule