module real_aes_11103_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_668;
wire n_237;
wire n_91;
AND2x2_ASAP7_75t_L g553 ( .A(n_0), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_0), .B(n_60), .Y(n_582) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_0), .Y(n_592) );
INVx1_ASAP7_75t_L g639 ( .A(n_0), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_1), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_2), .B(n_165), .Y(n_191) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_2), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_3), .B(n_126), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_4), .Y(n_561) );
INVx2_ASAP7_75t_L g518 ( .A(n_5), .Y(n_518) );
OR2x2_ASAP7_75t_L g680 ( .A(n_5), .B(n_533), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_6), .Y(n_632) );
INVx1_ASAP7_75t_L g552 ( .A(n_7), .Y(n_552) );
OR2x2_ASAP7_75t_L g581 ( .A(n_7), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g594 ( .A(n_7), .Y(n_594) );
BUFx2_ASAP7_75t_L g646 ( .A(n_7), .Y(n_646) );
INVx1_ASAP7_75t_L g602 ( .A(n_8), .Y(n_602) );
AOI221xp5_ASAP7_75t_SL g654 ( .A1(n_8), .A2(n_51), .B1(n_655), .B2(n_660), .C(n_665), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_9), .B(n_115), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_10), .B(n_107), .Y(n_257) );
INVx1_ASAP7_75t_L g566 ( .A(n_11), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_11), .A2(n_48), .B1(n_693), .B2(n_696), .C(n_699), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_12), .B(n_107), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_13), .B(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_14), .Y(n_555) );
INVx1_ASAP7_75t_L g615 ( .A(n_15), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_15), .A2(n_19), .B1(n_668), .B2(n_671), .Y(n_667) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_16), .Y(n_721) );
AOI22x1_ASAP7_75t_SL g724 ( .A1(n_17), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_17), .Y(n_727) );
AND2x2_ASAP7_75t_L g268 ( .A(n_18), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g596 ( .A(n_19), .Y(n_596) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_20), .Y(n_90) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_21), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_22), .B(n_185), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_23), .A2(n_538), .B1(n_722), .B2(n_741), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_23), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_24), .B(n_193), .Y(n_192) );
NAND2xp33_ASAP7_75t_L g255 ( .A(n_25), .B(n_193), .Y(n_255) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_27), .Y(n_114) );
INVx1_ASAP7_75t_L g517 ( .A(n_28), .Y(n_517) );
INVx1_ASAP7_75t_L g533 ( .A(n_28), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_29), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_30), .B(n_148), .Y(n_196) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_31), .A2(n_54), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_32), .A2(n_121), .B(n_273), .C(n_274), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_33), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_34), .B(n_119), .Y(n_142) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_35), .B(n_125), .Y(n_166) );
AND2x6_ASAP7_75t_L g84 ( .A(n_36), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_36), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_36), .B(n_510), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_37), .A2(n_45), .B1(n_574), .B2(n_583), .C(n_587), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_37), .A2(n_45), .B1(n_529), .B2(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_38), .B(n_118), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_39), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_40), .B(n_254), .Y(n_253) );
NAND2xp33_ASAP7_75t_L g209 ( .A(n_41), .B(n_125), .Y(n_209) );
INVx1_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_42), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_43), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_44), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_46), .B(n_125), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_47), .Y(n_629) );
INVx1_ASAP7_75t_L g542 ( .A(n_48), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_49), .Y(n_140) );
AND2x2_ASAP7_75t_L g276 ( .A(n_50), .B(n_185), .Y(n_276) );
INVx1_ASAP7_75t_L g610 ( .A(n_51), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_52), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g549 ( .A(n_53), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_55), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g177 ( .A(n_56), .B(n_93), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_57), .B(n_165), .Y(n_164) );
BUFx10_ASAP7_75t_L g527 ( .A(n_58), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_59), .B(n_92), .Y(n_251) );
INVx2_ASAP7_75t_L g554 ( .A(n_60), .Y(n_554) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_61), .B(n_115), .Y(n_183) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_62), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_63), .B(n_193), .Y(n_250) );
INVx1_ASAP7_75t_L g737 ( .A(n_64), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_65), .Y(n_275) );
INVx2_ASAP7_75t_L g110 ( .A(n_66), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_67), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_68), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_69), .B(n_152), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_70), .Y(n_204) );
INVx1_ASAP7_75t_L g267 ( .A(n_71), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_72), .Y(n_117) );
AND2x2_ASAP7_75t_L g132 ( .A(n_73), .B(n_107), .Y(n_132) );
INVx2_ASAP7_75t_L g550 ( .A(n_74), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_75), .B(n_185), .Y(n_184) );
BUFx3_ASAP7_75t_L g650 ( .A(n_76), .Y(n_650) );
INVx1_ASAP7_75t_L g675 ( .A(n_76), .Y(n_675) );
BUFx3_ASAP7_75t_L g525 ( .A(n_77), .Y(n_525) );
INVx1_ASAP7_75t_L g664 ( .A(n_77), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_95), .B(n_504), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_83), .A2(n_112), .B(n_122), .Y(n_111) );
INVx8_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
NOR2xp67_ASAP7_75t_L g262 ( .A(n_83), .B(n_263), .Y(n_262) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
BUFx2_ASAP7_75t_L g167 ( .A(n_84), .Y(n_167) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g753 ( .A1(n_87), .A2(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_88), .A2(n_266), .B(n_268), .Y(n_265) );
BUFx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_89), .Y(n_131) );
INVx3_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_89), .A2(n_164), .B(n_166), .Y(n_163) );
BUFx12f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx5_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_90), .A2(n_140), .B(n_141), .C(n_142), .Y(n_139) );
INVx5_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
INVx2_ASAP7_75t_L g179 ( .A(n_93), .Y(n_179) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_94), .Y(n_115) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_94), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_94), .Y(n_126) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g271 ( .A(n_94), .Y(n_271) );
INVx2_ASAP7_75t_SL g95 ( .A(n_96), .Y(n_95) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_403), .Y(n_96) );
NOR3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_321), .C(n_354), .Y(n_97) );
OAI211xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_133), .B(n_242), .C(n_306), .Y(n_98) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g328 ( .A(n_104), .B(n_260), .Y(n_328) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_105), .B(n_213), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_105), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g386 ( .A(n_105), .Y(n_386) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_132), .Y(n_105) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_106), .A2(n_111), .B(n_132), .Y(n_259) );
INVx3_ASAP7_75t_L g263 ( .A(n_106), .Y(n_263) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_L g137 ( .A(n_107), .Y(n_137) );
INVx3_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_107), .A2(n_175), .B(n_184), .Y(n_174) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_107), .A2(n_175), .B(n_184), .Y(n_219) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_107), .A2(n_175), .B(n_184), .Y(n_241) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g186 ( .A(n_109), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_120), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
INVx2_ASAP7_75t_L g165 ( .A(n_115), .Y(n_165) );
INVx2_ASAP7_75t_SL g254 ( .A(n_115), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx5_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
CKINVDCx6p67_ASAP7_75t_R g180 ( .A(n_121), .Y(n_180) );
OAI21xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B(n_131), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_124), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_124), .Y(n_738) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
INVx2_ASAP7_75t_L g193 ( .A(n_126), .Y(n_193) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_130), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_128), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_131), .A2(n_250), .B(n_251), .Y(n_249) );
AOI311xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_169), .A3(n_198), .B(n_211), .C(n_227), .Y(n_133) );
AND2x2_ASAP7_75t_L g283 ( .A(n_134), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g375 ( .A(n_134), .Y(n_375) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g337 ( .A(n_135), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_135), .B(n_172), .Y(n_489) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_154), .Y(n_135) );
AND2x2_ASAP7_75t_L g298 ( .A(n_136), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g308 ( .A(n_136), .B(n_225), .Y(n_308) );
INVx1_ASAP7_75t_L g319 ( .A(n_136), .Y(n_319) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_151), .Y(n_136) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_137), .A2(n_189), .B(n_197), .Y(n_188) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_137), .A2(n_202), .B(n_210), .Y(n_201) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_137), .A2(n_138), .B(n_151), .Y(n_218) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_189), .B(n_197), .Y(n_224) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_150), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_140), .A2(n_538), .B1(n_722), .B2(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_140), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_147), .C(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g751 ( .A(n_144), .Y(n_751) );
O2A1O1Ixp5_ASAP7_75t_L g194 ( .A1(n_145), .A2(n_149), .B(n_195), .C(n_196), .Y(n_194) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_L g203 ( .A1(n_149), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
OAI21x1_ASAP7_75t_L g175 ( .A1(n_150), .A2(n_176), .B(n_181), .Y(n_175) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_150), .A2(n_190), .B(n_194), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_150), .A2(n_203), .B(n_207), .Y(n_202) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_150), .A2(n_249), .B(n_252), .Y(n_248) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx2_ASAP7_75t_L g434 ( .A(n_154), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_168), .Y(n_154) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_155), .A2(n_157), .B(n_168), .Y(n_226) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_155), .A2(n_248), .B(n_257), .Y(n_247) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_163), .B(n_167), .Y(n_157) );
AOI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .Y(n_158) );
INVx1_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_162), .A2(n_182), .B(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g256 ( .A(n_162), .Y(n_256) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVxp67_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g449 ( .A(n_172), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_173), .B(n_187), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g340 ( .A(n_174), .B(n_299), .Y(n_340) );
AND2x2_ASAP7_75t_L g402 ( .A(n_174), .B(n_299), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_180), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_180), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_180), .A2(n_208), .B(n_209), .Y(n_207) );
BUFx5_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g284 ( .A(n_187), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_187), .B(n_217), .Y(n_452) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g479 ( .A(n_188), .B(n_294), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_193), .B(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x4_ASAP7_75t_L g367 ( .A(n_199), .B(n_368), .Y(n_367) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_199), .A2(n_394), .A3(n_397), .B1(n_398), .B2(n_400), .Y(n_393) );
AND2x4_ASAP7_75t_L g493 ( .A(n_199), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_200), .B(n_282), .Y(n_334) );
OR2x2_ASAP7_75t_L g345 ( .A(n_200), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_200), .B(n_281), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_200), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g416 ( .A(n_200), .B(n_246), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_200), .B(n_368), .Y(n_484) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g213 ( .A(n_201), .Y(n_213) );
AND2x2_ASAP7_75t_L g312 ( .A(n_201), .B(n_259), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .C(n_220), .Y(n_211) );
INVx1_ASAP7_75t_L g238 ( .A(n_212), .Y(n_238) );
AND2x2_ASAP7_75t_L g461 ( .A(n_212), .B(n_328), .Y(n_461) );
AND2x2_ASAP7_75t_L g469 ( .A(n_212), .B(n_430), .Y(n_469) );
BUFx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g325 ( .A(n_213), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g358 ( .A(n_213), .B(n_247), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
OAI211xp5_ASAP7_75t_SL g321 ( .A1(n_215), .A2(n_322), .B(n_329), .C(n_348), .Y(n_321) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g390 ( .A(n_217), .Y(n_390) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_217), .B(n_293), .Y(n_442) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_217), .B(n_377), .Y(n_474) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g232 ( .A(n_218), .Y(n_232) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_218), .Y(n_465) );
INVx2_ASAP7_75t_L g419 ( .A(n_219), .Y(n_419) );
INVx2_ASAP7_75t_L g430 ( .A(n_219), .Y(n_430) );
AND2x2_ASAP7_75t_L g498 ( .A(n_219), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g350 ( .A(n_221), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g347 ( .A(n_222), .B(n_231), .Y(n_347) );
AND2x2_ASAP7_75t_L g388 ( .A(n_222), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx2_ASAP7_75t_L g299 ( .A(n_223), .Y(n_299) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g236 ( .A(n_224), .B(n_225), .Y(n_236) );
INVx2_ASAP7_75t_L g294 ( .A(n_225), .Y(n_294) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_233), .C(n_237), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x4_ASAP7_75t_L g292 ( .A(n_231), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_233), .A2(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g427 ( .A(n_236), .B(n_240), .Y(n_427) );
NAND2xp33_ASAP7_75t_R g438 ( .A(n_236), .B(n_318), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g330 ( .A(n_240), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_SL g291 ( .A(n_241), .Y(n_291) );
INVx1_ASAP7_75t_L g351 ( .A(n_241), .Y(n_351) );
INVx1_ASAP7_75t_SL g396 ( .A(n_241), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_283), .B(n_285), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_277), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_258), .Y(n_244) );
OR2x2_ASAP7_75t_L g314 ( .A(n_245), .B(n_279), .Y(n_314) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g305 ( .A(n_247), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_247), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g326 ( .A(n_247), .Y(n_326) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_247), .Y(n_346) );
OR2x2_ASAP7_75t_L g369 ( .A(n_247), .B(n_259), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B(n_256), .Y(n_252) );
INVx2_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
AND2x2_ASAP7_75t_L g352 ( .A(n_258), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g423 ( .A(n_258), .Y(n_423) );
AND2x2_ASAP7_75t_L g443 ( .A(n_258), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g445 ( .A(n_258), .B(n_358), .Y(n_445) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g458 ( .A(n_259), .B(n_411), .Y(n_458) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
INVx1_ASAP7_75t_L g411 ( .A(n_260), .Y(n_411) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g282 ( .A(n_261), .Y(n_282) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_276), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_272), .Y(n_264) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI32xp33_ASAP7_75t_L g467 ( .A1(n_277), .A2(n_468), .A3(n_470), .B1(n_471), .B2(n_473), .Y(n_467) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g287 ( .A(n_279), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_282), .Y(n_344) );
OR2x2_ASAP7_75t_L g432 ( .A(n_284), .B(n_433), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_295), .B2(n_300), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_289), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g324 ( .A(n_290), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g362 ( .A(n_291), .B(n_299), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_291), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_292), .A2(n_383), .B1(n_388), .B2(n_391), .Y(n_382) );
AND2x2_ASAP7_75t_L g394 ( .A(n_292), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_294), .B(n_299), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_295), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g381 ( .A(n_298), .Y(n_381) );
INVx1_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_300), .A2(n_497), .B1(n_501), .B2(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g333 ( .A(n_304), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g379 ( .A(n_304), .B(n_374), .Y(n_379) );
INVx1_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B(n_313), .C(n_315), .Y(n_306) );
NAND2x1_ASAP7_75t_SL g360 ( .A(n_307), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_307), .B(n_339), .Y(n_407) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_308), .B(n_316), .C(n_320), .Y(n_315) );
OR2x6_ASAP7_75t_SL g418 ( .A(n_308), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_SL g331 ( .A(n_309), .Y(n_331) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g387 ( .A(n_310), .Y(n_387) );
AND2x2_ASAP7_75t_L g494 ( .A(n_310), .B(n_386), .Y(n_494) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_320), .A2(n_330), .B1(n_332), .B2(n_335), .C1(n_341), .C2(n_347), .Y(n_329) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
INVx1_ASAP7_75t_SL g399 ( .A(n_325), .Y(n_399) );
INVx1_ASAP7_75t_L g397 ( .A(n_327), .Y(n_397) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g398 ( .A(n_328), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g425 ( .A(n_328), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g436 ( .A(n_328), .B(n_358), .Y(n_436) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g392 ( .A(n_334), .Y(n_392) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g455 ( .A(n_336), .B(n_395), .Y(n_455) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_SL g412 ( .A(n_337), .B(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g466 ( .A(n_340), .Y(n_466) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_343), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g486 ( .A(n_343), .B(n_353), .Y(n_486) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
OR2x2_ASAP7_75t_L g453 ( .A(n_345), .B(n_423), .Y(n_453) );
AND2x2_ASAP7_75t_L g429 ( .A(n_347), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g451 ( .A(n_351), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g473 ( .A(n_351), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g502 ( .A(n_351), .B(n_503), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g354 ( .A(n_355), .B(n_370), .C(n_382), .D(n_393), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B1(n_363), .B2(n_365), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_409), .Y(n_408) );
NAND2xp67_ASAP7_75t_L g457 ( .A(n_358), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AO21x1_ASAP7_75t_L g477 ( .A1(n_361), .A2(n_442), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_362), .Y(n_364) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g391 ( .A(n_368), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_369), .Y(n_372) );
OR2x2_ASAP7_75t_L g462 ( .A(n_369), .B(n_410), .Y(n_462) );
AOI32xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .A3(n_376), .B1(n_378), .B2(n_380), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g501 ( .A(n_372), .Y(n_501) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_378), .A2(n_400), .B1(n_477), .B2(n_480), .C(n_482), .Y(n_476) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
BUFx2_ASAP7_75t_SL g472 ( .A(n_386), .Y(n_472) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g448 ( .A(n_390), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g495 ( .A(n_398), .B(n_478), .Y(n_495) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_475), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_428), .C(n_439), .D(n_454), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_412), .B2(n_413), .C(n_417), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_408), .A2(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g470 ( .A(n_409), .Y(n_470) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI31xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .A3(n_422), .B(n_424), .Y(n_417) );
NAND2xp33_ASAP7_75t_L g446 ( .A(n_418), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g478 ( .A(n_419), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_419), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
INVx1_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_430), .B(n_442), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B1(n_437), .B2(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_445), .B2(n_446), .C(n_450), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_442), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g492 ( .A(n_442), .Y(n_492) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_459), .B2(n_463), .C(n_467), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
INVx2_ASAP7_75t_L g503 ( .A(n_479), .Y(n_503) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_487), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_495), .C(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_536), .B1(n_740), .B2(n_742), .C(n_745), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .Y(n_508) );
OR2x4_ASAP7_75t_L g748 ( .A(n_509), .B(n_513), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_510), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g754 ( .A(n_510), .Y(n_754) );
INVx1_ASAP7_75t_L g744 ( .A(n_511), .Y(n_744) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AOI31xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_519), .A3(n_526), .B(n_528), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g666 ( .A(n_516), .Y(n_666) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x4_ASAP7_75t_L g710 ( .A(n_517), .B(n_534), .Y(n_710) );
INVx2_ASAP7_75t_L g534 ( .A(n_518), .Y(n_534) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g535 ( .A(n_522), .Y(n_535) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g648 ( .A(n_524), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g659 ( .A(n_525), .B(n_650), .Y(n_659) );
AND2x4_ASAP7_75t_L g674 ( .A(n_525), .B(n_675), .Y(n_674) );
INVx6_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
AND2x2_ASAP7_75t_L g647 ( .A(n_531), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g683 ( .A(n_531), .Y(n_683) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
XNOR2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_723), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_537) );
INVx1_ASAP7_75t_L g722 ( .A(n_538), .Y(n_722) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_640), .Y(n_538) );
NOR3xp33_ASAP7_75t_SL g539 ( .A(n_540), .B(n_573), .C(n_589), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_560), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B1(n_555), .B2(n_556), .Y(n_541) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_545), .B(n_551), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g619 ( .A(n_546), .Y(n_619) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_546), .Y(n_626) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x4_ASAP7_75t_L g558 ( .A(n_548), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g565 ( .A(n_549), .B(n_550), .Y(n_565) );
INVx1_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
INVx1_ASAP7_75t_L g579 ( .A(n_549), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_549), .B(n_550), .Y(n_601) );
INVx1_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_549), .B(n_570), .Y(n_614) );
INVx1_ASAP7_75t_L g559 ( .A(n_550), .Y(n_559) );
INVx2_ASAP7_75t_L g570 ( .A(n_550), .Y(n_570) );
INVx1_ASAP7_75t_L g608 ( .A(n_550), .Y(n_608) );
AND2x6_ASAP7_75t_L g556 ( .A(n_551), .B(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g562 ( .A(n_551), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_551), .B(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g636 ( .A(n_552), .Y(n_636) );
INVx1_ASAP7_75t_L g593 ( .A(n_554), .Y(n_593) );
INVx1_ASAP7_75t_L g638 ( .A(n_554), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_555), .A2(n_561), .B1(n_700), .B2(n_705), .C(n_708), .Y(n_699) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_557), .B(n_580), .Y(n_588) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_566), .B2(n_567), .Y(n_560) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g586 ( .A(n_570), .Y(n_586) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2x1_ASAP7_75t_SL g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_580), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g643 ( .A(n_581), .B(n_600), .Y(n_643) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI33xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .A3(n_609), .B1(n_620), .B2(n_628), .B3(n_633), .Y(n_589) );
OR2x6_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
BUFx2_ASAP7_75t_L g719 ( .A(n_594), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B1(n_602), .B2(n_603), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_597), .A2(n_629), .B1(n_630), .B2(n_632), .Y(n_628) );
BUFx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g631 ( .A(n_605), .Y(n_631) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_615), .B2(n_616), .Y(n_609) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx2_ASAP7_75t_L g622 ( .A(n_614), .Y(n_622) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B1(n_624), .B2(n_627), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_623), .A2(n_685), .B(n_687), .C(n_692), .Y(n_684) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_627), .A2(n_629), .B1(n_712), .B2(n_714), .Y(n_711) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_632), .A2(n_654), .B1(n_667), .B2(n_676), .C(n_681), .Y(n_653) );
CKINVDCx8_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
INVx5_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x6_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_651), .B(n_652), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx6_ASAP7_75t_L g670 ( .A(n_648), .Y(n_670) );
INVx1_ASAP7_75t_L g691 ( .A(n_649), .Y(n_691) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g663 ( .A(n_650), .B(n_664), .Y(n_663) );
AOI31xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_684), .A3(n_711), .B(n_717), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g681 ( .A(n_657), .B(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_659), .Y(n_678) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
BUFx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_663), .Y(n_686) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_663), .Y(n_695) );
INVx1_ASAP7_75t_L g704 ( .A(n_664), .Y(n_704) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g698 ( .A(n_674), .Y(n_698) );
INVx2_ASAP7_75t_L g716 ( .A(n_674), .Y(n_716) );
INVx1_ASAP7_75t_L g703 ( .A(n_675), .Y(n_703) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AND2x4_ASAP7_75t_L g685 ( .A(n_679), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g713 ( .A(n_680), .B(n_707), .Y(n_713) );
OR2x2_ASAP7_75t_L g715 ( .A(n_680), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g688 ( .A(n_683), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
BUFx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
BUFx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
OR2x2_ASAP7_75t_L g707 ( .A(n_703), .B(n_704), .Y(n_707) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx6_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx4_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_739), .Y(n_728) );
CKINVDCx14_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g739 ( .A(n_731), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx14_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B1(n_751), .B2(n_752), .Y(n_745) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx8_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
endmodule