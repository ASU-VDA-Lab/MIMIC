module real_aes_2877_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_774, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_773, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_775, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_774;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_773;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_775;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_461;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_639;
wire n_587;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
wire n_429;
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_0), .A2(n_224), .B1(n_451), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_1), .A2(n_221), .B1(n_461), .B2(n_473), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_2), .A2(n_239), .B1(n_516), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_3), .A2(n_130), .B1(n_332), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_4), .A2(n_107), .B1(n_463), .B2(n_540), .Y(n_539) );
AOI222xp33_ASAP7_75t_L g569 ( .A1(n_5), .A2(n_99), .B1(n_269), .B2(n_388), .C1(n_570), .C2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_6), .A2(n_160), .B1(n_389), .B2(n_598), .Y(n_597) );
OA22x2_ASAP7_75t_L g376 ( .A1(n_7), .A2(n_377), .B1(n_378), .B2(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_7), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_8), .A2(n_88), .B1(n_418), .B2(n_420), .Y(n_417) );
OA22x2_ASAP7_75t_L g749 ( .A1(n_9), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_9), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_10), .A2(n_75), .B1(n_319), .B2(n_324), .Y(n_318) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_11), .A2(n_196), .B1(n_296), .B2(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g727 ( .A(n_11), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_12), .A2(n_182), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_13), .A2(n_41), .B1(n_401), .B2(n_490), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_14), .A2(n_177), .B1(n_404), .B2(n_405), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_15), .A2(n_90), .B1(n_344), .B2(n_412), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_16), .A2(n_36), .B1(n_331), .B2(n_336), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_17), .B(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_18), .A2(n_199), .B1(n_359), .B2(n_487), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_19), .A2(n_91), .B1(n_693), .B2(n_702), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_20), .A2(n_21), .B1(n_367), .B2(n_369), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_22), .A2(n_82), .B1(n_337), .B2(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_23), .A2(n_136), .B1(n_566), .B2(n_567), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_24), .A2(n_195), .B1(n_385), .B2(n_574), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_25), .A2(n_120), .B1(n_352), .B2(n_540), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_26), .A2(n_134), .B1(n_401), .B2(n_589), .Y(n_588) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_27), .A2(n_63), .B1(n_229), .B2(n_290), .C1(n_314), .C2(n_451), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_28), .A2(n_47), .B1(n_382), .B2(n_383), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_29), .A2(n_219), .B1(n_319), .B2(n_324), .Y(n_738) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_30), .A2(n_77), .B1(n_296), .B2(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_30), .B(n_726), .Y(n_725) );
OA22x2_ASAP7_75t_L g509 ( .A1(n_31), .A2(n_510), .B1(n_524), .B2(n_525), .Y(n_509) );
INVx1_ASAP7_75t_L g524 ( .A(n_31), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_32), .A2(n_203), .B1(n_428), .B2(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_33), .A2(n_172), .B1(n_469), .B2(n_628), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_34), .A2(n_43), .B1(n_359), .B2(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g666 ( .A(n_35), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_37), .A2(n_202), .B1(n_466), .B2(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_38), .B(n_656), .Y(n_655) );
OA22x2_ASAP7_75t_L g407 ( .A1(n_39), .A2(n_408), .B1(n_409), .B2(n_436), .Y(n_407) );
INVx1_ASAP7_75t_L g436 ( .A(n_39), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_40), .A2(n_48), .B1(n_396), .B2(n_564), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_42), .A2(n_261), .B1(n_355), .B2(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_44), .B(n_446), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_45), .A2(n_133), .B1(n_344), .B2(n_348), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_46), .A2(n_234), .B1(n_388), .B2(n_570), .Y(n_607) );
INVx1_ASAP7_75t_L g691 ( .A(n_49), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_49), .A2(n_50), .B(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_49), .A2(n_706), .B1(n_714), .B2(n_775), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_50), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_51), .A2(n_235), .B1(n_385), .B2(n_574), .Y(n_611) );
AOI222xp33_ASAP7_75t_SL g710 ( .A1(n_52), .A2(n_129), .B1(n_180), .B2(n_514), .C1(n_711), .C2(n_712), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_53), .A2(n_94), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_54), .A2(n_210), .B1(n_332), .B2(n_426), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_55), .A2(n_58), .B1(n_320), .B2(n_516), .Y(n_515) );
AOI22x1_ASAP7_75t_L g480 ( .A1(n_56), .A2(n_481), .B1(n_504), .B2(n_505), .Y(n_480) );
CKINVDCx14_ASAP7_75t_R g505 ( .A(n_56), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_57), .A2(n_211), .B1(n_454), .B2(n_537), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_59), .A2(n_265), .B1(n_404), .B2(n_405), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_60), .A2(n_115), .B1(n_516), .B2(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_61), .A2(n_213), .B1(n_429), .B2(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_62), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_64), .A2(n_243), .B1(n_364), .B2(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_65), .A2(n_207), .B1(n_454), .B2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_66), .A2(n_268), .B1(n_522), .B2(n_636), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_67), .A2(n_188), .B1(n_471), .B2(n_473), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_68), .A2(n_76), .B1(n_431), .B2(n_433), .Y(n_430) );
OAI22x1_ASAP7_75t_SL g528 ( .A1(n_69), .A2(n_529), .B1(n_545), .B2(n_546), .Y(n_528) );
INVx1_ASAP7_75t_L g545 ( .A(n_69), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_70), .A2(n_81), .B1(n_319), .B2(n_324), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_71), .A2(n_109), .B1(n_471), .B2(n_473), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_72), .A2(n_118), .B1(n_398), .B2(n_399), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_73), .A2(n_217), .B1(n_367), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_74), .A2(n_205), .B1(n_449), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_78), .A2(n_121), .B1(n_451), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_79), .A2(n_237), .B1(n_463), .B2(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_80), .A2(n_104), .B1(n_422), .B2(n_423), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_83), .A2(n_191), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx3_ASAP7_75t_L g296 ( .A(n_84), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_85), .A2(n_169), .B1(n_382), .B2(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_86), .A2(n_154), .B1(n_348), .B2(n_414), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_87), .A2(n_193), .B1(n_352), .B2(n_589), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_89), .A2(n_267), .B1(n_352), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_92), .A2(n_95), .B1(n_344), .B2(n_346), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_93), .A2(n_254), .B1(n_492), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_96), .A2(n_170), .B1(n_398), .B2(n_399), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_97), .A2(n_122), .B1(n_371), .B2(n_485), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_98), .B(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_100), .A2(n_209), .B1(n_688), .B2(n_689), .Y(n_687) );
AO22x2_ASAP7_75t_L g441 ( .A1(n_101), .A2(n_442), .B1(n_443), .B2(n_474), .Y(n_441) );
INVx1_ASAP7_75t_L g474 ( .A(n_101), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_102), .A2(n_197), .B1(n_360), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_103), .A2(n_135), .B1(n_362), .B2(n_466), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_105), .A2(n_146), .B1(n_388), .B2(n_389), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_106), .A2(n_166), .B1(n_454), .B2(n_533), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_108), .A2(n_141), .B1(n_451), .B2(n_514), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_110), .A2(n_230), .B1(n_351), .B2(n_355), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_111), .A2(n_147), .B1(n_471), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_SL g297 ( .A(n_112), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_112), .B(n_144), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_113), .A2(n_216), .B1(n_370), .B2(n_636), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g734 ( .A1(n_114), .A2(n_139), .B1(n_253), .B2(n_449), .C1(n_456), .C2(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g278 ( .A(n_116), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_117), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_119), .A2(n_179), .B1(n_399), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_123), .A2(n_257), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_124), .A2(n_215), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_125), .A2(n_164), .B1(n_332), .B2(n_337), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_126), .A2(n_231), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_127), .A2(n_263), .B1(n_455), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_128), .A2(n_176), .B1(n_402), .B2(n_461), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_131), .A2(n_236), .B1(n_371), .B2(n_418), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_132), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_137), .A2(n_238), .B1(n_370), .B2(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_138), .A2(n_198), .B1(n_382), .B2(n_383), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_140), .A2(n_228), .B1(n_401), .B2(n_420), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_142), .A2(n_178), .B1(n_364), .B2(n_467), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_143), .A2(n_171), .B1(n_412), .B2(n_414), .Y(n_679) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_144), .A2(n_204), .B1(n_296), .B2(n_300), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_145), .A2(n_225), .B1(n_320), .B2(n_516), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_148), .A2(n_731), .B1(n_732), .B2(n_745), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_148), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_149), .A2(n_212), .B1(n_429), .B2(n_763), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_150), .A2(n_186), .B1(n_364), .B2(n_628), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_151), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_152), .A2(n_190), .B1(n_320), .B2(n_516), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_153), .Y(n_654) );
OA22x2_ASAP7_75t_L g284 ( .A1(n_155), .A2(n_285), .B1(n_286), .B2(n_372), .Y(n_284) );
INVx1_ASAP7_75t_L g372 ( .A(n_155), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_156), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_157), .A2(n_220), .B1(n_537), .B2(n_684), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_158), .A2(n_187), .B1(n_344), .B2(n_412), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_159), .A2(n_168), .B1(n_371), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_161), .A2(n_256), .B1(n_415), .B2(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_162), .B(n_735), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_163), .A2(n_262), .B1(n_319), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g298 ( .A(n_165), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_167), .B(n_391), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_173), .A2(n_227), .B1(n_309), .B2(n_503), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_174), .B(n_571), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_175), .A2(n_242), .B1(n_466), .B2(n_542), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_181), .A2(n_183), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_184), .A2(n_245), .B1(n_395), .B2(n_396), .Y(n_614) );
XNOR2x1_ASAP7_75t_L g620 ( .A(n_185), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_189), .B(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_192), .A2(n_201), .B1(n_309), .B2(n_314), .Y(n_308) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_194), .A2(n_206), .B1(n_467), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_200), .A2(n_246), .B1(n_364), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_208), .A2(n_260), .B1(n_463), .B2(n_464), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_214), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g723 ( .A(n_214), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_218), .A2(n_258), .B1(n_684), .B2(n_686), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_222), .A2(n_252), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
AND2x2_ASAP7_75t_R g747 ( .A(n_223), .B(n_723), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_226), .B(n_290), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_232), .B(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_233), .A2(n_244), .B1(n_337), .B2(n_455), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_240), .B(n_277), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_241), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_247), .B(n_516), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_248), .A2(n_266), .B1(n_343), .B2(n_346), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_249), .A2(n_264), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI211x1_ASAP7_75t_SL g270 ( .A1(n_250), .A2(n_271), .B(n_279), .C(n_729), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_251), .A2(n_255), .B1(n_332), .B2(n_426), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_259), .B(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g771 ( .A(n_274), .B(n_276), .Y(n_771) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_275), .B(n_723), .Y(n_722) );
AOI221xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_550), .B1(n_718), .B2(n_719), .C(n_720), .Y(n_279) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_280), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_476), .B1(n_477), .B2(n_549), .Y(n_280) );
INVx1_ASAP7_75t_L g549 ( .A(n_281), .Y(n_549) );
AOI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_440), .B1(n_441), .B2(n_475), .Y(n_281) );
INVx1_ASAP7_75t_L g475 ( .A(n_282), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_373), .B1(n_438), .B2(n_439), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g439 ( .A(n_284), .Y(n_439) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_341), .Y(n_286) );
NAND4xp25_ASAP7_75t_SL g287 ( .A(n_288), .B(n_308), .C(n_318), .D(n_330), .Y(n_287) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_SL g391 ( .A(n_291), .Y(n_391) );
INVx4_ASAP7_75t_SL g435 ( .A(n_291), .Y(n_435) );
INVx4_ASAP7_75t_SL g447 ( .A(n_291), .Y(n_447) );
BUFx2_ASAP7_75t_L g495 ( .A(n_291), .Y(n_495) );
INVx3_ASAP7_75t_L g711 ( .A(n_291), .Y(n_711) );
INVx6_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_301), .Y(n_292) );
AND2x4_ASAP7_75t_L g316 ( .A(n_293), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g338 ( .A(n_293), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g383 ( .A(n_293), .B(n_339), .Y(n_383) );
AND2x2_ASAP7_75t_L g389 ( .A(n_293), .B(n_317), .Y(n_389) );
AND2x2_ASAP7_75t_L g570 ( .A(n_293), .B(n_317), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_293), .B(n_301), .Y(n_571) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
INVx2_ASAP7_75t_L g313 ( .A(n_294), .Y(n_313) );
AND2x2_ASAP7_75t_L g322 ( .A(n_294), .B(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_294), .Y(n_329) );
OAI22x1_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B1(n_297), .B2(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
INVx2_ASAP7_75t_L g304 ( .A(n_296), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
AND2x2_ASAP7_75t_L g312 ( .A(n_299), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
BUFx2_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
AND2x4_ASAP7_75t_L g345 ( .A(n_301), .B(n_322), .Y(n_345) );
AND2x4_ASAP7_75t_L g354 ( .A(n_301), .B(n_349), .Y(n_354) );
AND2x2_ASAP7_75t_L g368 ( .A(n_301), .B(n_312), .Y(n_368) );
AND2x6_ASAP7_75t_L g398 ( .A(n_301), .B(n_312), .Y(n_398) );
AND2x2_ASAP7_75t_L g404 ( .A(n_301), .B(n_322), .Y(n_404) );
AND2x2_ASAP7_75t_L g567 ( .A(n_301), .B(n_349), .Y(n_567) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g311 ( .A(n_303), .B(n_305), .Y(n_311) );
AND2x2_ASAP7_75t_L g328 ( .A(n_303), .B(n_306), .Y(n_328) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
INVxp67_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g428 ( .A(n_310), .Y(n_428) );
BUFx3_ASAP7_75t_L g451 ( .A(n_310), .Y(n_451) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_310), .Y(n_712) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g321 ( .A(n_311), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g371 ( .A(n_311), .B(n_349), .Y(n_371) );
AND2x4_ASAP7_75t_L g385 ( .A(n_311), .B(n_322), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_311), .B(n_312), .Y(n_388) );
AND2x2_ASAP7_75t_L g566 ( .A(n_311), .B(n_349), .Y(n_566) );
AND2x2_ASAP7_75t_L g598 ( .A(n_311), .B(n_312), .Y(n_598) );
AND2x2_ASAP7_75t_L g361 ( .A(n_312), .B(n_334), .Y(n_361) );
AND2x2_ASAP7_75t_L g395 ( .A(n_312), .B(n_334), .Y(n_395) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_312), .B(n_334), .Y(n_564) );
AND2x4_ASAP7_75t_L g349 ( .A(n_313), .B(n_323), .Y(n_349) );
INVx2_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g429 ( .A(n_315), .Y(n_429) );
INVx2_ASAP7_75t_L g503 ( .A(n_315), .Y(n_503) );
INVx2_ASAP7_75t_L g514 ( .A(n_315), .Y(n_514) );
INVx2_ASAP7_75t_L g533 ( .A(n_315), .Y(n_533) );
INVx6_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g432 ( .A(n_321), .Y(n_432) );
BUFx3_ASAP7_75t_L g498 ( .A(n_321), .Y(n_498) );
BUFx5_ASAP7_75t_L g674 ( .A(n_321), .Y(n_674) );
AND2x2_ASAP7_75t_L g333 ( .A(n_322), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g382 ( .A(n_322), .B(n_334), .Y(n_382) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g433 ( .A(n_326), .Y(n_433) );
INVx3_ASAP7_75t_L g499 ( .A(n_326), .Y(n_499) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx12f_ASAP7_75t_L g516 ( .A(n_327), .Y(n_516) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x4_ASAP7_75t_L g348 ( .A(n_328), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g364 ( .A(n_328), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_SL g386 ( .A(n_328), .B(n_329), .Y(n_386) );
AND2x4_ASAP7_75t_L g396 ( .A(n_328), .B(n_365), .Y(n_396) );
AND2x4_ASAP7_75t_L g405 ( .A(n_328), .B(n_349), .Y(n_405) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_328), .B(n_329), .Y(n_574) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_333), .Y(n_455) );
INVx3_ASAP7_75t_L g672 ( .A(n_333), .Y(n_672) );
AND2x4_ASAP7_75t_L g357 ( .A(n_334), .B(n_349), .Y(n_357) );
AND2x6_ASAP7_75t_L g399 ( .A(n_334), .B(n_349), .Y(n_399) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_335), .Y(n_340) );
BUFx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g426 ( .A(n_338), .Y(n_426) );
INVx2_ASAP7_75t_L g458 ( .A(n_338), .Y(n_458) );
BUFx4f_ASAP7_75t_L g625 ( .A(n_338), .Y(n_625) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_342), .B(n_350), .C(n_358), .D(n_366), .Y(n_341) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g414 ( .A(n_345), .Y(n_414) );
INVx6_ASAP7_75t_L g472 ( .A(n_345), .Y(n_472) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g412 ( .A(n_348), .Y(n_412) );
BUFx3_ASAP7_75t_L g490 ( .A(n_348), .Y(n_490) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
INVx2_ASAP7_75t_L g461 ( .A(n_353), .Y(n_461) );
INVx2_ASAP7_75t_SL g703 ( .A(n_353), .Y(n_703) );
INVx3_ASAP7_75t_SL g742 ( .A(n_353), .Y(n_742) );
INVx8_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g420 ( .A(n_356), .Y(n_420) );
INVx2_ASAP7_75t_L g464 ( .A(n_356), .Y(n_464) );
INVx2_ASAP7_75t_L g522 ( .A(n_356), .Y(n_522) );
INVx2_ASAP7_75t_L g540 ( .A(n_356), .Y(n_540) );
INVx2_ASAP7_75t_L g688 ( .A(n_356), .Y(n_688) );
INVx2_ASAP7_75t_SL g759 ( .A(n_356), .Y(n_759) );
INVx8_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
INVx2_ASAP7_75t_L g468 ( .A(n_361), .Y(n_468) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g423 ( .A(n_363), .Y(n_423) );
INVx2_ASAP7_75t_L g469 ( .A(n_363), .Y(n_469) );
INVx2_ASAP7_75t_L g542 ( .A(n_363), .Y(n_542) );
INVx5_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g487 ( .A(n_364), .Y(n_487) );
BUFx2_ASAP7_75t_L g582 ( .A(n_364), .Y(n_582) );
BUFx3_ASAP7_75t_L g463 ( .A(n_367), .Y(n_463) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g419 ( .A(n_368), .Y(n_419) );
BUFx2_ASAP7_75t_L g636 ( .A(n_368), .Y(n_636) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx2_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
BUFx3_ASAP7_75t_L g694 ( .A(n_371), .Y(n_694) );
INVx1_ASAP7_75t_L g438 ( .A(n_373), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_406), .B2(n_437), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_380), .B(n_392), .Y(n_379) );
NAND4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .C(n_387), .D(n_390), .Y(n_380) );
INVx2_ASAP7_75t_L g736 ( .A(n_391), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_400), .C(n_403), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g585 ( .A(n_398), .Y(n_585) );
BUFx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_424), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .C(n_417), .D(n_421), .Y(n_410) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g589 ( .A(n_416), .Y(n_589) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g492 ( .A(n_419), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .C(n_430), .D(n_434), .Y(n_424) );
BUFx6f_ASAP7_75t_SL g686 ( .A(n_426), .Y(n_686) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g656 ( .A(n_432), .Y(n_656) );
INVx1_ASAP7_75t_L g698 ( .A(n_432), .Y(n_698) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_459), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_448), .C(n_452), .D(n_453), .Y(n_444) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g537 ( .A(n_458), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .C(n_465), .D(n_470), .Y(n_459) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g628 ( .A(n_468), .Y(n_628) );
INVx2_ASAP7_75t_L g709 ( .A(n_468), .Y(n_709) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g485 ( .A(n_472), .Y(n_485) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OA22x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_506), .B1(n_547), .B2(n_548), .Y(n_477) );
INVx1_ASAP7_75t_L g547 ( .A(n_478), .Y(n_547) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g504 ( .A(n_481), .Y(n_504) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g494 ( .A1(n_495), .A2(n_496), .B(n_497), .Y(n_494) );
BUFx6f_ASAP7_75t_SL g767 ( .A(n_498), .Y(n_767) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_499), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g548 ( .A(n_506), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_509), .B1(n_526), .B2(n_527), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g525 ( .A(n_510), .Y(n_525) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .C(n_515), .D(n_517), .Y(n_511) );
BUFx3_ASAP7_75t_L g766 ( .A(n_516), .Y(n_766) );
NAND4xp25_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .C(n_521), .D(n_523), .Y(n_518) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g546 ( .A(n_529), .Y(n_546) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_538), .Y(n_529) );
NAND4xp25_ASAP7_75t_SL g530 ( .A(n_531), .B(n_532), .C(n_534), .D(n_536), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .C(n_543), .D(n_544), .Y(n_538) );
INVx2_ASAP7_75t_SL g718 ( .A(n_550), .Y(n_718) );
XNOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_662), .Y(n_550) );
BUFx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_639), .B2(n_640), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
XNOR2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_601), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_576), .B(n_599), .Y(n_556) );
OA22x2_ASAP7_75t_L g641 ( .A1(n_557), .A2(n_558), .B1(n_642), .B2(n_643), .Y(n_641) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g600 ( .A(n_558), .Y(n_600) );
XNOR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_575), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_568), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .D(n_565), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .C(n_573), .Y(n_568) );
INVx2_ASAP7_75t_SL g592 ( .A(n_571), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_576), .B(n_600), .Y(n_599) );
XNOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_579), .B(n_590), .Y(n_578) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_586), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_595), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B(n_594), .Y(n_591) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_592), .A2(n_654), .B(n_655), .C(n_657), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AO22x2_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_620), .B1(n_637), .B2(n_638), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
XOR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_619), .Y(n_603) );
XOR2x2_ASAP7_75t_L g638 ( .A(n_604), .B(n_619), .Y(n_638) );
NAND2x1_ASAP7_75t_SL g604 ( .A(n_605), .B(n_612), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx2_ASAP7_75t_L g637 ( .A(n_620), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_630), .D(n_633), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g690 ( .A(n_636), .Y(n_690) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_661), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_652), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_658), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_664), .B1(n_680), .B2(n_717), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
XNOR2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_675), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .C(n_673), .Y(n_668) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g685 ( .A(n_672), .Y(n_685) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .C(n_678), .D(n_679), .Y(n_675) );
INVx2_ASAP7_75t_SL g717 ( .A(n_680), .Y(n_717) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_699), .Y(n_680) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_691), .B1(n_692), .B2(n_695), .C1(n_773), .C2(n_774), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_682), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_687), .Y(n_682) );
BUFx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_692), .B(n_695), .C(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_SL g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B(n_713), .Y(n_699) );
INVx1_ASAP7_75t_L g716 ( .A(n_702), .Y(n_716) );
BUFx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx3_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_722), .B(n_725), .Y(n_770) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_746), .B1(n_748), .B2(n_750), .C1(n_768), .C2(n_771), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_739), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .C(n_738), .Y(n_733) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .C(n_743), .D(n_744), .Y(n_739) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR3x1_ASAP7_75t_SL g752 ( .A(n_753), .B(n_756), .C(n_760), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NAND4xp25_ASAP7_75t_SL g760 ( .A(n_761), .B(n_762), .C(n_764), .D(n_765), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
CKINVDCx6p67_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
endmodule