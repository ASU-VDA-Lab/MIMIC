module fake_ariane_1988_n_887 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_887);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_887;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_712;
wire n_484;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_92),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_46),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_129),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_108),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_62),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_76),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_59),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_106),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_135),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

BUFx2_ASAP7_75t_SL g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_24),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_28),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_42),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_55),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_58),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_186),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_51),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_27),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_117),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_73),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_90),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_71),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_26),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_193),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_153),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_181),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_25),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_152),
.Y(n_257)
);

INVxp33_ASAP7_75t_R g258 ( 
.A(n_78),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_127),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_54),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_178),
.B(n_47),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_75),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_190),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_188),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_70),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_125),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_192),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_88),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_80),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_97),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_48),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_139),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_187),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_0),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_0),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_209),
.B(n_1),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_216),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_216),
.B(n_2),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_211),
.B(n_2),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_213),
.B(n_215),
.Y(n_292)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_203),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_3),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_203),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_202),
.B(n_30),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_3),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_225),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

BUFx8_ASAP7_75t_SL g303 ( 
.A(n_204),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_204),
.B(n_31),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_230),
.B(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_231),
.B(n_5),
.Y(n_307)
);

BUFx8_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_237),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_201),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_241),
.B(n_5),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_203),
.B(n_6),
.Y(n_315)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_199),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_251),
.B(n_6),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_202),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_240),
.B(n_7),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_262),
.B(n_8),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_8),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_9),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_199),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_243),
.B(n_9),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_205),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_244),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_205),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_200),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_207),
.B(n_10),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_206),
.B1(n_229),
.B2(n_279),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_206),
.B1(n_229),
.B2(n_256),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_293),
.B(n_207),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_290),
.A2(n_249),
.B1(n_273),
.B2(n_233),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_290),
.B(n_233),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_223),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_329),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_247),
.Y(n_345)
);

NAND3x1_ASAP7_75t_L g346 ( 
.A(n_281),
.B(n_261),
.C(n_10),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_247),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_270),
.B1(n_275),
.B2(n_272),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_287),
.A2(n_270),
.B1(n_277),
.B2(n_269),
.Y(n_349)
);

AND2x2_ASAP7_75t_SL g350 ( 
.A(n_281),
.B(n_208),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_282),
.A2(n_268),
.B1(n_266),
.B2(n_265),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_282),
.A2(n_263),
.B1(n_260),
.B2(n_259),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_286),
.B(n_210),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_212),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_214),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_312),
.A2(n_257),
.B1(n_254),
.B2(n_253),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_291),
.A2(n_252),
.B1(n_248),
.B2(n_236),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_307),
.A2(n_235),
.B1(n_234),
.B2(n_232),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_226),
.B1(n_224),
.B2(n_222),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_313),
.A2(n_218),
.B1(n_217),
.B2(n_13),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_323),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_364)
);

AO22x2_ASAP7_75t_L g365 ( 
.A1(n_315),
.A2(n_322),
.B1(n_328),
.B2(n_317),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_33),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_316),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_367)
);

OA22x2_ASAP7_75t_L g368 ( 
.A1(n_301),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g371 ( 
.A1(n_304),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_316),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_293),
.B(n_19),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_293),
.B(n_20),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_34),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_304),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_288),
.B(n_27),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_324),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_310),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_310),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_R g383 ( 
.A1(n_306),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_303),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_288),
.B(n_49),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_284),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_306),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_L g389 ( 
.A1(n_288),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_288),
.B(n_197),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_341),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_288),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_336),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_344),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_350),
.B(n_302),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_338),
.A2(n_325),
.B(n_330),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_334),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_351),
.B(n_334),
.Y(n_404)
);

OR2x6_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_365),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_302),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_302),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_376),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_369),
.Y(n_411)
);

BUFx6f_ASAP7_75t_SL g412 ( 
.A(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_337),
.B(n_300),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_302),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_388),
.B(n_308),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

XNOR2x2_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_372),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_358),
.B(n_302),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_357),
.B(n_285),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_339),
.B(n_315),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_352),
.B(n_300),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_374),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_308),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_349),
.B(n_285),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_373),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_366),
.A2(n_292),
.B(n_298),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_364),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_375),
.B(n_311),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

XOR2x2_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_308),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

NAND2x1p5_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_315),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_354),
.B(n_292),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_342),
.B(n_334),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_347),
.B(n_311),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_341),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_341),
.Y(n_458)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_347),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_350),
.B(n_303),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_342),
.B(n_289),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_350),
.B(n_335),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_397),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_396),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_405),
.B(n_317),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_397),
.B(n_289),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_391),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_460),
.B(n_319),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_425),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_319),
.B(n_335),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_404),
.B(n_289),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_320),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_320),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_318),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_402),
.B(n_318),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_404),
.B(n_331),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_414),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_436),
.A2(n_298),
.B(n_331),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_412),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_309),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_402),
.B(n_280),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_327),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_412),
.Y(n_496)
);

CKINVDCx11_ASAP7_75t_R g497 ( 
.A(n_393),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_428),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_395),
.B(n_445),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_417),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_395),
.B(n_280),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_434),
.B(n_298),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_333),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_392),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_455),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_449),
.B(n_333),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_450),
.B(n_333),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_457),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_283),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_454),
.B(n_283),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_298),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_447),
.B(n_333),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_451),
.A2(n_298),
.B(n_296),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_424),
.B(n_283),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_429),
.B(n_284),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_409),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_392),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_461),
.B(n_283),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_409),
.B(n_296),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_439),
.B(n_321),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_446),
.B(n_321),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_446),
.B(n_321),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_452),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_493),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_406),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_495),
.B(n_516),
.Y(n_539)
);

BUFx6f_ASAP7_75t_SL g540 ( 
.A(n_465),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_401),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_522),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_401),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_522),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_532),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_469),
.B(n_422),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_463),
.B(n_442),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_487),
.B(n_394),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_476),
.B(n_427),
.Y(n_551)
);

INVx6_ASAP7_75t_SL g552 ( 
.A(n_476),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_463),
.B(n_442),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_532),
.B(n_394),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_476),
.B(n_427),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_465),
.B(n_411),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_465),
.B(n_411),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_472),
.B(n_393),
.Y(n_560)
);

BUFx4f_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_467),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_509),
.B(n_451),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_489),
.B(n_416),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_498),
.B(n_475),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_524),
.B(n_430),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_464),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_498),
.B(n_448),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_478),
.B(n_419),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_492),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_493),
.B(n_321),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_485),
.B(n_321),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_523),
.B(n_63),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_468),
.B(n_64),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_510),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_508),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_523),
.B(n_65),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_479),
.B(n_66),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_497),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_485),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_496),
.B(n_67),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_506),
.B(n_196),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_509),
.B(n_68),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_69),
.Y(n_593)
);

BUFx4_ASAP7_75t_SL g594 ( 
.A(n_588),
.Y(n_594)
);

INVx8_ASAP7_75t_L g595 ( 
.A(n_540),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_548),
.A2(n_530),
.B1(n_506),
.B2(n_519),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_537),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_579),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_535),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_561),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_565),
.B(n_486),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_556),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_541),
.Y(n_604)
);

INVx5_ASAP7_75t_SL g605 ( 
.A(n_535),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_568),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_535),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_543),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_540),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_551),
.B(n_479),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_543),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_563),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_541),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_562),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

BUFx2_ASAP7_75t_SL g618 ( 
.A(n_582),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_547),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_590),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_544),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_578),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_569),
.Y(n_625)
);

BUFx4_ASAP7_75t_SL g626 ( 
.A(n_590),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_549),
.B(n_479),
.Y(n_627)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_569),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_591),
.Y(n_629)
);

BUFx2_ASAP7_75t_SL g630 ( 
.A(n_582),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_553),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_574),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_566),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_574),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_567),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_554),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_617),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_618),
.A2(n_630),
.B1(n_536),
.B2(n_545),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_594),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_624),
.A2(n_577),
.B1(n_573),
.B2(n_539),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_627),
.A2(n_539),
.B1(n_470),
.B2(n_564),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_598),
.Y(n_644)
);

CKINVDCx11_ASAP7_75t_R g645 ( 
.A(n_614),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_627),
.A2(n_470),
.B1(n_564),
.B2(n_538),
.Y(n_646)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_614),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_638),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_603),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_613),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_595),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_610),
.Y(n_652)
);

BUFx2_ASAP7_75t_SL g653 ( 
.A(n_616),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_636),
.A2(n_545),
.B1(n_558),
.B2(n_559),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_623),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_SL g657 ( 
.A1(n_620),
.A2(n_551),
.B1(n_557),
.B2(n_583),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_595),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

BUFx2_ASAP7_75t_SL g660 ( 
.A(n_616),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_620),
.A2(n_558),
.B1(n_559),
.B2(n_550),
.Y(n_662)
);

BUFx8_ASAP7_75t_L g663 ( 
.A(n_631),
.Y(n_663)
);

BUFx8_ASAP7_75t_L g664 ( 
.A(n_626),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_SL g665 ( 
.A1(n_629),
.A2(n_583),
.B1(n_557),
.B2(n_551),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_619),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_632),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_596),
.A2(n_550),
.B1(n_571),
.B2(n_542),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_622),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_599),
.Y(n_671)
);

CKINVDCx6p67_ASAP7_75t_R g672 ( 
.A(n_595),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

INVx3_ASAP7_75t_SL g674 ( 
.A(n_599),
.Y(n_674)
);

INVx6_ASAP7_75t_L g675 ( 
.A(n_595),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_628),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_638),
.Y(n_677)
);

CKINVDCx11_ASAP7_75t_R g678 ( 
.A(n_629),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_611),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_677),
.Y(n_680)
);

BUFx12f_ASAP7_75t_SL g681 ( 
.A(n_651),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_648),
.B(n_611),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_665),
.A2(n_586),
.B(n_490),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_642),
.A2(n_634),
.B1(n_557),
.B2(n_611),
.Y(n_684)
);

BUFx4f_ASAP7_75t_SL g685 ( 
.A(n_664),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_646),
.A2(n_538),
.B1(n_590),
.B2(n_593),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_648),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_646),
.A2(n_483),
.B1(n_514),
.B2(n_480),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_642),
.A2(n_505),
.B1(n_560),
.B2(n_552),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_644),
.B(n_615),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_649),
.B(n_615),
.Y(n_691)
);

BUFx8_ASAP7_75t_SL g692 ( 
.A(n_641),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_665),
.A2(n_505),
.B1(n_552),
.B2(n_580),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_662),
.A2(n_657),
.B1(n_654),
.B2(n_669),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_643),
.A2(n_503),
.B1(n_511),
.B2(n_483),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_615),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_643),
.A2(n_518),
.B1(n_600),
.B2(n_530),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_675),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_518),
.B1(n_600),
.B2(n_629),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_666),
.B(n_607),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_673),
.A2(n_600),
.B1(n_520),
.B2(n_607),
.Y(n_701)
);

BUFx4f_ASAP7_75t_SL g702 ( 
.A(n_664),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_674),
.A2(n_503),
.B1(n_514),
.B2(n_511),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_651),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_655),
.B(n_605),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_674),
.A2(n_584),
.B1(n_600),
.B2(n_605),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_679),
.B(n_632),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_639),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_SL g709 ( 
.A1(n_651),
.A2(n_471),
.B(n_488),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_663),
.A2(n_600),
.B1(n_605),
.B2(n_587),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_650),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_668),
.A2(n_520),
.B1(n_519),
.B2(n_546),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_670),
.A2(n_519),
.B1(n_474),
.B2(n_481),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_639),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_663),
.A2(n_519),
.B1(n_474),
.B2(n_481),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_678),
.A2(n_500),
.B1(n_501),
.B2(n_507),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_671),
.A2(n_466),
.B1(n_601),
.B2(n_675),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_661),
.A2(n_494),
.B(n_512),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_653),
.A2(n_605),
.B1(n_601),
.B2(n_592),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_678),
.A2(n_507),
.B1(n_501),
.B2(n_500),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_660),
.A2(n_592),
.B1(n_597),
.B2(n_608),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_671),
.A2(n_597),
.B1(n_608),
.B2(n_554),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_645),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_645),
.B(n_585),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_647),
.A2(n_531),
.B1(n_521),
.B2(n_525),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_667),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_694),
.A2(n_612),
.B1(n_675),
.B2(n_659),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_680),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_680),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_686),
.A2(n_609),
.B1(n_651),
.B2(n_612),
.Y(n_731)
);

OAI222xp33_ASAP7_75t_L g732 ( 
.A1(n_689),
.A2(n_609),
.B1(n_521),
.B2(n_525),
.C1(n_527),
.C2(n_531),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_726),
.A2(n_656),
.B1(n_672),
.B2(n_658),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_723),
.A2(n_609),
.B1(n_502),
.B2(n_656),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_684),
.A2(n_527),
.B1(n_526),
.B2(n_491),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_693),
.A2(n_526),
.B1(n_491),
.B2(n_647),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_722),
.A2(n_667),
.B1(n_515),
.B2(n_517),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_687),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_711),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_717),
.A2(n_676),
.B1(n_602),
.B2(n_637),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_720),
.A2(n_515),
.B1(n_504),
.B2(n_635),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_711),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_716),
.A2(n_676),
.B1(n_602),
.B2(n_637),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_SL g744 ( 
.A1(n_703),
.A2(n_515),
.B1(n_504),
.B2(n_635),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_697),
.A2(n_491),
.B1(n_528),
.B2(n_515),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_683),
.A2(n_529),
.B(n_513),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_700),
.B(n_625),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_712),
.A2(n_491),
.B1(n_528),
.B2(n_484),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_700),
.B(n_625),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_713),
.B1(n_721),
.B2(n_701),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_682),
.A2(n_491),
.B1(n_528),
.B2(n_533),
.Y(n_751)
);

OAI22x1_ASAP7_75t_L g752 ( 
.A1(n_725),
.A2(n_633),
.B1(n_565),
.B2(n_589),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_715),
.A2(n_528),
.B1(n_534),
.B2(n_484),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_688),
.A2(n_528),
.B1(n_484),
.B2(n_504),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_695),
.A2(n_724),
.B1(n_710),
.B2(n_699),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_708),
.A2(n_637),
.B1(n_628),
.B2(n_589),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_690),
.B(n_606),
.Y(n_757)
);

AOI222xp33_ASAP7_75t_L g758 ( 
.A1(n_685),
.A2(n_702),
.B1(n_691),
.B2(n_690),
.C1(n_696),
.C2(n_724),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_705),
.A2(n_707),
.B1(n_691),
.B2(n_696),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_705),
.A2(n_504),
.B1(n_486),
.B2(n_628),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_707),
.A2(n_633),
.B1(n_621),
.B2(n_606),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_633),
.B1(n_621),
.B2(n_606),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_714),
.A2(n_621),
.B1(n_606),
.B2(n_576),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_719),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_681),
.A2(n_621),
.B1(n_576),
.B2(n_575),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_738),
.B(n_719),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_727),
.B(n_698),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_758),
.B(n_704),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_747),
.B(n_698),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_733),
.B(n_709),
.C(n_718),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_732),
.B(n_681),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_L g772 ( 
.A1(n_728),
.A2(n_704),
.B1(n_581),
.B2(n_576),
.C(n_575),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_749),
.B(n_704),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_746),
.A2(n_704),
.B1(n_482),
.B2(n_581),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_759),
.B(n_704),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_755),
.A2(n_482),
.B1(n_692),
.B2(n_79),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_757),
.B(n_482),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_746),
.B(n_482),
.C(n_692),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_739),
.B(n_482),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_736),
.A2(n_72),
.B1(n_77),
.B2(n_81),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_764),
.B(n_82),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_729),
.B(n_194),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_SL g783 ( 
.A1(n_755),
.A2(n_83),
.B(n_84),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_730),
.B(n_85),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_752),
.B(n_86),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_742),
.B(n_87),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_762),
.B(n_89),
.Y(n_787)
);

XNOR2xp5_ASAP7_75t_L g788 ( 
.A(n_740),
.B(n_91),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_746),
.B(n_191),
.Y(n_789)
);

NAND4xp25_ASAP7_75t_L g790 ( 
.A(n_734),
.B(n_731),
.C(n_750),
.D(n_744),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_763),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_761),
.B(n_93),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_737),
.B(n_94),
.C(n_95),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_L g794 ( 
.A1(n_762),
.A2(n_96),
.B(n_98),
.Y(n_794)
);

OA211x2_ASAP7_75t_L g795 ( 
.A1(n_778),
.A2(n_765),
.B(n_754),
.C(n_751),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_783),
.B(n_776),
.C(n_787),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_766),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_767),
.B(n_756),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_773),
.B(n_765),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_768),
.B(n_741),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_769),
.B(n_743),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_791),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_770),
.B(n_748),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_775),
.B(n_760),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_779),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_777),
.B(n_748),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_789),
.A2(n_735),
.B(n_753),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_790),
.A2(n_774),
.B1(n_785),
.B2(n_787),
.C(n_794),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_785),
.B(n_745),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_803),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_806),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_803),
.B(n_771),
.Y(n_813)
);

XNOR2xp5_ASAP7_75t_L g814 ( 
.A(n_801),
.B(n_788),
.Y(n_814)
);

XOR2x2_ASAP7_75t_L g815 ( 
.A(n_809),
.B(n_793),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_806),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_797),
.B(n_774),
.Y(n_817)
);

AND2x4_ASAP7_75t_SL g818 ( 
.A(n_800),
.B(n_784),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_798),
.Y(n_819)
);

NAND4xp75_ASAP7_75t_L g820 ( 
.A(n_795),
.B(n_786),
.C(n_792),
.D(n_782),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_796),
.A2(n_780),
.B1(n_772),
.B2(n_781),
.Y(n_821)
);

XNOR2xp5_ASAP7_75t_L g822 ( 
.A(n_815),
.B(n_796),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_818),
.B(n_798),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_816),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_816),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_818),
.Y(n_826)
);

OA22x2_ASAP7_75t_L g827 ( 
.A1(n_822),
.A2(n_814),
.B1(n_813),
.B2(n_811),
.Y(n_827)
);

XNOR2xp5_ASAP7_75t_L g828 ( 
.A(n_822),
.B(n_820),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_824),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_826),
.A2(n_821),
.B1(n_804),
.B2(n_799),
.Y(n_830)
);

XNOR2x1_ASAP7_75t_L g831 ( 
.A(n_826),
.B(n_810),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_823),
.A2(n_821),
.B1(n_810),
.B2(n_802),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_829),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_830),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_832),
.Y(n_836)
);

AO22x2_ASAP7_75t_L g837 ( 
.A1(n_833),
.A2(n_828),
.B1(n_827),
.B2(n_825),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_834),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_835),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_839),
.Y(n_840)
);

O2A1O1Ixp5_ASAP7_75t_SL g841 ( 
.A1(n_838),
.A2(n_836),
.B(n_798),
.C(n_780),
.Y(n_841)
);

O2A1O1Ixp5_ASAP7_75t_SL g842 ( 
.A1(n_837),
.A2(n_819),
.B(n_817),
.C(n_801),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_SL g843 ( 
.A(n_837),
.B(n_800),
.Y(n_843)
);

OA22x2_ASAP7_75t_L g844 ( 
.A1(n_840),
.A2(n_843),
.B1(n_842),
.B2(n_841),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_840),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_840),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_840),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_843),
.A2(n_808),
.B1(n_805),
.B2(n_807),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_843),
.A2(n_819),
.B1(n_812),
.B2(n_808),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_843),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_845),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_846),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_844),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_847),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_848),
.B(n_850),
.Y(n_855)
);

OA22x2_ASAP7_75t_L g856 ( 
.A1(n_849),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_856)
);

NOR2x1_ASAP7_75t_L g857 ( 
.A(n_845),
.B(n_113),
.Y(n_857)
);

AND4x1_ASAP7_75t_L g858 ( 
.A(n_853),
.B(n_114),
.C(n_115),
.D(n_116),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_852),
.B(n_118),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_851),
.B(n_119),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_855),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_861)
);

AND4x1_ASAP7_75t_L g862 ( 
.A(n_857),
.B(n_124),
.C(n_126),
.D(n_128),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_854),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_856),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

XNOR2xp5_ASAP7_75t_L g866 ( 
.A(n_862),
.B(n_189),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_863),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_867)
);

OA22x2_ASAP7_75t_L g868 ( 
.A1(n_864),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_860),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_858),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_861),
.Y(n_871)
);

OAI22x1_ASAP7_75t_L g872 ( 
.A1(n_869),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_865),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_870),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_185),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_866),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_875),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_876),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_872),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_873),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_SL g881 ( 
.A1(n_879),
.A2(n_874),
.B1(n_868),
.B2(n_867),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_880),
.A2(n_184),
.B1(n_159),
.B2(n_162),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_881),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_883),
.A2(n_878),
.B1(n_877),
.B2(n_882),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_884),
.Y(n_885)
);

AOI221xp5_ASAP7_75t_L g886 ( 
.A1(n_885),
.A2(n_158),
.B1(n_163),
.B2(n_166),
.C(n_168),
.Y(n_886)
);

AOI211xp5_ASAP7_75t_L g887 ( 
.A1(n_886),
.A2(n_169),
.B(n_170),
.C(n_171),
.Y(n_887)
);


endmodule