module real_jpeg_31661_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_299;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_273;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_0),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_148),
.B1(n_152),
.B2(n_155),
.Y(n_147)
);

INVx2_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g191 ( 
.A1(n_1),
.A2(n_155),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_155),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_2),
.A2(n_122),
.B1(n_126),
.B2(n_130),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_2),
.A2(n_130),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_130),
.B1(n_259),
.B2(n_264),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_7),
.A2(n_81),
.B1(n_251),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_73),
.B1(n_106),
.B2(n_111),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_10),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_12),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.A3(n_27),
.B1(n_32),
.B2(n_39),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_13),
.A2(n_33),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_13),
.A2(n_64),
.B1(n_205),
.B2(n_211),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_13),
.B(n_157),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_198),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_197),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_179),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_18),
.B(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_118),
.B2(n_119),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_78),
.B1(n_116),
.B2(n_117),
.Y(n_20)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_47),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_22),
.B(n_47),
.Y(n_181)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_25),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_26),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_26),
.Y(n_194)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_26),
.Y(n_263)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_29),
.Y(n_188)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_R g167 ( 
.A(n_33),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_33),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_33),
.B(n_115),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_33),
.B(n_248),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_33),
.A2(n_247),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_39),
.A2(n_132),
.B(n_138),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_41),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_42),
.Y(n_134)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_46),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_46),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_63),
.B2(n_70),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_52),
.A2(n_63),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_62),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_63),
.A2(n_219),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_64),
.A2(n_205),
.B1(n_226),
.B2(n_232),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_64),
.A2(n_274),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

BUFx2_ASAP7_75t_SL g223 ( 
.A(n_68),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_70),
.Y(n_285)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_77),
.Y(n_229)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_84),
.B1(n_105),
.B2(n_115),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22x1_ASAP7_75t_L g189 ( 
.A1(n_80),
.A2(n_190),
.B1(n_191),
.B2(n_196),
.Y(n_189)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

AO21x2_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B(n_98),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_90),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_158),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_131),
.B1(n_147),
.B2(n_156),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_121),
.A2(n_131),
.B1(n_156),
.B2(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_138)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

BUFx4f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.C(n_189),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_181),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_182),
.A2(n_183),
.B1(n_189),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_190),
.A2(n_196),
.B1(n_258),
.B2(n_268),
.Y(n_257)
);

NAND2x1_ASAP7_75t_SL g288 ( 
.A(n_190),
.B(n_191),
.Y(n_288)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2x1_ASAP7_75t_L g287 ( 
.A(n_196),
.B(n_258),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_291),
.B(n_299),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_280),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_236),
.B(n_277),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_224),
.B(n_235),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_216),
.Y(n_203)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_215),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_234),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_272),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_256),
.B1(n_257),
.B2(n_271),
.Y(n_237)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_238),
.B(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_246),
.B1(n_250),
.B2(n_255),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_256),
.B(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_271),
.Y(n_279)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_289),
.C(n_295),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B(n_289),
.C(n_290),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_R g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

NOR2x1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_296),
.Y(n_299)
);


endmodule