module fake_jpeg_28626_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_0),
.C(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_0),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_2),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_73),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_61),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_49),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_55),
.B1(n_65),
.B2(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_64),
.B1(n_51),
.B2(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_65),
.B1(n_64),
.B2(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_56),
.Y(n_107)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_55),
.B(n_47),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_4),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_7),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_50),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_120),
.C(n_125),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_21),
.C(n_22),
.Y(n_136)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_36),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_13),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_129)
);

XOR2x2_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_114),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_14),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_24),
.C(n_26),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_28),
.C(n_29),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.C(n_143),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_31),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_121),
.A2(n_117),
.B(n_115),
.C(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_144),
.B1(n_122),
.B2(n_113),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_33),
.C(n_34),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_148),
.B1(n_127),
.B2(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_142),
.B(n_131),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_134),
.C(n_131),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_151),
.C(n_148),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_146),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_40),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_42),
.Y(n_160)
);


endmodule