module fake_jpeg_11145_n_639 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_639);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_639;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_29),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_69),
.B(n_73),
.Y(n_147)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_76),
.B(n_79),
.Y(n_157)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g192 ( 
.A(n_78),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_85),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

CKINVDCx9p33_ASAP7_75t_R g91 ( 
.A(n_29),
.Y(n_91)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_93),
.Y(n_182)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_102),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_98),
.Y(n_201)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_100),
.Y(n_214)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_23),
.B(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_110),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_16),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_121),
.Y(n_181)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_37),
.Y(n_119)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_59),
.B(n_0),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_44),
.Y(n_124)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_119),
.A2(n_36),
.B1(n_43),
.B2(n_57),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_135),
.A2(n_173),
.B(n_145),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_30),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_137),
.B(n_160),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_32),
.C(n_55),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_143),
.B(n_166),
.C(n_182),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_30),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_153),
.B(n_161),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_28),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_86),
.B(n_28),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_46),
.C(n_55),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_78),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_25),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_171),
.B(n_180),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_62),
.A2(n_36),
.B1(n_57),
.B2(n_43),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_124),
.B(n_25),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_67),
.B(n_50),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_183),
.B(n_190),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_70),
.A2(n_33),
.B1(n_107),
.B2(n_125),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_189),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_67),
.B(n_50),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_65),
.B(n_53),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_197),
.B(n_205),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_85),
.B(n_53),
.Y(n_205)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_92),
.Y(n_208)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_106),
.B(n_38),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_155),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_147),
.A2(n_42),
.B1(n_38),
.B2(n_48),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_216),
.A2(n_239),
.B(n_256),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_157),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_217),
.B(n_229),
.Y(n_298)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_42),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_221),
.B(n_241),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_222),
.Y(n_332)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_147),
.A2(n_127),
.B1(n_126),
.B2(n_123),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_226),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_230),
.B(n_237),
.Y(n_312)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_232),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_174),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_233),
.B(n_234),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_164),
.B(n_174),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_170),
.A2(n_48),
.B1(n_45),
.B2(n_46),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_235),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_130),
.B(n_45),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_192),
.B(n_41),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_240),
.B(n_248),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_41),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_242),
.Y(n_313)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_244),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_245),
.Y(n_321)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_134),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_246),
.Y(n_348)
);

BUFx16f_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_1),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_249),
.B(n_251),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_2),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_252),
.A2(n_133),
.B1(n_214),
.B2(n_213),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_132),
.B(n_64),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_168),
.B(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_254),
.B(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_184),
.A2(n_57),
.B1(n_43),
.B2(n_114),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_158),
.B(n_57),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_263),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_259),
.Y(n_327)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_176),
.Y(n_261)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_261),
.Y(n_346)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_188),
.B(n_43),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_199),
.B(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_267),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_190),
.B(n_3),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_131),
.B(n_115),
.Y(n_268)
);

NAND2x1_ASAP7_75t_L g337 ( 
.A(n_268),
.B(n_202),
.Y(n_337)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_173),
.A2(n_117),
.B1(n_5),
.B2(n_6),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_145),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_140),
.B(n_152),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_273),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_141),
.B(n_4),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_274),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_135),
.A2(n_15),
.B1(n_6),
.B2(n_9),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_148),
.B(n_5),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_14),
.B(n_213),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_149),
.A2(n_6),
.B(n_9),
.C(n_10),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_279),
.A2(n_282),
.B(n_241),
.C(n_221),
.Y(n_339)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_195),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_280),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g281 ( 
.A(n_159),
.Y(n_281)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_154),
.A2(n_9),
.B(n_11),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_286),
.C(n_277),
.Y(n_306)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_142),
.Y(n_283)
);

BUFx4f_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_129),
.B(n_9),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_284),
.Y(n_343)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_156),
.B(n_11),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_133),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_177),
.B(n_11),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_151),
.Y(n_290)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_159),
.A2(n_14),
.B1(n_178),
.B2(n_210),
.Y(n_291)
);

AOI22x1_ASAP7_75t_SL g305 ( 
.A1(n_226),
.A2(n_186),
.B1(n_187),
.B2(n_193),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_305),
.A2(n_306),
.B(n_239),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_252),
.A2(n_207),
.B1(n_203),
.B2(n_198),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_307),
.A2(n_338),
.B1(n_269),
.B2(n_215),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_185),
.C(n_146),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_329),
.C(n_231),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_SL g369 ( 
.A1(n_318),
.A2(n_288),
.B(n_276),
.C(n_223),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_240),
.B(n_138),
.C(n_139),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_163),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_337),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_256),
.A2(n_139),
.B1(n_202),
.B2(n_142),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_268),
.Y(n_380)
);

OR2x2_ASAP7_75t_SL g353 ( 
.A(n_340),
.B(n_279),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_271),
.A2(n_150),
.B1(n_213),
.B2(n_214),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_229),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_353),
.B(n_380),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_249),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_384),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_300),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_360),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_298),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_217),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_361),
.B(n_362),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_247),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_299),
.B(n_236),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_364),
.B(n_365),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_293),
.B(n_247),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_367),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_293),
.B(n_238),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_371),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_369),
.A2(n_388),
.B(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_317),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_328),
.A2(n_251),
.B1(n_254),
.B2(n_270),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_374),
.B1(n_333),
.B2(n_307),
.Y(n_401)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_373),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_328),
.A2(n_216),
.B1(n_286),
.B2(n_281),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_376),
.Y(n_408)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_219),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_382),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_344),
.A2(n_288),
.B1(n_232),
.B2(n_260),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_378),
.A2(n_396),
.B1(n_245),
.B2(n_316),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_268),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_387),
.Y(n_414)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_383),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_322),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_325),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_385),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_299),
.B(n_301),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_391),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_272),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_344),
.A2(n_228),
.B(n_288),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_265),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_392),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_310),
.B(n_224),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_395),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_330),
.B(n_220),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_347),
.B(n_294),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_220),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_406),
.Y(n_439)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_365),
.A2(n_309),
.A3(n_311),
.B1(n_305),
.B2(n_306),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_329),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_422),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_379),
.A2(n_334),
.B1(n_343),
.B2(n_350),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_411),
.A2(n_425),
.B1(n_434),
.B2(n_389),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_338),
.B1(n_333),
.B2(n_340),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_412),
.A2(n_416),
.B1(n_433),
.B2(n_390),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_314),
.B1(n_341),
.B2(n_319),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_303),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_412),
.Y(n_444)
);

OAI32xp33_ASAP7_75t_L g422 ( 
.A1(n_379),
.A2(n_266),
.A3(n_341),
.B1(n_315),
.B2(n_337),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_396),
.A2(n_314),
.B1(n_218),
.B2(n_262),
.Y(n_425)
);

OAI32xp33_ASAP7_75t_L g429 ( 
.A1(n_362),
.A2(n_315),
.A3(n_292),
.B1(n_316),
.B2(n_227),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_354),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_387),
.B(n_394),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_380),
.A2(n_319),
.B1(n_295),
.B2(n_326),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_388),
.A2(n_215),
.B1(n_283),
.B2(n_225),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_367),
.Y(n_435)
);

INVx13_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_368),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_442),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_441),
.B(n_449),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_417),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_381),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_456),
.C(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_320),
.Y(n_449)
);

AOI31xp33_ASAP7_75t_L g451 ( 
.A1(n_432),
.A2(n_417),
.A3(n_397),
.B(n_421),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_457),
.Y(n_472)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_401),
.A2(n_359),
.B1(n_390),
.B2(n_369),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_458),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

INVx13_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_455),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_403),
.B(n_381),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_402),
.B(n_352),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_399),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_400),
.A2(n_359),
.B1(n_353),
.B2(n_394),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_466),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_409),
.A2(n_389),
.B1(n_369),
.B2(n_356),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_461),
.B(n_467),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_399),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_464),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_424),
.B(n_363),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_398),
.B(n_324),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_469),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_400),
.A2(n_397),
.B1(n_398),
.B2(n_416),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_403),
.B(n_421),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_296),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_470),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_456),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_497),
.Y(n_524)
);

OAI32xp33_ASAP7_75t_L g482 ( 
.A1(n_439),
.A2(n_420),
.A3(n_424),
.B1(n_429),
.B2(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_440),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_444),
.A2(n_410),
.B1(n_406),
.B2(n_433),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_484),
.A2(n_499),
.B1(n_445),
.B2(n_443),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_414),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_486),
.B(n_453),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_423),
.C(n_414),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_490),
.C(n_492),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_410),
.C(n_434),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_430),
.C(n_369),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_458),
.A2(n_462),
.B(n_439),
.Y(n_494)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_422),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_404),
.C(n_413),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_447),
.C(n_454),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_444),
.A2(n_404),
.B1(n_425),
.B2(n_405),
.Y(n_499)
);

XOR2x2_ASAP7_75t_L g500 ( 
.A(n_438),
.B(n_413),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_500),
.B(n_464),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_460),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_504),
.B(n_512),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_507),
.A2(n_520),
.B1(n_523),
.B2(n_525),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_483),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_519),
.Y(n_540)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_473),
.Y(n_509)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_509),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_522),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_511),
.A2(n_516),
.B1(n_503),
.B2(n_487),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_513),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_472),
.A2(n_445),
.B1(n_442),
.B2(n_437),
.Y(n_515)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_515),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_491),
.A2(n_470),
.B1(n_467),
.B2(n_459),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_503),
.A2(n_448),
.B(n_450),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_517),
.A2(n_487),
.B(n_501),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_347),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_518),
.B(n_521),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_435),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_489),
.A2(n_450),
.B1(n_405),
.B2(n_419),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_347),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_486),
.B(n_455),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_405),
.B1(n_419),
.B2(n_428),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_480),
.A2(n_455),
.B1(n_426),
.B2(n_376),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_383),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_531),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_480),
.A2(n_426),
.B1(n_382),
.B2(n_355),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_527),
.A2(n_529),
.B1(n_530),
.B2(n_532),
.Y(n_558)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_528),
.Y(n_556)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_471),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_348),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_371),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_481),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_490),
.B(n_345),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_521),
.Y(n_546)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_534),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_506),
.A2(n_481),
.B(n_474),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_537),
.B(n_543),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_500),
.C(n_474),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_538),
.B(n_542),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_541),
.A2(n_547),
.B1(n_550),
.B2(n_553),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_492),
.C(n_484),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_495),
.C(n_477),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_544),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_505),
.A2(n_499),
.B1(n_495),
.B2(n_501),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_545),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_531),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_511),
.A2(n_482),
.B1(n_479),
.B2(n_477),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_533),
.C(n_504),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_524),
.C(n_510),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_507),
.A2(n_471),
.B1(n_502),
.B2(n_493),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_517),
.A2(n_502),
.B1(n_332),
.B2(n_346),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_516),
.A2(n_332),
.B1(n_327),
.B2(n_317),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_562),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_522),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_514),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_563),
.B(n_348),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_576),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_557),
.A2(n_514),
.B(n_345),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_567),
.A2(n_570),
.B(n_549),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_550),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_568),
.B(n_575),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_555),
.A2(n_308),
.B(n_373),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_554),
.B(n_392),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_571),
.B(n_574),
.Y(n_581)
);

BUFx12_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_572),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_392),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_552),
.A2(n_346),
.B1(n_327),
.B2(n_295),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_536),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_577),
.A2(n_578),
.B1(n_541),
.B2(n_556),
.Y(n_584)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_547),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_542),
.C(n_551),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_580),
.A2(n_582),
.B(n_585),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_551),
.C(n_539),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_584),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_579),
.B(n_574),
.C(n_564),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_543),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_592),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_587),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_575),
.A2(n_555),
.B1(n_544),
.B2(n_553),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_588),
.A2(n_589),
.B1(n_593),
.B2(n_569),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_560),
.A2(n_538),
.B1(n_535),
.B2(n_545),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_559),
.A2(n_535),
.B(n_546),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_590),
.A2(n_595),
.B(n_573),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_567),
.B(n_244),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_264),
.C(n_246),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_596),
.B(n_321),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_580),
.B(n_570),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_597),
.B(n_609),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_594),
.B(n_565),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_598),
.A2(n_606),
.B(n_297),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_600),
.A2(n_583),
.B1(n_595),
.B2(n_592),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_586),
.B(n_562),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_602),
.B(n_605),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_576),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_603),
.B(n_608),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_565),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_572),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_607),
.B(n_321),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_582),
.B(n_573),
.Y(n_609)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_611),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_583),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_613),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_604),
.A2(n_572),
.B(n_581),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_618),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_617),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_227),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_610),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_620),
.B(n_621),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_250),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_616),
.B(n_612),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_602),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_628),
.B(n_607),
.Y(n_629)
);

AOI322xp5_ASAP7_75t_L g633 ( 
.A1(n_629),
.A2(n_630),
.A3(n_631),
.B1(n_632),
.B2(n_625),
.C1(n_627),
.C2(n_626),
.Y(n_633)
);

AO21x1_ASAP7_75t_L g630 ( 
.A1(n_622),
.A2(n_613),
.B(n_615),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_624),
.A2(n_619),
.B(n_259),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_633),
.A2(n_634),
.B(n_242),
.Y(n_635)
);

AOI322xp5_ASAP7_75t_L g634 ( 
.A1(n_631),
.A2(n_627),
.A3(n_261),
.B1(n_222),
.B2(n_280),
.C1(n_285),
.C2(n_297),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_287),
.B(n_297),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_636),
.A2(n_243),
.B(n_248),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_637),
.B(n_248),
.Y(n_638)
);

AO21x1_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_280),
.B(n_214),
.Y(n_639)
);


endmodule