module fake_jpeg_7226_n_221 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_221);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_33),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_13),
.B(n_14),
.C(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_13),
.B1(n_20),
.B2(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_34),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_66),
.Y(n_82)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_29),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_45),
.C(n_40),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_30),
.B1(n_35),
.B2(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_32),
.B1(n_62),
.B2(n_63),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_54),
.B(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_36),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_45),
.C(n_29),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.C(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_29),
.C(n_49),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_42),
.C(n_37),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_32),
.B1(n_51),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_36),
.B1(n_28),
.B2(n_55),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_37),
.C(n_33),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_68),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_28),
.C(n_22),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_67),
.B1(n_59),
.B2(n_61),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_92),
.B1(n_101),
.B2(n_63),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_64),
.B1(n_36),
.B2(n_28),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_56),
.B(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_99),
.B1(n_102),
.B2(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_104),
.Y(n_108)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_32),
.B1(n_63),
.B2(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_79),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_81),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_112),
.C(n_119),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_113),
.B(n_104),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_83),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_71),
.B(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_118),
.B1(n_95),
.B2(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_55),
.B1(n_72),
.B2(n_28),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_17),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_123),
.C(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_75),
.C(n_22),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_17),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_113),
.C(n_112),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_124),
.B1(n_108),
.B2(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_138),
.B1(n_119),
.B2(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_17),
.C(n_18),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_139),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_25),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_108),
.C(n_121),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_126),
.C(n_136),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_25),
.C(n_17),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_24),
.C(n_23),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_135),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_24),
.C(n_16),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_137),
.B1(n_128),
.B2(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_148),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_164),
.B(n_168),
.C(n_169),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_141),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_140),
.B1(n_139),
.B2(n_132),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_171),
.B1(n_2),
.B2(n_1),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_146),
.C(n_145),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_182),
.C(n_165),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_144),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_16),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_125),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_127),
.C(n_125),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_8),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_162),
.B(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_195),
.B1(n_185),
.B2(n_174),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_189),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_194),
.B(n_5),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_5),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_9),
.C(n_12),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_192),
.C(n_9),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_15),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_179),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_6),
.B(n_12),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_175),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_4),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_3),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_189),
.C(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.C(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_15),
.C(n_4),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_10),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_213),
.B1(n_205),
.B2(n_10),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_205),
.C(n_213),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_217),
.B1(n_11),
.B2(n_1),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_11),
.C(n_1),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_2),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_2),
.Y(n_221)
);


endmodule