module fake_jpeg_13199_n_260 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_2),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_73),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_30),
.B(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_29),
.B(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_26),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_32),
.Y(n_106)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_28),
.B1(n_37),
.B2(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_82),
.B1(n_93),
.B2(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_33),
.B(n_32),
.C(n_28),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_115),
.B(n_104),
.C(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_26),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_106),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_121),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_78),
.B(n_74),
.C(n_10),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_47),
.B(n_6),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_67),
.B(n_6),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_66),
.B1(n_64),
.B2(n_50),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_125),
.B1(n_157),
.B2(n_155),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_148),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_70),
.B1(n_44),
.B2(n_46),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_84),
.B1(n_105),
.B2(n_144),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_131),
.B1(n_155),
.B2(n_84),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_12),
.B1(n_8),
.B2(n_11),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_143),
.Y(n_178)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_88),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_153),
.Y(n_162)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_94),
.B(n_90),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_104),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_104),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_158),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_101),
.B1(n_118),
.B2(n_111),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_117),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_155),
.B1(n_131),
.B2(n_135),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_138),
.C(n_140),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_181),
.C(n_124),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_182),
.B1(n_184),
.B2(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_84),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_105),
.B1(n_134),
.B2(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_126),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_153),
.B1(n_127),
.B2(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_189),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_159),
.B(n_133),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_147),
.B1(n_148),
.B2(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_202),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

OAI211xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_159),
.B(n_183),
.C(n_172),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_199),
.B(n_190),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_203),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_128),
.B(n_139),
.C(n_162),
.D(n_178),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_193),
.B(n_204),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_181),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_175),
.B1(n_176),
.B2(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_164),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

BUFx4f_ASAP7_75t_SL g220 ( 
.A(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_169),
.B(n_167),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_213),
.B(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_198),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.C(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_161),
.C(n_169),
.Y(n_221)
);

AOI221xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_187),
.B1(n_192),
.B2(n_197),
.C(n_203),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_209),
.A3(n_216),
.B1(n_213),
.B2(n_221),
.C1(n_219),
.C2(n_207),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_188),
.B1(n_214),
.B2(n_200),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_191),
.C(n_220),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_217),
.Y(n_228)
);

OA21x2_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_231),
.B(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_206),
.B1(n_201),
.B2(n_185),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_202),
.Y(n_231)
);

AOI31xp67_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_234),
.A3(n_232),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_212),
.C(n_185),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_224),
.C(n_170),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_223),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_242),
.B(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_246),
.Y(n_248)
);

AOI22x1_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_232),
.B1(n_225),
.B2(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_240),
.B1(n_239),
.B2(n_220),
.Y(n_250)
);

AOI31xp33_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_239),
.A3(n_220),
.B(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_249),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_246),
.B1(n_244),
.B2(n_160),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_250),
.B(n_248),
.Y(n_255)
);

NOR2x1_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_165),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_255),
.A2(n_160),
.B(n_170),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_253),
.C(n_180),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_258),
.A2(n_257),
.B(n_180),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_165),
.Y(n_260)
);


endmodule