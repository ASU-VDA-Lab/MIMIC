module fake_jpeg_1012_n_101 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_29),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_34),
.B1(n_31),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_48),
.B1(n_39),
.B2(n_1),
.Y(n_54)
);

OA22x2_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_39),
.B1(n_37),
.B2(n_33),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.C(n_11),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_8),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_64),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_3),
.C(n_5),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_52),
.B(n_7),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_62),
.C(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_14),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_6),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_17),
.C(n_25),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_73),
.C(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_23),
.B1(n_26),
.B2(n_83),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_85),
.B1(n_82),
.B2(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_93),
.C(n_90),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_91),
.C(n_88),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_81),
.Y(n_101)
);


endmodule