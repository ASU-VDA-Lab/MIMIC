module fake_jpeg_8261_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_22),
.B1(n_19),
.B2(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_46),
.B(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_22),
.B1(n_19),
.B2(n_26),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_48),
.B1(n_20),
.B2(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_22),
.B1(n_19),
.B2(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_31),
.B1(n_18),
.B2(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_18),
.B1(n_21),
.B2(n_28),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_30),
.B(n_29),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_16),
.B(n_38),
.C(n_39),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_64),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_58),
.Y(n_85)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_67),
.Y(n_96)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_16),
.B1(n_17),
.B2(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_72),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_74),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_17),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_37),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_34),
.C(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_36),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_36),
.B1(n_37),
.B2(n_20),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_80),
.B1(n_57),
.B2(n_81),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_36),
.B1(n_34),
.B2(n_9),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_66),
.B1(n_67),
.B2(n_76),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_101),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_77),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_34),
.B(n_2),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_86),
.B(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_113),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_75),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_108),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_13),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_12),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_104),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_0),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_139),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_83),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_127),
.C(n_109),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_135),
.B(n_137),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_84),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_146),
.B(n_123),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_123),
.B(n_115),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_102),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_91),
.B(n_84),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_101),
.B1(n_100),
.B2(n_105),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_105),
.B1(n_100),
.B2(n_94),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_160),
.C(n_128),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_133),
.C(n_141),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_158),
.C(n_134),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_162),
.B1(n_139),
.B2(n_97),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_122),
.B1(n_120),
.B2(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_117),
.C(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_157),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_143),
.B(n_146),
.C(n_137),
.D(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_130),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_109),
.C(n_128),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_9),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_164),
.B1(n_170),
.B2(n_165),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_140),
.A3(n_129),
.B1(n_89),
.B2(n_113),
.C1(n_82),
.C2(n_10),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_153),
.B(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_153),
.B1(n_154),
.B2(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_94),
.B1(n_10),
.B2(n_14),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_166),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_180),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_0),
.C(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_192),
.Y(n_196)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_4),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_4),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_188),
.C(n_189),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_6),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_6),
.C(n_7),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_187),
.C(n_192),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_195),
.B(n_191),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_201),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_199),
.B(n_202),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);


endmodule