module fake_netlist_1_2329_n_622 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_622);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_622;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_42), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_8), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_2), .Y(n_78) );
NOR2xp33_ASAP7_75t_L g79 ( .A(n_52), .B(n_69), .Y(n_79) );
BUFx8_ASAP7_75t_SL g80 ( .A(n_15), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_75), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_0), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_28), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_43), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_29), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
INVx1_ASAP7_75t_SL g89 ( .A(n_3), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_8), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_27), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_40), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_6), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_11), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_21), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_23), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_51), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_60), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_65), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_30), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_31), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_55), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_57), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_68), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_20), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_39), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_50), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_54), .Y(n_116) );
INVx3_ASAP7_75t_L g117 ( .A(n_49), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_5), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_64), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_22), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_24), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_117), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_112), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_118), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_76), .A2(n_34), .B(n_72), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_112), .B(n_1), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_94), .B(n_2), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_76), .A2(n_35), .B(n_71), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_118), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_115), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_115), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_78), .B(n_4), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_117), .B(n_5), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_117), .B(n_6), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_117), .B(n_7), .Y(n_137) );
BUFx8_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_92), .B(n_7), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_108), .B(n_9), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_81), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_88), .Y(n_148) );
INVx4_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_88), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_107), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_77), .B(n_9), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_87), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_90), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_77), .B(n_10), .Y(n_162) );
INVxp67_ASAP7_75t_SL g163 ( .A(n_138), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_141), .B(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_155), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_149), .B(n_99), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_141), .B(n_95), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_155), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_122), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_139), .A2(n_93), .B1(n_95), .B2(n_90), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_149), .B(n_121), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_141), .B(n_93), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_149), .B(n_120), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_139), .A2(n_90), .B1(n_104), .B2(n_105), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_149), .B(n_110), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_153), .B(n_110), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_141), .B(n_120), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_143), .A2(n_90), .B1(n_116), .B2(n_114), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_153), .B(n_83), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_162), .B(n_89), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_143), .B(n_119), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_138), .Y(n_187) );
AND3x4_ASAP7_75t_L g188 ( .A(n_162), .B(n_80), .C(n_148), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_161), .B(n_119), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_122), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_161), .B(n_116), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_150), .A2(n_156), .B1(n_159), .B2(n_154), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_122), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_122), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_150), .A2(n_90), .B1(n_113), .B2(n_114), .Y(n_198) );
INVx4_ASAP7_75t_SL g199 ( .A(n_122), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_154), .B(n_113), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_140), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_156), .B(n_102), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_157), .B(n_98), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_157), .B(n_91), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_127), .A2(n_89), .B1(n_86), .B2(n_111), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_137), .B(n_109), .Y(n_215) );
INVx6_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_147), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_123), .B(n_109), .Y(n_219) );
INVx5_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_128), .B(n_106), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_202), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_187), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_163), .B(n_138), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_171), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_191), .B(n_128), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_193), .B(n_133), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_174), .B(n_145), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_171), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_174), .B(n_145), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_171), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
AOI21x1_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_129), .B(n_126), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_180), .A2(n_130), .B1(n_125), .B2(n_124), .Y(n_237) );
BUFx12f_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_189), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_195), .B(n_103), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_195), .B(n_102), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_219), .B(n_136), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_206), .A2(n_130), .B1(n_124), .B2(n_125), .Y(n_244) );
NOR2xp67_ASAP7_75t_L g245 ( .A(n_209), .B(n_151), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
AND2x2_ASAP7_75t_SL g248 ( .A(n_181), .B(n_168), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_189), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_192), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
BUFx12f_ASAP7_75t_SL g252 ( .A(n_167), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_177), .B(n_145), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_185), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_179), .A2(n_101), .B1(n_96), .B2(n_100), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_196), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_197), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g261 ( .A1(n_183), .A2(n_126), .B1(n_129), .B2(n_100), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_165), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_219), .B(n_136), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_219), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_177), .B(n_97), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_168), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_166), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_168), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_175), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_221), .B(n_131), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_197), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_172), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_176), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_175), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_190), .B(n_132), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_212), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_210), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_211), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_188), .Y(n_282) );
OR2x4_ASAP7_75t_L g283 ( .A(n_186), .B(n_188), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_227), .B(n_190), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_255), .B(n_175), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_232), .Y(n_286) );
OR2x6_ASAP7_75t_L g287 ( .A(n_238), .B(n_181), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_239), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_239), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_252), .B(n_204), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_238), .Y(n_291) );
CKINVDCx8_ASAP7_75t_R g292 ( .A(n_256), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_248), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_228), .A2(n_186), .B(n_164), .C(n_201), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_255), .B(n_190), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_268), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_239), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_248), .B(n_194), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_273), .B(n_194), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g302 ( .A1(n_265), .A2(n_215), .B1(n_207), .B2(n_214), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_222), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_256), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_262), .B(n_194), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_248), .A2(n_201), .B1(n_203), .B2(n_178), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_225), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_265), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_242), .A2(n_203), .B(n_201), .C(n_173), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_282), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_273), .B(n_178), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_249), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_282), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_268), .B(n_131), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_233), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_243), .B(n_215), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_270), .Y(n_320) );
O2A1O1Ixp5_ASAP7_75t_L g321 ( .A1(n_224), .A2(n_218), .B(n_212), .C(n_79), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_249), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_270), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_243), .B(n_158), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_264), .B(n_173), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_263), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_264), .B(n_158), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_263), .Y(n_330) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_270), .B(n_216), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_300), .B(n_264), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_284), .A2(n_229), .B(n_254), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_303), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_291), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_300), .A2(n_252), .B1(n_271), .B2(n_277), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_301), .B(n_237), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_294), .A2(n_277), .B1(n_266), .B2(n_223), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_294), .B(n_271), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_321), .A2(n_236), .B(n_126), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_287), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_327), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_294), .A2(n_322), .B1(n_286), .B2(n_319), .Y(n_343) );
CKINVDCx11_ASAP7_75t_R g344 ( .A(n_291), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_SL g346 ( .A1(n_295), .A2(n_223), .B(n_231), .C(n_280), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_244), .B1(n_278), .B2(n_271), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_287), .B(n_269), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_306), .B(n_269), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_327), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_290), .A2(n_257), .B1(n_275), .B2(n_276), .C(n_272), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_330), .A2(n_275), .B1(n_272), .B2(n_276), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
CKINVDCx11_ASAP7_75t_R g355 ( .A(n_304), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_292), .A2(n_283), .B1(n_245), .B2(n_241), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_314), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_292), .A2(n_283), .B1(n_281), .B2(n_280), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_287), .B(n_281), .Y(n_360) );
CKINVDCx6p67_ASAP7_75t_R g361 ( .A(n_287), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_347), .A2(n_302), .B1(n_330), .B2(n_283), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_332), .B(n_306), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_332), .B(n_342), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_355), .A2(n_304), .B1(n_309), .B2(n_306), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_359), .A2(n_309), .B1(n_315), .B2(n_311), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_352), .A2(n_312), .B1(n_319), .B2(n_325), .C(n_329), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_353), .A2(n_296), .B1(n_285), .B2(n_326), .Y(n_369) );
CKINVDCx10_ASAP7_75t_R g370 ( .A(n_344), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_334), .A2(n_311), .B1(n_315), .B2(n_296), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_351), .B(n_325), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_345), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_353), .A2(n_296), .B1(n_285), .B2(n_317), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_351), .B(n_314), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_361), .A2(n_323), .B1(n_285), .B2(n_298), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_337), .A2(n_329), .B1(n_317), .B2(n_323), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_348), .A2(n_317), .B1(n_324), .B2(n_313), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_356), .A2(n_310), .B1(n_305), .B2(n_320), .C(n_316), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_348), .A2(n_324), .B1(n_313), .B2(n_298), .Y(n_381) );
AOI33xp33_ASAP7_75t_L g382 ( .A1(n_343), .A2(n_132), .A3(n_198), .B1(n_182), .B2(n_106), .B3(n_97), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_350), .B(n_293), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_348), .A2(n_298), .B1(n_313), .B2(n_324), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_341), .B1(n_338), .B2(n_360), .C1(n_348), .C2(n_335), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_360), .A2(n_126), .B1(n_129), .B2(n_288), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_335), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_375), .A2(n_360), .B1(n_341), .B2(n_339), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_370), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_367), .A2(n_360), .B1(n_361), .B2(n_350), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_373), .B(n_345), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_362), .A2(n_336), .B1(n_339), .B2(n_346), .C(n_261), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_365), .B(n_349), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_388), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_374), .A2(n_358), .B1(n_357), .B2(n_354), .C(n_349), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_358), .B1(n_357), .B2(n_354), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_362), .A2(n_198), .B1(n_182), .B2(n_333), .C(n_331), .Y(n_398) );
NAND3xp33_ASAP7_75t_SL g399 ( .A(n_371), .B(n_146), .C(n_151), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_378), .A2(n_331), .B1(n_357), .B2(n_354), .C(n_349), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_369), .A2(n_358), .B1(n_299), .B2(n_289), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_364), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_373), .B(n_288), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_377), .A2(n_146), .A3(n_151), .B1(n_158), .B2(n_218), .B3(n_289), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_383), .B(n_299), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_383), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_376), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_376), .B(n_340), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_365), .B(n_129), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_376), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_372), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_146), .A3(n_152), .B(n_279), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_363), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_384), .A2(n_340), .B(n_236), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_368), .A2(n_147), .B1(n_142), .B2(n_152), .C1(n_160), .C2(n_199), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_363), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_366), .B(n_10), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_385), .B(n_147), .Y(n_421) );
OAI21x1_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_226), .B(n_230), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_413), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_420), .A2(n_380), .B1(n_379), .B2(n_142), .C(n_152), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_415), .B(n_11), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_395), .A2(n_152), .B1(n_387), .B2(n_160), .C(n_205), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_396), .B(n_160), .C(n_382), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_392), .Y(n_428) );
NOR3xp33_ASAP7_75t_L g429 ( .A(n_399), .B(n_370), .C(n_279), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_397), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_415), .B(n_12), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_415), .B(n_13), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_392), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
OAI33xp33_ASAP7_75t_L g438 ( .A1(n_404), .A2(n_14), .A3(n_16), .B1(n_160), .B2(n_251), .B3(n_250), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_408), .B(n_160), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_230), .B(n_226), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_419), .B(n_220), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_417), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_411), .B(n_17), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_205), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_416), .B(n_18), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_421), .B(n_208), .C(n_217), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_419), .B(n_220), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_417), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_416), .B(n_220), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_403), .B(n_208), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_416), .B(n_25), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_391), .B(n_220), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_389), .A2(n_328), .B1(n_318), .B2(n_208), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_26), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_421), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_406), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_400), .B(n_208), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_393), .B(n_213), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_422), .B(n_33), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_414), .A2(n_216), .B1(n_213), .B2(n_217), .C(n_259), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_405), .A2(n_328), .B1(n_318), .B2(n_213), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_422), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_418), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_425), .B(n_398), .C(n_217), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_455), .B(n_213), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_436), .B(n_390), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_455), .B(n_217), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_441), .B(n_390), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_455), .B(n_36), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_423), .B(n_37), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_457), .B(n_38), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_436), .B(n_44), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_428), .B(n_216), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_462), .B(n_45), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_427), .A2(n_328), .B(n_318), .C(n_53), .Y(n_484) );
NAND5xp2_ASAP7_75t_L g485 ( .A(n_469), .B(n_46), .C(n_48), .D(n_58), .E(n_59), .Y(n_485) );
NAND4xp75_ASAP7_75t_L g486 ( .A(n_425), .B(n_63), .C(n_66), .D(n_67), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_462), .B(n_70), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_459), .B(n_74), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_457), .B(n_199), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_459), .B(n_328), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_457), .B(n_199), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_423), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_433), .B(n_328), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_461), .B(n_318), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_443), .B(n_318), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_433), .B(n_251), .Y(n_496) );
AOI21xp5_ASAP7_75t_SL g497 ( .A1(n_449), .A2(n_233), .B(n_234), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_434), .B(n_250), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_469), .B(n_274), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_443), .B(n_274), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_443), .B(n_246), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_460), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_437), .B(n_246), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_432), .A2(n_260), .B1(n_259), .B2(n_235), .C(n_240), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_431), .B(n_235), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_431), .B(n_233), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_460), .B(n_240), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_431), .B(n_234), .Y(n_512) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_445), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_448), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_439), .B(n_234), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_431), .B(n_440), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_440), .B(n_234), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_478), .B(n_440), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_473), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_475), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_498), .B(n_440), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_473), .B(n_438), .Y(n_523) );
OA22x2_ASAP7_75t_L g524 ( .A1(n_492), .A2(n_448), .B1(n_454), .B2(n_465), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_507), .B(n_445), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_504), .B(n_445), .Y(n_526) );
OAI21xp5_ASAP7_75t_SL g527 ( .A1(n_484), .A2(n_429), .B(n_427), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_514), .A2(n_464), .B1(n_466), .B2(n_454), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_476), .Y(n_529) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_500), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_501), .B(n_445), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_516), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_484), .A2(n_458), .B1(n_456), .B2(n_424), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g535 ( .A1(n_481), .A2(n_464), .A3(n_450), .B1(n_444), .B2(n_452), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_481), .A2(n_426), .B1(n_465), .B2(n_467), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_516), .B(n_468), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_508), .B(n_442), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_508), .B(n_442), .Y(n_539) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_479), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_453), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_502), .B(n_446), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_486), .B(n_446), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_490), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_495), .B(n_442), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_502), .B(n_468), .Y(n_547) );
XNOR2x1_ASAP7_75t_L g548 ( .A(n_477), .B(n_447), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_471), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_513), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_503), .B(n_465), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_494), .B(n_447), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
NAND2xp33_ASAP7_75t_SL g554 ( .A(n_548), .B(n_483), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_523), .B(n_485), .C(n_470), .D(n_487), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_521), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_546), .B(n_471), .Y(n_557) );
OAI211xp5_ASAP7_75t_SL g558 ( .A1(n_523), .A2(n_488), .B(n_496), .C(n_499), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_532), .A2(n_477), .B1(n_480), .B2(n_510), .C(n_474), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_524), .A2(n_480), .B1(n_517), .B2(n_512), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_529), .B(n_493), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_525), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_522), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_550), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_533), .B(n_509), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_533), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_550), .Y(n_567) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_548), .B(n_491), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_518), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_537), .B(n_509), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_524), .A2(n_463), .B(n_515), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_540), .B(n_491), .Y(n_572) );
AOI321xp33_ASAP7_75t_L g573 ( .A1(n_535), .A2(n_489), .A3(n_505), .B1(n_506), .B2(n_497), .C(n_234), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
NAND3xp33_ASAP7_75t_SL g575 ( .A(n_527), .B(n_489), .C(n_497), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g576 ( .A1(n_543), .A2(n_253), .B(n_258), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_536), .A2(n_253), .B1(n_258), .B2(n_539), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g578 ( .A(n_552), .B(n_253), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_538), .A2(n_253), .B1(n_258), .B2(n_534), .Y(n_579) );
NAND2xp33_ASAP7_75t_SL g580 ( .A(n_526), .B(n_258), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_530), .B(n_549), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_528), .B(n_531), .Y(n_582) );
AOI31xp33_ASAP7_75t_L g583 ( .A1(n_528), .A2(n_551), .A3(n_542), .B(n_545), .Y(n_583) );
NOR2xp33_ASAP7_75t_SL g584 ( .A(n_541), .B(n_547), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_523), .A2(n_546), .B1(n_519), .B2(n_485), .Y(n_585) );
XNOR2xp5_ASAP7_75t_L g586 ( .A(n_519), .B(n_390), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_546), .B(n_544), .Y(n_587) );
OAI211xp5_ASAP7_75t_SL g588 ( .A1(n_546), .A2(n_355), .B(n_473), .C(n_523), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_523), .A2(n_546), .B1(n_519), .B2(n_485), .Y(n_589) );
AOI211xp5_ASAP7_75t_L g590 ( .A1(n_527), .A2(n_523), .B(n_485), .C(n_535), .Y(n_590) );
AOI211xp5_ASAP7_75t_L g591 ( .A1(n_590), .A2(n_588), .B(n_554), .C(n_555), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_583), .A2(n_582), .B(n_558), .C(n_587), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_554), .A2(n_582), .B1(n_561), .B2(n_562), .C(n_567), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_575), .B(n_571), .C(n_564), .Y(n_594) );
XOR2xp5_ASAP7_75t_L g595 ( .A(n_586), .B(n_568), .Y(n_595) );
INVxp33_ASAP7_75t_L g596 ( .A(n_578), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_563), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_567), .A2(n_564), .B(n_589), .C(n_585), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_561), .B(n_569), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_560), .A2(n_585), .B1(n_589), .B2(n_574), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_584), .A2(n_573), .B1(n_577), .B2(n_572), .C(n_579), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_596), .A2(n_572), .B1(n_559), .B2(n_565), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_597), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_601), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_593), .B(n_576), .Y(n_607) );
NAND3xp33_ASAP7_75t_SL g608 ( .A(n_591), .B(n_579), .C(n_580), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_603), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_592), .A2(n_566), .B(n_581), .C(n_570), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_610), .A2(n_600), .B1(n_598), .B2(n_594), .C(n_595), .Y(n_611) );
XOR2xp5_ASAP7_75t_L g612 ( .A(n_608), .B(n_557), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_605), .B(n_594), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_604), .B(n_599), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_611), .A2(n_607), .B1(n_602), .B2(n_606), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_613), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_616), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_615), .Y(n_618) );
OR3x1_ASAP7_75t_L g619 ( .A(n_618), .B(n_612), .C(n_614), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_619), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_620), .B(n_617), .Y(n_621) );
AO21x2_ASAP7_75t_L g622 ( .A1(n_621), .A2(n_607), .B(n_609), .Y(n_622) );
endmodule