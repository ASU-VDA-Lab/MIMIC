module fake_jpeg_13579_n_407 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_54),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_21),
.B(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_60),
.Y(n_127)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_14),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_62),
.B(n_66),
.Y(n_141)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_67),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_22),
.B(n_8),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_69),
.Y(n_144)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_72),
.Y(n_159)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_18),
.Y(n_74)
);

CKINVDCx9p33_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_20),
.A2(n_11),
.B1(n_3),
.B2(n_6),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_75),
.A2(n_51),
.B1(n_37),
.B2(n_31),
.Y(n_145)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_79),
.B(n_81),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_18),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_80),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_0),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_23),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_83),
.B(n_87),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_36),
.B(n_0),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_23),
.B(n_11),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_97),
.Y(n_114)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_27),
.B(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_94),
.B(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_28),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_28),
.B(n_51),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_29),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_105),
.B(n_107),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_33),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_33),
.B(n_13),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_110),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_35),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_31),
.Y(n_146)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_44),
.B1(n_49),
.B2(n_45),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_113),
.A2(n_177),
.B1(n_141),
.B2(n_159),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_39),
.B1(n_26),
.B2(n_30),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_145),
.B1(n_153),
.B2(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_120),
.B(n_170),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_56),
.A2(n_38),
.B1(n_26),
.B2(n_30),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_149),
.B1(n_177),
.B2(n_58),
.Y(n_183)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_42),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_134),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_42),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_154),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_85),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_77),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_50),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_155),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_58),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_73),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_67),
.A2(n_93),
.B1(n_99),
.B2(n_88),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_92),
.A2(n_76),
.B1(n_109),
.B2(n_74),
.Y(n_177)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_183),
.B(n_219),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_199),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_84),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_186),
.B(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_84),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_117),
.B(n_90),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_193),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_78),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_194),
.B(n_196),
.Y(n_273)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_90),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_134),
.A2(n_61),
.B1(n_118),
.B2(n_153),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_114),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_198),
.B(n_202),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_144),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_144),
.B1(n_149),
.B2(n_125),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_116),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_208),
.B(n_215),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_130),
.A2(n_137),
.B1(n_169),
.B2(n_128),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_113),
.B(n_141),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_214),
.C(n_224),
.Y(n_268)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_113),
.B(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_122),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_119),
.B(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_221),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_142),
.A2(n_172),
.B1(n_115),
.B2(n_159),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_240),
.B1(n_199),
.B2(n_223),
.Y(n_248)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_126),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_151),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_179),
.A2(n_176),
.B1(n_178),
.B2(n_166),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_138),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_231),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_123),
.C(n_132),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_227),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_124),
.Y(n_227)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_147),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_150),
.B(n_129),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_239),
.Y(n_250)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_127),
.B(n_117),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_121),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_116),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_167),
.B(n_143),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_184),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_256),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_192),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_197),
.B1(n_209),
.B2(n_232),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_258),
.A2(n_271),
.B1(n_281),
.B2(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_201),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_261),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_213),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_222),
.A2(n_187),
.B1(n_214),
.B2(n_210),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_263),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_235),
.B1(n_233),
.B2(n_228),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_272),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_191),
.B(n_204),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_218),
.A2(n_207),
.B1(n_212),
.B2(n_195),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_200),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_221),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_282),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_205),
.A2(n_240),
.B1(n_203),
.B2(n_238),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_188),
.B(n_185),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_188),
.B(n_215),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_230),
.A2(n_201),
.B1(n_197),
.B2(n_211),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_229),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_290),
.Y(n_320)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_278),
.B(n_273),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_252),
.A3(n_296),
.B1(n_306),
.B2(n_291),
.C1(n_308),
.C2(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_254),
.A2(n_268),
.B(n_264),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_301),
.A2(n_307),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_246),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_309),
.Y(n_327)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_SL g306 ( 
.A(n_256),
.B(n_246),
.C(n_278),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_315),
.C(n_275),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_254),
.B(n_284),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_247),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_286),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_258),
.B1(n_253),
.B2(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_317),
.B1(n_319),
.B2(n_279),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_261),
.A2(n_244),
.B(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_250),
.C(n_249),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_274),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_259),
.A2(n_243),
.B1(n_249),
.B2(n_271),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_251),
.A2(n_277),
.B1(n_265),
.B2(n_275),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_325),
.B1(n_341),
.B2(n_293),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_318),
.A2(n_286),
.B1(n_285),
.B2(n_269),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_311),
.A2(n_277),
.B1(n_274),
.B2(n_257),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_329),
.C(n_342),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_330),
.B(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_281),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_336),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_252),
.B1(n_303),
.B2(n_297),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_334),
.A2(n_289),
.B1(n_333),
.B2(n_331),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_298),
.B(n_252),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_307),
.A2(n_301),
.B(n_303),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_293),
.B(n_294),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_308),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_335),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_299),
.B1(n_296),
.B2(n_314),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_312),
.C(n_305),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_322),
.B(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

AOI221xp5_ASAP7_75t_L g348 ( 
.A1(n_323),
.A2(n_310),
.B1(n_316),
.B2(n_302),
.C(n_299),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_348),
.B(n_336),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_360),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_300),
.Y(n_351)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_341),
.Y(n_353)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_313),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_359),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_357),
.A2(n_358),
.B1(n_325),
.B2(n_339),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_333),
.B1(n_335),
.B2(n_320),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_342),
.C(n_321),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_363),
.A2(n_365),
.B1(n_372),
.B2(n_352),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_337),
.B1(n_321),
.B2(n_328),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_327),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_378),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_376),
.B(n_380),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_344),
.C(n_360),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_383),
.C(n_381),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_350),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_379),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_344),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_370),
.A2(n_349),
.B(n_343),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_371),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_360),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_370),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_345),
.C(n_359),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_386),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_374),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_390),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_363),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_394),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_387),
.A2(n_362),
.B1(n_374),
.B2(n_367),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_353),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_397),
.C(n_391),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_388),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_385),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_361),
.B1(n_351),
.B2(n_354),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_394),
.A2(n_348),
.B1(n_373),
.B2(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_401),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_399),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.C(n_398),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_396),
.Y(n_405)
);

XNOR2x2_ASAP7_75t_SL g407 ( 
.A(n_406),
.B(n_405),
.Y(n_407)
);


endmodule