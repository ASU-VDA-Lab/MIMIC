module fake_jpeg_27347_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_53),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_42),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_55),
.B1(n_62),
.B2(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_45),
.B1(n_51),
.B2(n_49),
.Y(n_92)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_86),
.Y(n_90)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_42),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_48),
.B1(n_56),
.B2(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_84),
.B1(n_64),
.B2(n_76),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_1),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_2),
.B(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_80),
.B1(n_83),
.B2(n_81),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_88),
.B1(n_89),
.B2(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_60),
.B1(n_86),
.B2(n_8),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_5),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_105),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

AOI21x1_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_7),
.B(n_9),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_16),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_19),
.B(n_25),
.C(n_26),
.Y(n_117)
);

OAI21x1_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_27),
.B(n_28),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_35),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_37),
.Y(n_121)
);


endmodule