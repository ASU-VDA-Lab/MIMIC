module fake_jpeg_10504_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_18),
.B1(n_14),
.B2(n_22),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_46),
.B1(n_22),
.B2(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_47),
.Y(n_59)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_18),
.B1(n_15),
.B2(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_61),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_62),
.C(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_25),
.B1(n_48),
.B2(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_36),
.C(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_40),
.B1(n_51),
.B2(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_43),
.B1(n_25),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_81),
.B1(n_48),
.B2(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_60),
.C(n_56),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_82),
.C(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.C(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_57),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_54),
.B(n_51),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_26),
.B(n_13),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_53),
.C(n_52),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_73),
.B1(n_79),
.B2(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_43),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_19),
.C(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_101),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_99),
.C(n_107),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_69),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_24),
.B(n_23),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_90),
.B1(n_81),
.B2(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_23),
.B1(n_20),
.B2(n_13),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_105),
.B(n_84),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_111),
.B1(n_105),
.B2(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_90),
.C(n_89),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_98),
.C(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_109),
.Y(n_122)
);

OA21x2_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_109),
.B(n_114),
.Y(n_118)
);

AOI31xp67_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_50),
.A3(n_38),
.B(n_12),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_119),
.B1(n_26),
.B2(n_3),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_106),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_50),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_10),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_132),
.B1(n_4),
.B2(n_6),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_26),
.B1(n_10),
.B2(n_7),
.C(n_8),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_4),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_130),
.B(n_6),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_7),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_7),
.Y(n_138)
);


endmodule