module fake_jpeg_5463_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_14),
.B1(n_18),
.B2(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_14),
.B1(n_12),
.B2(n_10),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_24),
.B1(n_22),
.B2(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_27),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_32),
.B1(n_38),
.B2(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_55),
.B1(n_44),
.B2(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_44),
.B1(n_40),
.B2(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_42),
.B1(n_48),
.B2(n_26),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_29),
.B1(n_37),
.B2(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_23),
.C(n_36),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_62),
.B1(n_52),
.B2(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_36),
.B1(n_25),
.B2(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_17),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_75),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_50),
.C(n_65),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_78),
.B1(n_71),
.B2(n_69),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_65),
.C(n_57),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_77),
.C(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_89),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_92),
.B1(n_88),
.B2(n_87),
.C(n_17),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_73),
.C(n_17),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_17),
.B(n_8),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_3),
.B(n_4),
.Y(n_95)
);

AOI321xp33_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_84),
.A3(n_83),
.B1(n_80),
.B2(n_81),
.C(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_17),
.B1(n_19),
.B2(n_5),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_98),
.B1(n_9),
.B2(n_5),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_102),
.C(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_105),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_3),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_4),
.C(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule