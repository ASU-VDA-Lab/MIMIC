module fake_jpeg_11414_n_197 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_0),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_57),
.B1(n_68),
.B2(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_110),
.B1(n_71),
.B2(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_73),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_77),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_76),
.B1(n_68),
.B2(n_57),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_108),
.B1(n_84),
.B2(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_62),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_71),
.B1(n_74),
.B2(n_84),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_60),
.B1(n_80),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_120),
.B1(n_131),
.B2(n_132),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_102),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_10),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_93),
.B1(n_59),
.B2(n_69),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_71),
.A3(n_79),
.B1(n_82),
.B2(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_124),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_75),
.B1(n_61),
.B2(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_122),
.B1(n_131),
.B2(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_1),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_33),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_27),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_61),
.B1(n_94),
.B2(n_85),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_85),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_28),
.C(n_53),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_39),
.CI(n_40),
.CON(n_168),
.SN(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_12),
.B(n_13),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_31),
.B(n_34),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_155),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_167),
.B(n_172),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_36),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_163),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_41),
.B(n_44),
.Y(n_181)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

AOI22x1_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_181),
.B(n_158),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_138),
.B1(n_152),
.B2(n_142),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_135),
.C(n_43),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_179),
.C(n_175),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_166),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_185),
.B(n_180),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_189),
.B(n_180),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_174),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_156),
.B(n_173),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_157),
.C(n_163),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_46),
.CI(n_49),
.CON(n_195),
.SN(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_50),
.B(n_52),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_54),
.Y(n_197)
);


endmodule