module fake_ariane_2660_n_1966 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1966);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1966;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_103),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_84),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_60),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_20),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_119),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_38),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_126),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_5),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_55),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_65),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_44),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_3),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_21),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_60),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_83),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_38),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_87),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_61),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_42),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_58),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_4),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_21),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_94),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_28),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_181),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_167),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_5),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_111),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_64),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_65),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_183),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_82),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_89),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_59),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_196),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_42),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_44),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_131),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_96),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_180),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_72),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_78),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_7),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_29),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_41),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_2),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_86),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_53),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_104),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_58),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_33),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_64),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_69),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_51),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_34),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_57),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_105),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_75),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_115),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_140),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_142),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_162),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_32),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_146),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_15),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_125),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_10),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_141),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_156),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_59),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_6),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_97),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_184),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_107),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_80),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_31),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_154),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_13),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_165),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_188),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_71),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_79),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_48),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_50),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_30),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_85),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_17),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_17),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_6),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_172),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_19),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_81),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_185),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_4),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_54),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_66),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_122),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_72),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_92),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_143),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_25),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_187),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_110),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_157),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_47),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_31),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_178),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_114),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_32),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_88),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_132),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_139),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_135),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_69),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_61),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_63),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_18),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_55),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_52),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_71),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_63),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_193),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_192),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_161),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_74),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_116),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_128),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_56),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_30),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_70),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_102),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_171),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_176),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_182),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_158),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_170),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_29),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_39),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_136),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_169),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_8),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_138),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_186),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_109),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_35),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_144),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_1),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_73),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_201),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_270),
.B(n_0),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_244),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_267),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_200),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_270),
.B(n_0),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_200),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_313),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_307),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_231),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_223),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_307),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_231),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_323),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_323),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_3),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_223),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_227),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_225),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_225),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_204),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_7),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_8),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_229),
.B(n_9),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_229),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_213),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_237),
.B(n_9),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_221),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_260),
.B(n_266),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_245),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_245),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_217),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_232),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_237),
.B(n_326),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_234),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_242),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_234),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_240),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_220),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_224),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_240),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_274),
.Y(n_437)
);

INVx4_ASAP7_75t_SL g438 ( 
.A(n_219),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_215),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_326),
.B(n_11),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_258),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_258),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_235),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_236),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_238),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_269),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_239),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_269),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_294),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_249),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_311),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_286),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_221),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_294),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_302),
.B(n_11),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_302),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_250),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_310),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_251),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_254),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_310),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_255),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_318),
.B(n_13),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_318),
.B(n_14),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_256),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_263),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_271),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_324),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_324),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_288),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_221),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_328),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_328),
.Y(n_473)
);

BUFx2_ASAP7_75t_SL g474 ( 
.A(n_215),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_332),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_272),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_205),
.B(n_14),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_332),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_322),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_339),
.B(n_16),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_276),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_339),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_R g483 ( 
.A(n_199),
.B(n_194),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_219),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_219),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_205),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_268),
.Y(n_487)
);

BUFx6f_ASAP7_75t_SL g488 ( 
.A(n_215),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_278),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_282),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_396),
.B(n_344),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_463),
.A2(n_197),
.B(n_344),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_418),
.B(n_242),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_396),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_395),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_412),
.A2(n_390),
.B1(n_308),
.B2(n_359),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_428),
.A2(n_452),
.B1(n_470),
.B2(n_437),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_405),
.B(n_268),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_413),
.B(n_347),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_406),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_471),
.B(n_268),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_420),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_430),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_432),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_436),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_424),
.B(n_347),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_410),
.B(n_242),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_442),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_446),
.B(n_350),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_446),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_471),
.B(n_341),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_448),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_480),
.A2(n_365),
.B(n_350),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_449),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_454),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_474),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_454),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_456),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_283),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_456),
.B(n_341),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_392),
.A2(n_209),
.B1(n_216),
.B2(n_218),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_474),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_458),
.B(n_461),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_426),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_458),
.B(n_341),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_365),
.Y(n_555)
);

AND3x1_ASAP7_75t_L g556 ( 
.A(n_417),
.B(n_216),
.C(n_209),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_469),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_472),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_475),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_404),
.A2(n_280),
.B1(n_391),
.B2(n_329),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_488),
.B(n_215),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_495),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_556),
.A2(n_425),
.B1(n_489),
.B2(n_397),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_544),
.B(n_488),
.Y(n_575)
);

AOI22x1_ASAP7_75t_L g576 ( 
.A1(n_498),
.A2(n_477),
.B1(n_440),
.B2(n_482),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_544),
.B(n_415),
.Y(n_577)
);

AND2x2_ASAP7_75t_SL g578 ( 
.A(n_568),
.B(n_197),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_495),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_501),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_497),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_570),
.Y(n_584)
);

INVxp33_ASAP7_75t_L g585 ( 
.A(n_547),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_550),
.B(n_488),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_501),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_550),
.B(n_439),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_551),
.B(n_423),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_568),
.B(n_421),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_503),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_501),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_551),
.B(n_453),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_530),
.A2(n_416),
.B1(n_455),
.B2(n_419),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_570),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_509),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_551),
.B(n_507),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_SL g601 ( 
.A1(n_530),
.A2(n_477),
.B(n_440),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_509),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_514),
.B(n_451),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_503),
.B(n_427),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_509),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_509),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_516),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_516),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_508),
.B(n_487),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_541),
.A2(n_416),
.B1(n_464),
.B2(n_486),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_507),
.B(n_482),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_507),
.B(n_434),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_549),
.A2(n_393),
.B1(n_422),
.B2(n_483),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_514),
.B(n_435),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_553),
.B(n_429),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_516),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_514),
.B(n_443),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_518),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_518),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_518),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_498),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_498),
.B(n_502),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_498),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_518),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_518),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_518),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_520),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_498),
.B(n_444),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_552),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_520),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_537),
.B(n_445),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_520),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_547),
.A2(n_394),
.B1(n_399),
.B2(n_401),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_520),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_537),
.B(n_447),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_537),
.B(n_450),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_520),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_197),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_520),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_502),
.B(n_457),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_520),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_526),
.B(n_366),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_512),
.B(n_459),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_523),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_502),
.B(n_460),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_541),
.A2(n_484),
.B1(n_485),
.B2(n_290),
.Y(n_659)
);

INVx8_ASAP7_75t_L g660 ( 
.A(n_508),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_553),
.B(n_508),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_505),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_553),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_512),
.B(n_462),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_513),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_496),
.B(n_465),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_515),
.B(n_466),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_523),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_515),
.B(n_467),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_523),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

NAND2xp33_ASAP7_75t_SL g674 ( 
.A(n_496),
.B(n_476),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_523),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_566),
.B(n_481),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_523),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_502),
.B(n_490),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_566),
.B(n_311),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_523),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_541),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_536),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_502),
.B(n_311),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_557),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_547),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_557),
.B(n_311),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_SL g690 ( 
.A(n_499),
.B(n_284),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_541),
.A2(n_338),
.B1(n_364),
.B2(n_335),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_508),
.B(n_429),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_536),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_557),
.B(n_508),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_557),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_438),
.Y(n_697)
);

XNOR2x2_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_218),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_536),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_548),
.B(n_499),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_506),
.B(n_438),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_506),
.B(n_330),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_536),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_504),
.B(n_377),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_510),
.B(n_438),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_526),
.B(n_366),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_567),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_532),
.A2(n_289),
.B1(n_303),
.B2(n_287),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_567),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_548),
.B(n_306),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_567),
.B(n_242),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_567),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_541),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_510),
.B(n_348),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_548),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_548),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_567),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_505),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_493),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_667),
.B(n_517),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_593),
.B(n_548),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_620),
.A2(n_511),
.B1(n_535),
.B2(n_491),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_590),
.B(n_517),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_601),
.A2(n_532),
.B1(n_494),
.B2(n_569),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_575),
.B(n_586),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_663),
.B(n_519),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_604),
.B(n_500),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_631),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_578),
.A2(n_494),
.B1(n_504),
.B2(n_519),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_627),
.B(n_522),
.C(n_521),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_571),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_663),
.B(n_521),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_616),
.B(n_522),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_616),
.B(n_591),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_578),
.B(n_525),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_597),
.A2(n_569),
.B1(n_565),
.B2(n_564),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_631),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_578),
.B(n_601),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_631),
.B(n_525),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_634),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_576),
.A2(n_565),
.B1(n_564),
.B2(n_563),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_660),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_634),
.B(n_527),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_621),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_582),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_634),
.B(n_527),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_591),
.A2(n_528),
.B(n_546),
.C(n_526),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_665),
.B(n_529),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_692),
.A2(n_554),
.B1(n_562),
.B2(n_561),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_685),
.B(n_529),
.Y(n_754)
);

AND2x6_ASAP7_75t_SL g755 ( 
.A(n_698),
.B(n_228),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_607),
.B(n_500),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_685),
.B(n_531),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_685),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_698),
.A2(n_563),
.B1(n_562),
.B2(n_561),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_616),
.B(n_531),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_616),
.B(n_591),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_579),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_579),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_668),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_580),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_580),
.Y(n_766)
);

BUFx6f_ASAP7_75t_SL g767 ( 
.A(n_591),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_577),
.B(n_533),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_668),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_596),
.B(n_533),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_717),
.B(n_560),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_623),
.B(n_643),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_696),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_617),
.A2(n_539),
.B1(n_559),
.B2(n_558),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_584),
.B(n_534),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_702),
.A2(n_492),
.B(n_559),
.C(n_558),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_696),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_534),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_615),
.B(n_539),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_716),
.B(n_540),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_640),
.B(n_540),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_652),
.B(n_543),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_704),
.A2(n_377),
.B1(n_555),
.B2(n_491),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_696),
.B(n_543),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_581),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_584),
.B(n_545),
.Y(n_786)
);

AOI22x1_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_687),
.B1(n_603),
.B2(n_672),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_658),
.B(n_545),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_678),
.B(n_619),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_632),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_600),
.B(n_554),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_615),
.B(n_528),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_717),
.B(n_500),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_647),
.B(n_511),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_576),
.A2(n_555),
.B1(n_535),
.B2(n_546),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_719),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_615),
.B(n_528),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_615),
.B(n_528),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_581),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_546),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_719),
.B(n_524),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_SL g802 ( 
.A1(n_662),
.A2(n_316),
.B1(n_314),
.B2(n_388),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_661),
.B(n_524),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_626),
.B(n_546),
.Y(n_804)
);

INVx8_ASAP7_75t_L g805 ( 
.A(n_660),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_626),
.B(n_689),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_626),
.B(n_524),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_598),
.B(n_538),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_660),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_538),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_625),
.B(n_538),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_635),
.A2(n_492),
.B(n_542),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_625),
.B(n_542),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_648),
.B(n_542),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_626),
.B(n_560),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_689),
.B(n_560),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_645),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_693),
.B(n_700),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_693),
.B(n_492),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_674),
.A2(n_383),
.B1(n_374),
.B2(n_369),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_592),
.B(n_325),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_618),
.B(n_292),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_689),
.B(n_367),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_583),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_588),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_659),
.A2(n_377),
.B1(n_242),
.B2(n_300),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_588),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_689),
.B(n_367),
.Y(n_830)
);

BUFx8_ASAP7_75t_L g831 ( 
.A(n_641),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_695),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_636),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_641),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_620),
.B(n_333),
.C(n_327),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_598),
.B(n_228),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_636),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_689),
.B(n_369),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_660),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_660),
.Y(n_840)
);

BUFx5_ASAP7_75t_L g841 ( 
.A(n_650),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_621),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_621),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_681),
.B(n_320),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_574),
.B(n_264),
.C(n_261),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_681),
.B(n_374),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_572),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_645),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_715),
.B(n_375),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_715),
.B(n_375),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_638),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_707),
.B(n_383),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_655),
.B(n_334),
.Y(n_853)
);

AOI221xp5_ASAP7_75t_L g854 ( 
.A1(n_676),
.A2(n_338),
.B1(n_290),
.B2(n_281),
.C(n_335),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_606),
.B(n_345),
.C(n_337),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_707),
.B(n_635),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_664),
.B(n_346),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_683),
.B(n_385),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_712),
.A2(n_354),
.B(n_362),
.C(n_273),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_385),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_654),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_669),
.B(n_349),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_599),
.B(n_273),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_671),
.B(n_281),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_679),
.B(n_355),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_709),
.B(n_624),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_638),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_721),
.A2(n_360),
.B1(n_362),
.B2(n_321),
.C(n_364),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_690),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_707),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_707),
.B(n_198),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_624),
.B(n_357),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_599),
.B(n_298),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_642),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_599),
.B(n_298),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_707),
.B(n_248),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_599),
.B(n_319),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_572),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_603),
.B(n_319),
.Y(n_879)
);

O2A1O1Ixp5_ASAP7_75t_L g880 ( 
.A1(n_714),
.A2(n_360),
.B(n_368),
.C(n_321),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_642),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_714),
.A2(n_493),
.B(n_304),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_686),
.A2(n_368),
.B1(n_361),
.B2(n_371),
.C(n_384),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_587),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_587),
.A2(n_304),
.B(n_296),
.C(n_265),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_714),
.B(n_265),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_603),
.B(n_358),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_603),
.B(n_372),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_654),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_624),
.B(n_296),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_672),
.B(n_687),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_814),
.A2(n_602),
.B(n_589),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_789),
.A2(n_697),
.B(n_602),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_741),
.A2(n_672),
.B(n_610),
.C(n_718),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_723),
.B(n_687),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_767),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_821),
.A2(n_605),
.B(n_589),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_856),
.A2(n_705),
.B(n_701),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_891),
.A2(n_806),
.B(n_782),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_806),
.A2(n_608),
.B(n_605),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_781),
.A2(n_609),
.B(n_608),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_745),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_832),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_726),
.B(n_687),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_805),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_745),
.B(n_573),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_788),
.A2(n_611),
.B(n_609),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_734),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_741),
.A2(n_672),
.B1(n_720),
.B2(n_612),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_803),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_750),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_840),
.B(n_594),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_767),
.B(n_585),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_812),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_770),
.A2(n_611),
.B(n_720),
.C(n_612),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_745),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_794),
.B(n_594),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_778),
.A2(n_670),
.B(n_628),
.C(n_629),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_725),
.B(n_594),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_737),
.B(n_595),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_831),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_769),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_853),
.B(n_380),
.C(n_373),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_SL g924 ( 
.A1(n_728),
.A2(n_628),
.B(n_629),
.C(n_633),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_761),
.B(n_595),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_776),
.A2(n_614),
.B(n_613),
.Y(n_926)
);

BUFx4f_ASAP7_75t_L g927 ( 
.A(n_805),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_815),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_809),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_857),
.A2(n_381),
.B(n_613),
.Y(n_930)
);

AND2x4_ASAP7_75t_SL g931 ( 
.A(n_752),
.B(n_377),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_783),
.A2(n_670),
.B1(n_633),
.B2(n_637),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_856),
.A2(n_637),
.B(n_614),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_780),
.B(n_595),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_738),
.A2(n_673),
.B(n_639),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_835),
.B(n_722),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_820),
.B(n_722),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_808),
.B(n_610),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_792),
.A2(n_673),
.B(n_639),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_790),
.A2(n_751),
.B(n_792),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_796),
.A2(n_760),
.B1(n_736),
.B2(n_866),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_745),
.B(n_610),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_724),
.B(n_654),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_730),
.B(n_759),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_810),
.B(n_722),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_729),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_772),
.B(n_722),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_775),
.B(n_622),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_797),
.A2(n_684),
.B(n_680),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_810),
.B(n_573),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_786),
.B(n_654),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_797),
.A2(n_684),
.B(n_680),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_798),
.A2(n_699),
.B(n_691),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_810),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_861),
.B(n_644),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_791),
.A2(n_691),
.B1(n_699),
.B2(n_710),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_768),
.A2(n_718),
.B(n_622),
.C(n_711),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_748),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_839),
.B(n_573),
.Y(n_961)
);

NAND3xp33_ASAP7_75t_SL g962 ( 
.A(n_862),
.B(n_203),
.C(n_202),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_798),
.A2(n_804),
.B(n_807),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_804),
.A2(n_818),
.B(n_807),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_839),
.A2(n_733),
.B1(n_771),
.B2(n_777),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_818),
.A2(n_703),
.B(n_708),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_865),
.A2(n_703),
.B1(n_710),
.B2(n_708),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_764),
.B(n_644),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_750),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_732),
.B(n_622),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_834),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_816),
.B(n_630),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_742),
.A2(n_649),
.B(n_651),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_869),
.B(n_649),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_756),
.B(n_630),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_742),
.A2(n_651),
.B(n_675),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_746),
.A2(n_675),
.B(n_677),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_831),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_828),
.B(n_242),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_831),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_839),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_839),
.B(n_573),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_836),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_735),
.B(n_630),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_751),
.A2(n_677),
.B(n_682),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_863),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_738),
.A2(n_682),
.B(n_694),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_746),
.A2(n_694),
.B(n_657),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_848),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_771),
.A2(n_711),
.B1(n_666),
.B2(n_657),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_749),
.A2(n_718),
.B(n_657),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_855),
.B(n_646),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_749),
.A2(n_757),
.B(n_754),
.Y(n_993)
);

O2A1O1Ixp5_ASAP7_75t_L g994 ( 
.A1(n_795),
.A2(n_646),
.B(n_711),
.C(n_653),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_873),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_754),
.A2(n_666),
.B(n_656),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_844),
.B(n_646),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_889),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_747),
.Y(n_999)
);

OAI321xp33_ASAP7_75t_L g1000 ( 
.A1(n_868),
.A2(n_300),
.A3(n_493),
.B1(n_666),
.B2(n_653),
.C(n_656),
.Y(n_1000)
);

AO21x1_ASAP7_75t_L g1001 ( 
.A1(n_886),
.A2(n_656),
.B(n_653),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_824),
.B(n_654),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_739),
.B(n_654),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_889),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_822),
.B(n_573),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_757),
.A2(n_573),
.B(n_713),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_774),
.B(n_654),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_784),
.A2(n_210),
.B(n_207),
.Y(n_1008)
);

NOR2x2_ASAP7_75t_L g1009 ( 
.A(n_755),
.B(n_16),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_727),
.B(n_706),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_753),
.B(n_864),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_747),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_819),
.B(n_706),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_777),
.A2(n_300),
.B1(n_275),
.B2(n_279),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_870),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_861),
.Y(n_1016)
);

NAND2x1p5_ASAP7_75t_L g1017 ( 
.A(n_870),
.B(n_493),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_706),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_823),
.B(n_793),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_801),
.B(n_706),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_870),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_784),
.A2(n_212),
.B(n_206),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_845),
.B(n_211),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_785),
.A2(n_214),
.B(n_226),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_731),
.B(n_706),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_802),
.Y(n_1026)
);

O2A1O1Ixp5_ASAP7_75t_L g1027 ( 
.A1(n_744),
.A2(n_880),
.B(n_890),
.C(n_871),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_870),
.B(n_222),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_875),
.A2(n_305),
.B(n_293),
.C(n_279),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_740),
.B(n_706),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_841),
.B(n_300),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_886),
.A2(n_650),
.B(n_706),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_785),
.A2(n_230),
.B(n_253),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_861),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_743),
.B(n_20),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_883),
.B(n_305),
.C(n_247),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_877),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_799),
.A2(n_309),
.B(n_241),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_758),
.B(n_650),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_847),
.A2(n_650),
.B(n_312),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_841),
.B(n_300),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_889),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_799),
.A2(n_315),
.B(n_243),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_854),
.B(n_650),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_879),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_813),
.A2(n_317),
.B(n_246),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_773),
.B(n_650),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_841),
.B(n_300),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_842),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_887),
.A2(n_293),
.B(n_279),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_878),
.A2(n_650),
.B(n_336),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_843),
.B(n_22),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_762),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_888),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_825),
.B(n_438),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_846),
.B(n_233),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_859),
.B(n_252),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_825),
.B(n_247),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_884),
.A2(n_340),
.B(n_389),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_849),
.B(n_850),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_813),
.A2(n_331),
.B(n_387),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_826),
.A2(n_342),
.B(n_379),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_890),
.A2(n_493),
.B(n_23),
.C(n_24),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_858),
.B(n_257),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_841),
.B(n_493),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_860),
.B(n_259),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_763),
.B(n_765),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_765),
.B(n_493),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_830),
.A2(n_378),
.B(n_376),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_841),
.B(n_291),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_826),
.A2(n_363),
.B(n_356),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_766),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_827),
.B(n_22),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_766),
.B(n_353),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_827),
.B(n_352),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_829),
.A2(n_351),
.B(n_262),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_833),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_983),
.B(n_971),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1042),
.B(n_833),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_960),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_923),
.A2(n_852),
.B(n_838),
.C(n_830),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_947),
.B(n_837),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_957),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_949),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_994),
.A2(n_837),
.B(n_881),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_922),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_921),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_929),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_979),
.B(n_841),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_949),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1016),
.B(n_851),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1042),
.B(n_851),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_914),
.B(n_867),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_928),
.B(n_867),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1016),
.B(n_874),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_971),
.B(n_838),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_904),
.A2(n_800),
.B(n_811),
.Y(n_1097)
);

INVx8_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1053),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_904),
.A2(n_817),
.B(n_779),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_927),
.B(n_841),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_910),
.B(n_874),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_978),
.B(n_852),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1016),
.B(n_881),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_896),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_931),
.B(n_871),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1011),
.B(n_876),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_927),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1018),
.A2(n_787),
.B(n_876),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_979),
.A2(n_882),
.B(n_24),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_895),
.A2(n_885),
.B(n_297),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_892),
.A2(n_343),
.B(n_291),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1026),
.B(n_989),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_942),
.A2(n_301),
.B(n_299),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_953),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_899),
.A2(n_295),
.B(n_285),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_913),
.B(n_23),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_939),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_903),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1015),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_934),
.A2(n_277),
.B(n_343),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_939),
.B(n_343),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1019),
.B(n_25),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1054),
.B(n_26),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1072),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_897),
.A2(n_343),
.B(n_291),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_896),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_917),
.A2(n_343),
.B(n_291),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_980),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1077),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1013),
.B(n_1023),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_923),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1132)
);

OAI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_962),
.A2(n_343),
.B(n_291),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_962),
.A2(n_291),
.B1(n_33),
.B2(n_36),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_893),
.A2(n_179),
.B(n_168),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_905),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_919),
.A2(n_166),
.B(n_160),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_905),
.B(n_27),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_932),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1036),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_948),
.B(n_43),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1003),
.A2(n_950),
.B1(n_948),
.B2(n_1010),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1015),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_913),
.B(n_45),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_978),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_968),
.B(n_45),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_958),
.A2(n_77),
.B(n_151),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_944),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_998),
.B(n_76),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1004),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_902),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_943),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_926),
.A2(n_153),
.B(n_150),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1036),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_986),
.B(n_995),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1035),
.A2(n_945),
.B1(n_1052),
.B2(n_938),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_46),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1058),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_902),
.B(n_101),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_994),
.A2(n_49),
.B(n_50),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1015),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_999),
.B(n_52),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1035),
.B(n_54),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_984),
.A2(n_95),
.B(n_133),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1037),
.B(n_57),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1045),
.B(n_62),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_908),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_902),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1044),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1073),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_936),
.A2(n_67),
.B(n_68),
.C(n_70),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1058),
.B(n_73),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_1009),
.A2(n_74),
.B1(n_91),
.B2(n_98),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_999),
.B(n_99),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1016),
.B(n_106),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_911),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_943),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_937),
.B(n_113),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_969),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1049),
.Y(n_1181)
);

INVx3_ASAP7_75t_SL g1182 ( 
.A(n_957),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_937),
.B(n_118),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1034),
.B(n_148),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_902),
.B(n_916),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1034),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_1052),
.B(n_1073),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_L g1188 ( 
.A1(n_1028),
.A2(n_1027),
.B(n_1040),
.C(n_1051),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_924),
.A2(n_963),
.B(n_964),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1057),
.A2(n_918),
.B(n_915),
.C(n_959),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_967),
.A2(n_1007),
.B1(n_925),
.B2(n_920),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1034),
.B(n_916),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1063),
.B(n_965),
.C(n_1027),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_SL g1194 ( 
.A(n_930),
.B(n_1066),
.C(n_1064),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1049),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1012),
.B(n_974),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_936),
.A2(n_974),
.B(n_941),
.C(n_1002),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1069),
.B(n_1008),
.C(n_1022),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_912),
.A2(n_1056),
.B1(n_1012),
.B2(n_1005),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_901),
.A2(n_907),
.B(n_933),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_916),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1060),
.B(n_970),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1049),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1074),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_909),
.A2(n_1020),
.B1(n_993),
.B2(n_1025),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_916),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1049),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_894),
.A2(n_996),
.B(n_991),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1067),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_R g1210 ( 
.A(n_956),
.B(n_981),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_900),
.A2(n_988),
.B(n_976),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_975),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1034),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1030),
.A2(n_912),
.B1(n_972),
.B2(n_981),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_956),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1021),
.B(n_1075),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1021),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_935),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1068),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_992),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1039),
.A2(n_1047),
.B(n_1038),
.C(n_1076),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_997),
.B(n_956),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_956),
.B(n_981),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_981),
.B(n_1000),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_990),
.B(n_906),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1001),
.A2(n_985),
.B(n_987),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1024),
.B(n_1071),
.C(n_1062),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_946),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_906),
.B(n_1017),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_973),
.A2(n_977),
.B(n_940),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1017),
.A2(n_961),
.B1(n_952),
.B2(n_982),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1055),
.B(n_1065),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_951),
.A2(n_954),
.B(n_955),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1055),
.B(n_1065),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1050),
.A2(n_1014),
.B1(n_1061),
.B2(n_1046),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1029),
.B(n_1043),
.C(n_1033),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1113),
.B(n_1032),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1156),
.B(n_1123),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1179),
.A2(n_966),
.B(n_1070),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1139),
.A2(n_1006),
.B1(n_1031),
.B2(n_1041),
.C(n_1048),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1084),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1086),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1078),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1112),
.A2(n_898),
.B(n_1031),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1183),
.A2(n_1070),
.B(n_1041),
.Y(n_1245)
);

NAND3x1_ASAP7_75t_L g1246 ( 
.A(n_1144),
.B(n_1048),
.C(n_1170),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1089),
.A2(n_1140),
.B1(n_1134),
.B2(n_1139),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1164),
.A2(n_1159),
.B1(n_1158),
.B2(n_1124),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1156),
.B(n_1171),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1130),
.B(n_1096),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1189),
.A2(n_1208),
.B(n_1230),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_SL g1252 ( 
.A(n_1083),
.B(n_1186),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_1196),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1204),
.B(n_1202),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_1157),
.A2(n_1115),
.B1(n_1142),
.B2(n_1218),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_SL g1256 ( 
.A(n_1083),
.B(n_1186),
.Y(n_1256)
);

A2O1A1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1089),
.A2(n_1133),
.B(n_1157),
.C(n_1110),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1097),
.A2(n_1100),
.B(n_1197),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1142),
.A2(n_1191),
.A3(n_1126),
.B(n_1205),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1200),
.A2(n_1211),
.B(n_1109),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1141),
.A2(n_1146),
.B1(n_1115),
.B2(n_1081),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1233),
.A2(n_1085),
.B(n_1205),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1225),
.A2(n_1191),
.B(n_1085),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1161),
.A2(n_1188),
.B(n_1128),
.Y(n_1264)
);

O2A1O1Ixp5_ASAP7_75t_L g1265 ( 
.A1(n_1141),
.A2(n_1161),
.B(n_1147),
.C(n_1154),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1135),
.A2(n_1221),
.B(n_1214),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1193),
.A2(n_1190),
.B(n_1224),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1088),
.B(n_1119),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1194),
.A2(n_1121),
.B(n_1111),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1166),
.A2(n_1167),
.B1(n_1199),
.B2(n_1172),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1125),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1132),
.A2(n_1155),
.B(n_1138),
.C(n_1117),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1137),
.A2(n_1229),
.B(n_1175),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1214),
.A2(n_1220),
.A3(n_1107),
.B(n_1212),
.Y(n_1274)
);

OAI22x1_ASAP7_75t_L g1275 ( 
.A1(n_1131),
.A2(n_1106),
.B1(n_1173),
.B2(n_1127),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1168),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1108),
.B(n_1178),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1084),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1231),
.A2(n_1165),
.B(n_1094),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1084),
.B(n_1090),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1231),
.A2(n_1093),
.B(n_1094),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1148),
.A2(n_1174),
.B1(n_1163),
.B2(n_1103),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1105),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1093),
.A2(n_1222),
.B(n_1216),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1145),
.B(n_1150),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1080),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1114),
.A2(n_1176),
.B(n_1116),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1177),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1101),
.A2(n_1185),
.B(n_1223),
.C(n_1122),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1226),
.A2(n_1091),
.B(n_1235),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1198),
.A2(n_1082),
.B(n_1227),
.C(n_1079),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1180),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1118),
.A2(n_1136),
.B1(n_1182),
.B2(n_1153),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1102),
.A2(n_1223),
.B(n_1209),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1219),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1079),
.A2(n_1092),
.B(n_1207),
.C(n_1234),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1091),
.A2(n_1215),
.B(n_1213),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1099),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1232),
.A2(n_1234),
.B(n_1092),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1232),
.A2(n_1203),
.B(n_1181),
.C(n_1195),
.Y(n_1300)
);

OAI22x1_ASAP7_75t_L g1301 ( 
.A1(n_1129),
.A2(n_1087),
.B1(n_1153),
.B2(n_1184),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1184),
.A2(n_1090),
.B1(n_1098),
.B2(n_1217),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1210),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1095),
.A2(n_1104),
.B(n_1098),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1090),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1098),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1118),
.B(n_1083),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1151),
.A2(n_1192),
.B1(n_1095),
.B2(n_1104),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1169),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1186),
.B(n_1192),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1136),
.A2(n_1083),
.B(n_1120),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1186),
.A2(n_1206),
.B1(n_1201),
.B2(n_1120),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1149),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1143),
.B(n_1152),
.Y(n_1314)
);

AO32x2_ASAP7_75t_L g1315 ( 
.A1(n_1160),
.A2(n_1143),
.A3(n_1152),
.B1(n_1162),
.B2(n_1201),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1152),
.B(n_1162),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1228),
.A2(n_1162),
.B1(n_1201),
.B2(n_1206),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1228),
.A2(n_1112),
.B(n_1189),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1206),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1228),
.A2(n_1187),
.B1(n_1158),
.B2(n_1141),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1118),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1119),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1156),
.B(n_752),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1187),
.A2(n_1158),
.B(n_1123),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1156),
.B(n_752),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1084),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1119),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1086),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1119),
.Y(n_1330)
);

AO32x2_ASAP7_75t_L g1331 ( 
.A1(n_1139),
.A2(n_1142),
.A3(n_1157),
.B1(n_1191),
.B2(n_1205),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1187),
.B(n_1158),
.C(n_923),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1156),
.B(n_752),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1118),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1156),
.B(n_752),
.Y(n_1335)
);

AO21x1_ASAP7_75t_L g1336 ( 
.A1(n_1089),
.A2(n_1157),
.B(n_1139),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1187),
.A2(n_1123),
.B(n_923),
.C(n_1158),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1119),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1218),
.A2(n_1001),
.A3(n_1142),
.B(n_1197),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1112),
.A2(n_1189),
.B(n_1208),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1218),
.A2(n_1001),
.A3(n_1142),
.B(n_1197),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1080),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1089),
.A2(n_1157),
.B(n_1139),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1187),
.A2(n_530),
.B1(n_556),
.B2(n_404),
.C(n_574),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1119),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1112),
.A2(n_1189),
.B(n_1208),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1157),
.B(n_593),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1087),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1158),
.A2(n_1187),
.B1(n_1089),
.B2(n_1123),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1204),
.B(n_582),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1084),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1118),
.B(n_1108),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1080),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1156),
.B(n_752),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1119),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1084),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1084),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1187),
.A2(n_1123),
.B(n_923),
.C(n_1158),
.Y(n_1359)
);

OAI22x1_ASAP7_75t_L g1360 ( 
.A1(n_1170),
.A2(n_620),
.B1(n_547),
.B2(n_1134),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1112),
.A2(n_1189),
.B(n_1208),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1119),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1139),
.A2(n_1187),
.B1(n_1133),
.B2(n_1193),
.C(n_1161),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1204),
.B(n_582),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1187),
.A2(n_1158),
.B(n_1123),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1080),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1156),
.B(n_752),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1139),
.A2(n_1187),
.B1(n_601),
.B2(n_1132),
.C(n_1155),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1084),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1118),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1187),
.A2(n_1158),
.B(n_1123),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1373)
);

NAND2xp33_ASAP7_75t_SL g1374 ( 
.A(n_1118),
.B(n_905),
.Y(n_1374)
);

AOI31xp67_ASAP7_75t_L g1375 ( 
.A1(n_1225),
.A2(n_1229),
.A3(n_1183),
.B(n_1179),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1112),
.A2(n_1189),
.B(n_1208),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1187),
.A2(n_1158),
.B(n_1123),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1086),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1119),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1218),
.A2(n_1001),
.A3(n_1142),
.B(n_1197),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1139),
.A2(n_1187),
.B1(n_601),
.B2(n_1132),
.C(n_1155),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1187),
.A2(n_1018),
.B(n_1179),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1089),
.A2(n_620),
.B1(n_704),
.B2(n_1140),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1078),
.B(n_769),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1156),
.B(n_752),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1112),
.A2(n_1189),
.B(n_1208),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1158),
.A2(n_1187),
.B1(n_1089),
.B2(n_1123),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1324),
.A2(n_1372),
.B(n_1365),
.Y(n_1393)
);

AOI21xp33_ASAP7_75t_L g1394 ( 
.A1(n_1377),
.A2(n_1332),
.B(n_1337),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1366),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1342),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1348),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1360),
.A2(n_1388),
.B1(n_1332),
.B2(n_1336),
.Y(n_1398)
);

INVx3_ASAP7_75t_SL g1399 ( 
.A(n_1353),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1285),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1322),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1359),
.A2(n_1392),
.B1(n_1349),
.B2(n_1282),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1282),
.A2(n_1392),
.B1(n_1349),
.B2(n_1238),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1389),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1381),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1328),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1344),
.A2(n_1272),
.B(n_1247),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1343),
.A2(n_1347),
.B1(n_1248),
.B2(n_1261),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1363),
.A2(n_1354),
.B1(n_1325),
.B2(n_1367),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1303),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1307),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1303),
.Y(n_1412)
);

BUFx10_ASAP7_75t_L g1413 ( 
.A(n_1350),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1330),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1242),
.Y(n_1416)
);

AOI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1270),
.A2(n_1386),
.B(n_1368),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1338),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1323),
.A2(n_1390),
.B1(n_1333),
.B2(n_1335),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1253),
.A2(n_1320),
.B1(n_1257),
.B2(n_1267),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1265),
.A2(n_1327),
.B(n_1387),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1255),
.A2(n_1275),
.B1(n_1301),
.B2(n_1295),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1255),
.A2(n_1263),
.B1(n_1384),
.B2(n_1355),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1339),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1286),
.A2(n_1283),
.B1(n_1364),
.B2(n_1246),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1306),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1250),
.A2(n_1302),
.B1(n_1345),
.B2(n_1362),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1313),
.A2(n_1329),
.B1(n_1237),
.B2(n_1368),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_1352),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1319),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1243),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1241),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1386),
.A2(n_1299),
.B1(n_1331),
.B2(n_1277),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1241),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1299),
.A2(n_1331),
.B1(n_1288),
.B2(n_1276),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1278),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1326),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1271),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1278),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1284),
.B(n_1292),
.Y(n_1440)
);

INVx6_ASAP7_75t_L g1441 ( 
.A(n_1326),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1351),
.Y(n_1442)
);

CKINVDCx6p67_ASAP7_75t_R g1443 ( 
.A(n_1278),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1315),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1321),
.A2(n_1334),
.B1(n_1370),
.B2(n_1302),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1298),
.A2(n_1378),
.B1(n_1371),
.B2(n_1373),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1331),
.A2(n_1281),
.B1(n_1382),
.B2(n_1358),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1305),
.Y(n_1448)
);

NAND2x1p5_ASAP7_75t_L g1449 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1379),
.A2(n_1380),
.B1(n_1383),
.B2(n_1294),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1309),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1305),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1315),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1287),
.A2(n_1293),
.B1(n_1264),
.B2(n_1279),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1356),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1240),
.A2(n_1308),
.B1(n_1334),
.B2(n_1321),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1252),
.A2(n_1256),
.B1(n_1264),
.B2(n_1273),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1356),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1274),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1357),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1357),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1304),
.A2(n_1369),
.B1(n_1280),
.B2(n_1308),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1369),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1311),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1269),
.A2(n_1245),
.B1(n_1258),
.B2(n_1266),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1262),
.A2(n_1239),
.B1(n_1374),
.B2(n_1316),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1314),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1290),
.A2(n_1312),
.B1(n_1317),
.B2(n_1260),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1259),
.A2(n_1297),
.B1(n_1375),
.B2(n_1251),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1300),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1259),
.A2(n_1244),
.B1(n_1318),
.B2(n_1376),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1289),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1259),
.A2(n_1391),
.B1(n_1361),
.B2(n_1346),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1340),
.A2(n_1296),
.B1(n_1341),
.B2(n_1385),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1291),
.A2(n_1236),
.B1(n_1341),
.B2(n_1385),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1385),
.A2(n_698),
.B1(n_1360),
.B2(n_549),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1339),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1332),
.A2(n_645),
.B1(n_698),
.B2(n_704),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1282),
.A2(n_704),
.B1(n_1347),
.B2(n_1238),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1324),
.A2(n_1372),
.B(n_1365),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1332),
.A2(n_645),
.B1(n_698),
.B2(n_704),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1353),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1342),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1342),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1315),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1268),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1238),
.B(n_1249),
.Y(n_1490)
);

BUFx8_ASAP7_75t_SL g1491 ( 
.A(n_1348),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1332),
.A2(n_645),
.B1(n_698),
.B2(n_704),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1268),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1324),
.A2(n_1372),
.B(n_1365),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1332),
.A2(n_645),
.B1(n_698),
.B2(n_704),
.Y(n_1495)
);

BUFx12f_ASAP7_75t_L g1496 ( 
.A(n_1366),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1337),
.A2(n_1359),
.B1(n_1332),
.B2(n_1324),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1366),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1337),
.A2(n_1359),
.B1(n_1332),
.B2(n_1324),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1282),
.A2(n_704),
.B1(n_1347),
.B2(n_1238),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1268),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1243),
.B(n_1253),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1306),
.B(n_1299),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1268),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1342),
.Y(n_1507)
);

CKINVDCx6p67_ASAP7_75t_R g1508 ( 
.A(n_1366),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1238),
.B(n_1249),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1360),
.A2(n_698),
.B1(n_549),
.B2(n_1324),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1360),
.A2(n_1248),
.B1(n_582),
.B2(n_1301),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1282),
.A2(n_1089),
.B1(n_1392),
.B2(n_1349),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1238),
.B(n_1249),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1366),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1238),
.B(n_1249),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1285),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1348),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1353),
.Y(n_1519)
);

CKINVDCx14_ASAP7_75t_R g1520 ( 
.A(n_1366),
.Y(n_1520)
);

INVx4_ASAP7_75t_L g1521 ( 
.A(n_1353),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1444),
.B(n_1453),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1400),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1421),
.A2(n_1465),
.B(n_1454),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1440),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1407),
.A2(n_1499),
.B(n_1497),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1478),
.A2(n_1495),
.B1(n_1492),
.B2(n_1482),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1427),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1459),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1424),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1504),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1477),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1477),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1491),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1486),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1465),
.A2(n_1473),
.B(n_1454),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1513),
.A2(n_1447),
.B(n_1403),
.Y(n_1538)
);

CKINVDCx14_ASAP7_75t_R g1539 ( 
.A(n_1520),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1414),
.B(n_1418),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1438),
.B(n_1433),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1464),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1505),
.B(n_1402),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1451),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1449),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1464),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1395),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1490),
.B(n_1509),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1423),
.B(n_1435),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1423),
.B(n_1398),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1470),
.B(n_1449),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1450),
.A2(n_1473),
.B(n_1469),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1430),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1394),
.A2(n_1393),
.B(n_1494),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1447),
.A2(n_1417),
.B(n_1450),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1471),
.A2(n_1469),
.B(n_1446),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1558)
);

AND2x2_ASAP7_75t_SL g1559 ( 
.A(n_1398),
.B(n_1408),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1472),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1420),
.A2(n_1445),
.B(n_1425),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1475),
.B(n_1474),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1487),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1472),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1493),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1503),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1506),
.B(n_1408),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1429),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1446),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1427),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1468),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1468),
.Y(n_1572)
);

AOI21xp33_ASAP7_75t_L g1573 ( 
.A1(n_1513),
.A2(n_1403),
.B(n_1479),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1500),
.B(n_1409),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1485),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1485),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1467),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1409),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1471),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1480),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1466),
.Y(n_1581)
);

INVx3_ASAP7_75t_SL g1582 ( 
.A(n_1443),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1466),
.Y(n_1584)
);

BUFx12f_ASAP7_75t_L g1585 ( 
.A(n_1412),
.Y(n_1585)
);

BUFx4f_ASAP7_75t_SL g1586 ( 
.A(n_1496),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1422),
.A2(n_1462),
.B(n_1411),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1456),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1515),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1422),
.A2(n_1462),
.B(n_1411),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1476),
.B(n_1428),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1456),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1457),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1419),
.B(n_1415),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1426),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1481),
.A2(n_1489),
.B(n_1488),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1481),
.A2(n_1489),
.B(n_1488),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1501),
.A2(n_1511),
.B1(n_1502),
.B2(n_1510),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1484),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1512),
.B(n_1404),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1501),
.A2(n_1511),
.B1(n_1510),
.B2(n_1502),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1405),
.B(n_1452),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1410),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1518),
.B(n_1396),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1432),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1507),
.B(n_1413),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1525),
.B(n_1416),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1532),
.B(n_1413),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1545),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1599),
.B(n_1521),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1599),
.B(n_1575),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1526),
.A2(n_1520),
.B1(n_1431),
.B2(n_1397),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1523),
.B(n_1399),
.Y(n_1614)
);

INVx6_ASAP7_75t_L g1615 ( 
.A(n_1605),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1585),
.Y(n_1616)
);

OR2x6_ASAP7_75t_L g1617 ( 
.A(n_1544),
.B(n_1460),
.Y(n_1617)
);

AOI221x1_ASAP7_75t_L g1618 ( 
.A1(n_1526),
.A2(n_1519),
.B1(n_1483),
.B2(n_1460),
.C(n_1458),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1576),
.B(n_1483),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1602),
.Y(n_1620)
);

AOI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1598),
.A2(n_1455),
.B1(n_1439),
.B2(n_1434),
.C(n_1448),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1399),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1525),
.B(n_1397),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1602),
.B(n_1508),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1555),
.A2(n_1498),
.B(n_1461),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1555),
.A2(n_1528),
.B(n_1573),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1546),
.B(n_1436),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1585),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1601),
.A2(n_1463),
.B(n_1441),
.C(n_1442),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1601),
.A2(n_1437),
.B(n_1441),
.C(n_1442),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1556),
.A2(n_1437),
.B(n_1441),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1578),
.A2(n_1574),
.B1(n_1592),
.B2(n_1588),
.C(n_1580),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1559),
.C(n_1527),
.Y(n_1633)
);

AO32x2_ASAP7_75t_L g1634 ( 
.A1(n_1543),
.A2(n_1547),
.A3(n_1595),
.B1(n_1568),
.B2(n_1522),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1554),
.B(n_1530),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1564),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1530),
.B(n_1541),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1559),
.C(n_1591),
.Y(n_1638)
);

AO32x2_ASAP7_75t_L g1639 ( 
.A1(n_1543),
.A2(n_1547),
.A3(n_1595),
.B1(n_1568),
.B2(n_1522),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1564),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1559),
.A2(n_1591),
.B1(n_1551),
.B2(n_1550),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1573),
.A2(n_1556),
.B(n_1580),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1594),
.B(n_1549),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1551),
.A2(n_1578),
.B(n_1550),
.C(n_1562),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1561),
.A2(n_1570),
.B(n_1569),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1541),
.B(n_1606),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1561),
.A2(n_1570),
.B(n_1569),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1581),
.A2(n_1584),
.B(n_1588),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1606),
.B(n_1603),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1594),
.B(n_1549),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1585),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1544),
.B(n_1552),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1604),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1581),
.A2(n_1584),
.B(n_1592),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1603),
.B(n_1604),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_R g1656 ( 
.A(n_1548),
.B(n_1589),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1535),
.B(n_1539),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1563),
.B(n_1565),
.Y(n_1658)
);

AOI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1562),
.A2(n_1593),
.B(n_1567),
.C(n_1542),
.Y(n_1659)
);

BUFx8_ASAP7_75t_L g1660 ( 
.A(n_1586),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1577),
.B(n_1558),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1538),
.A2(n_1567),
.B1(n_1583),
.B2(n_1542),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1538),
.A2(n_1583),
.B1(n_1544),
.B2(n_1572),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1529),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1593),
.A2(n_1600),
.B(n_1587),
.C(n_1590),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1553),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1646),
.B(n_1553),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1537),
.B(n_1557),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1613),
.B(n_1560),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1611),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1666),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1643),
.B(n_1538),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1639),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1634),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1658),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1627),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1658),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1661),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1662),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1661),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1609),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1634),
.B(n_1639),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1639),
.B(n_1553),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1524),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1635),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1655),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1524),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1647),
.B(n_1524),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1641),
.A2(n_1600),
.B1(n_1552),
.B2(n_1579),
.Y(n_1692)
);

BUFx4f_ASAP7_75t_L g1693 ( 
.A(n_1627),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1665),
.B(n_1537),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1631),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1663),
.B(n_1531),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1664),
.B(n_1536),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1665),
.B(n_1537),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1642),
.B(n_1534),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1664),
.B(n_1540),
.Y(n_1700)
);

INVxp67_ASAP7_75t_SL g1701 ( 
.A(n_1631),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1649),
.Y(n_1702)
);

NAND3xp33_ASAP7_75t_L g1703 ( 
.A(n_1699),
.B(n_1632),
.C(n_1659),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1675),
.B(n_1620),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1693),
.Y(n_1705)
);

NAND2x1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.B(n_1636),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1638),
.B1(n_1659),
.B2(n_1633),
.C(n_1644),
.Y(n_1707)
);

NAND5xp2_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1625),
.C(n_1657),
.D(n_1624),
.E(n_1622),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1673),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1684),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1636),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1682),
.B(n_1653),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1679),
.B(n_1617),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1685),
.B(n_1612),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1673),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1672),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1684),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1612),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1695),
.Y(n_1722)
);

AO21x2_ASAP7_75t_L g1723 ( 
.A1(n_1670),
.A2(n_1667),
.B(n_1654),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1670),
.A2(n_1625),
.B1(n_1654),
.B2(n_1648),
.C(n_1613),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1668),
.B(n_1608),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1668),
.B(n_1669),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1673),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1678),
.B(n_1607),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1694),
.A2(n_1621),
.B1(n_1648),
.B2(n_1627),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1693),
.B(n_1640),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1693),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1682),
.B(n_1607),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1693),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_L g1734 ( 
.A(n_1699),
.B(n_1690),
.C(n_1687),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1678),
.B(n_1623),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1669),
.B(n_1623),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1674),
.B(n_1614),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1672),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1692),
.A2(n_1629),
.B1(n_1630),
.B2(n_1652),
.C(n_1628),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1674),
.B(n_1533),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1677),
.B(n_1533),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1726),
.B(n_1676),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1677),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1676),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1717),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1722),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1734),
.B(n_1677),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1737),
.B(n_1696),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1726),
.B(n_1686),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1740),
.B(n_1680),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1686),
.Y(n_1752)
);

NAND2x1_ASAP7_75t_SL g1753 ( 
.A(n_1733),
.B(n_1686),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1703),
.B(n_1671),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

NAND2xp33_ASAP7_75t_R g1756 ( 
.A(n_1731),
.B(n_1616),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1709),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1741),
.B(n_1680),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1741),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1722),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1680),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1709),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1712),
.B(n_1681),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1732),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1733),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1681),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1713),
.B(n_1694),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1716),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1736),
.B(n_1681),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1683),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1722),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1713),
.B(n_1694),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1727),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1757),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1756),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1757),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1766),
.B(n_1728),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1754),
.B(n_1735),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1766),
.B(n_1728),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1717),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1748),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1750),
.B(n_1752),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1766),
.B(n_1732),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1743),
.B(n_1735),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1746),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1748),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1763),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1743),
.B(n_1703),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1746),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1763),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1747),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.B(n_1718),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1749),
.B(n_1718),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1750),
.B(n_1717),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1753),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1801)
);

AOI32xp33_ASAP7_75t_L g1802 ( 
.A1(n_1742),
.A2(n_1724),
.A3(n_1707),
.B1(n_1698),
.B2(n_1700),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1765),
.B(n_1720),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1765),
.B(n_1725),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1752),
.B(n_1725),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1742),
.B(n_1704),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1772),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1749),
.B(n_1738),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1769),
.B(n_1777),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1744),
.B(n_1738),
.Y(n_1810)
);

AOI32xp33_ASAP7_75t_L g1811 ( 
.A1(n_1742),
.A2(n_1724),
.A3(n_1707),
.B1(n_1698),
.B2(n_1700),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1772),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1770),
.B(n_1704),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1759),
.B(n_1689),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1759),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1753),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1770),
.B(n_1704),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1773),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1770),
.B(n_1714),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1778),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1746),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1793),
.B(n_1780),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_SL g1824 ( 
.A(n_1800),
.B(n_1656),
.C(n_1651),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1783),
.B(n_1744),
.Y(n_1826)
);

INVxp67_ASAP7_75t_SL g1827 ( 
.A(n_1796),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1809),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1802),
.B(n_1771),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1809),
.B(n_1771),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1797),
.A2(n_1723),
.B1(n_1698),
.B2(n_1691),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1802),
.B(n_1768),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1782),
.B(n_1768),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1786),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1811),
.A2(n_1708),
.B(n_1761),
.Y(n_1835)
);

OR2x6_ASAP7_75t_L g1836 ( 
.A(n_1810),
.B(n_1767),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1782),
.B(n_1784),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1784),
.B(n_1774),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1789),
.B(n_1798),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1791),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1774),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1797),
.B(n_1775),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1798),
.B(n_1775),
.Y(n_1844)
);

XOR2xp5_ASAP7_75t_L g1845 ( 
.A(n_1810),
.B(n_1729),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1808),
.B(n_1758),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1792),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1803),
.B(n_1708),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1792),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1788),
.B(n_1815),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1788),
.B(n_1751),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1814),
.B(n_1751),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1809),
.B(n_1767),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1785),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1813),
.B(n_1758),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1809),
.B(n_1769),
.Y(n_1856)
);

AOI221x1_ASAP7_75t_L g1857 ( 
.A1(n_1779),
.A2(n_1767),
.B1(n_1761),
.B2(n_1764),
.C(n_1769),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1779),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1806),
.B(n_1767),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1831),
.A2(n_1723),
.B1(n_1729),
.B2(n_1816),
.Y(n_1860)
);

AOI31xp33_ASAP7_75t_SL g1861 ( 
.A1(n_1829),
.A2(n_1804),
.A3(n_1702),
.B(n_1751),
.Y(n_1861)
);

AOI222xp33_ASAP7_75t_L g1862 ( 
.A1(n_1831),
.A2(n_1690),
.B1(n_1691),
.B2(n_1687),
.C1(n_1700),
.C2(n_1806),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1858),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1823),
.B(n_1660),
.Y(n_1864)
);

OAI31xp33_ASAP7_75t_L g1865 ( 
.A1(n_1835),
.A2(n_1739),
.A3(n_1764),
.B(n_1761),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1813),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1832),
.A2(n_1787),
.B1(n_1817),
.B2(n_1777),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1858),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1827),
.B(n_1817),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1827),
.B(n_1801),
.Y(n_1870)
);

NAND3xp33_ASAP7_75t_L g1871 ( 
.A(n_1857),
.B(n_1781),
.C(n_1795),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1845),
.A2(n_1781),
.B(n_1755),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1853),
.B(n_1787),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1837),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1842),
.A2(n_1805),
.B(n_1801),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1847),
.Y(n_1876)
);

OAI32xp33_ASAP7_75t_L g1877 ( 
.A1(n_1848),
.A2(n_1785),
.A3(n_1799),
.B1(n_1739),
.B2(n_1805),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1828),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1828),
.B(n_1799),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1839),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1848),
.A2(n_1723),
.B1(n_1818),
.B2(n_1821),
.C(n_1795),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1824),
.B(n_1820),
.Y(n_1882)
);

OAI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1826),
.A2(n_1697),
.B1(n_1733),
.B2(n_1715),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1850),
.A2(n_1755),
.B(n_1745),
.Y(n_1884)
);

INVxp67_ASAP7_75t_SL g1885 ( 
.A(n_1825),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1833),
.B(n_1762),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1880),
.B(n_1851),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1870),
.B(n_1838),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1879),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1864),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1874),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1860),
.A2(n_1723),
.B1(n_1761),
.B2(n_1764),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1881),
.A2(n_1764),
.B1(n_1761),
.B2(n_1777),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1879),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1866),
.A2(n_1824),
.B1(n_1836),
.B2(n_1843),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1878),
.B(n_1834),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1864),
.B(n_1859),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_L g1898 ( 
.A(n_1865),
.B(n_1872),
.C(n_1871),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1882),
.A2(n_1856),
.B(n_1830),
.Y(n_1899)
);

BUFx2_ASAP7_75t_SL g1900 ( 
.A(n_1878),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1885),
.B(n_1840),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1885),
.B(n_1841),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1869),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1863),
.Y(n_1904)
);

NAND2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1879),
.B(n_1856),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1868),
.Y(n_1906)
);

INVxp67_ASAP7_75t_SL g1907 ( 
.A(n_1901),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1898),
.A2(n_1875),
.B(n_1877),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1887),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1889),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1893),
.A2(n_1892),
.B1(n_1903),
.B2(n_1888),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1905),
.A2(n_1862),
.B1(n_1883),
.B2(n_1867),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1894),
.B(n_1886),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1900),
.B(n_1873),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1896),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1901),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1902),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1902),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1913),
.Y(n_1919)
);

NOR4xp25_ASAP7_75t_L g1920 ( 
.A(n_1908),
.B(n_1906),
.C(n_1890),
.D(n_1904),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1909),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1910),
.Y(n_1922)
);

NAND4xp25_ASAP7_75t_L g1923 ( 
.A(n_1914),
.B(n_1895),
.C(n_1899),
.D(n_1891),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_L g1924 ( 
.A(n_1907),
.B(n_1895),
.C(n_1884),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1915),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1907),
.A2(n_1897),
.B(n_1883),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1912),
.B(n_1856),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1916),
.B(n_1836),
.Y(n_1928)
);

OAI211xp5_ASAP7_75t_SL g1929 ( 
.A1(n_1916),
.A2(n_1861),
.B(n_1876),
.C(n_1854),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1911),
.B(n_1917),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1919),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1929),
.A2(n_1918),
.B(n_1854),
.Y(n_1932)
);

AOI322xp5_ASAP7_75t_L g1933 ( 
.A1(n_1930),
.A2(n_1794),
.A3(n_1849),
.B1(n_1846),
.B2(n_1790),
.C1(n_1822),
.C2(n_1855),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1920),
.A2(n_1836),
.B1(n_1852),
.B2(n_1844),
.C(n_1794),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1921),
.B(n_1820),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_R g1936 ( 
.A(n_1928),
.B(n_1660),
.Y(n_1936)
);

AOI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1932),
.A2(n_1924),
.B1(n_1926),
.B2(n_1922),
.C(n_1925),
.Y(n_1937)
);

OAI33xp33_ASAP7_75t_L g1938 ( 
.A1(n_1931),
.A2(n_1923),
.A3(n_1927),
.B1(n_1807),
.B2(n_1812),
.B3(n_1818),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_SL g1939 ( 
.A(n_1936),
.B(n_1935),
.C(n_1933),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1934),
.A2(n_1821),
.B1(n_1819),
.B2(n_1812),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1931),
.A2(n_1764),
.B1(n_1794),
.B2(n_1790),
.Y(n_1941)
);

AOI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1932),
.A2(n_1582),
.B(n_1819),
.C(n_1807),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1935),
.B(n_1745),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1943),
.Y(n_1944)
);

NAND4xp75_ASAP7_75t_L g1945 ( 
.A(n_1937),
.B(n_1618),
.C(n_1719),
.D(n_1711),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1939),
.Y(n_1946)
);

NOR2xp67_ASAP7_75t_SL g1947 ( 
.A(n_1938),
.B(n_1705),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1941),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1940),
.B(n_1733),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1944),
.B(n_1942),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1946),
.Y(n_1951)
);

OAI211xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1946),
.A2(n_1719),
.B(n_1711),
.C(n_1822),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1947),
.A2(n_1777),
.B1(n_1769),
.B2(n_1760),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1951),
.Y(n_1954)
);

OAI22x1_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1950),
.B1(n_1948),
.B2(n_1949),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1954),
.B1(n_1953),
.B2(n_1945),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1955),
.A2(n_1954),
.B1(n_1952),
.B2(n_1760),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1957),
.B(n_1954),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_1956),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1958),
.Y(n_1960)
);

O2A1O1Ixp33_ASAP7_75t_SL g1961 ( 
.A1(n_1959),
.A2(n_1706),
.B(n_1730),
.C(n_1762),
.Y(n_1961)
);

INVx4_ASAP7_75t_L g1962 ( 
.A(n_1960),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1961),
.B(n_1776),
.Y(n_1963)
);

XOR2xp5_ASAP7_75t_L g1964 ( 
.A(n_1963),
.B(n_1705),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1964),
.A2(n_1582),
.B1(n_1615),
.B2(n_1715),
.C(n_1705),
.Y(n_1965)
);

AOI211xp5_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1582),
.B(n_1610),
.C(n_1619),
.Y(n_1966)
);


endmodule