module fake_netlist_6_1229_n_955 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_955);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_955;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_69),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_21),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_99),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_101),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_17),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_60),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_89),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_38),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_31),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_66),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_88),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_26),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_123),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_70),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_84),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_23),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_85),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_24),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_40),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_21),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_95),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_180),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_54),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_173),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_151),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_53),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_150),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_118),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_183),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_119),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_115),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_72),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_106),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_43),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_104),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_91),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_189),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_187),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_0),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_225),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_0),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_1),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_186),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_225),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_189),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g276 ( 
.A(n_197),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_203),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_204),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_213),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_214),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_221),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_203),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_196),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_228),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_230),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_234),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_198),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_211),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_212),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_212),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_201),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_210),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_236),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_226),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_258),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_238),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_263),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_309),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_190),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_R g320 ( 
.A(n_262),
.B(n_226),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

AND3x1_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_246),
.C(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_309),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_261),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_271),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_246),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_269),
.B(n_233),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_188),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

BUFx8_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_279),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_260),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_281),
.B(n_191),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_194),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_275),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_292),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_292),
.B(n_206),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_306),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_277),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_319),
.B(n_207),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_233),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_240),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_240),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_338),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_311),
.B(n_364),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_34),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_35),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_208),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_209),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_314),
.B(n_297),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_215),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_319),
.B(n_217),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_330),
.A2(n_244),
.B1(n_219),
.B2(n_224),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

AO21x2_ASAP7_75t_L g409 ( 
.A1(n_313),
.A2(n_227),
.B(n_218),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_248),
.B1(n_232),
.B2(n_235),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_229),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_354),
.A2(n_237),
.B1(n_239),
.B2(n_241),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_247),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_249),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_252),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_36),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_336),
.B(n_253),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_336),
.B(n_254),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_316),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_37),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_334),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_362),
.B(n_296),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_321),
.B(n_41),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_348),
.B(n_352),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_312),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_321),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_383),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_430),
.A2(n_352),
.B1(n_358),
.B2(n_332),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_352),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_358),
.B1(n_361),
.B2(n_363),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_433),
.B(n_322),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_358),
.B1(n_361),
.B2(n_363),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_383),
.A2(n_342),
.B1(n_365),
.B2(n_347),
.Y(n_447)
);

O2A1O1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_369),
.A2(n_438),
.B(n_403),
.C(n_398),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_391),
.B(n_361),
.Y(n_450)
);

AND2x6_ASAP7_75t_SL g451 ( 
.A(n_400),
.B(n_366),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_327),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_432),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_363),
.B1(n_324),
.B2(n_335),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

AND2x6_ASAP7_75t_SL g458 ( 
.A(n_414),
.B(n_366),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_398),
.B(n_312),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_376),
.B(n_351),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_325),
.B1(n_327),
.B2(n_350),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_412),
.A2(n_325),
.B(n_342),
.Y(n_463)
);

AO22x1_ASAP7_75t_L g464 ( 
.A1(n_371),
.A2(n_365),
.B1(n_350),
.B2(n_347),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_343),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_343),
.B1(n_341),
.B2(n_283),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_375),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_415),
.B(n_315),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_374),
.B(n_397),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_341),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_367),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_379),
.B(n_341),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_415),
.B(n_317),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_360),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_369),
.B(n_290),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_381),
.B(n_295),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_SL g481 ( 
.A(n_433),
.B(n_317),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_397),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_395),
.B(n_323),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_409),
.A2(n_323),
.B1(n_92),
.B2(n_93),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_409),
.A2(n_373),
.B1(n_371),
.B2(n_434),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_412),
.B(n_42),
.Y(n_486)
);

INVx8_ASAP7_75t_L g487 ( 
.A(n_371),
.Y(n_487)
);

OR2x6_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_3),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_395),
.B(n_3),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_401),
.B(n_5),
.C(n_6),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_368),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_411),
.B(n_416),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_371),
.A2(n_94),
.B1(n_182),
.B2(n_181),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_5),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_420),
.B(n_45),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_420),
.B(n_46),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g498 ( 
.A(n_413),
.B(n_7),
.C(n_8),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_367),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_427),
.B(n_48),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_425),
.B(n_429),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_425),
.A2(n_97),
.B(n_179),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_429),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_399),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_429),
.B(n_7),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_424),
.B(n_49),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_424),
.B(n_8),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_424),
.B(n_50),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

NOR2x2_ASAP7_75t_L g512 ( 
.A(n_371),
.B(n_9),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_436),
.B(n_51),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_384),
.B(n_55),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_385),
.B(n_56),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_427),
.B(n_9),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_373),
.B(n_10),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_373),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_373),
.B(n_10),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_394),
.B(n_58),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_386),
.A2(n_105),
.B(n_177),
.Y(n_523)
);

INVx8_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_451),
.Y(n_526)
);

INVx3_ASAP7_75t_SL g527 ( 
.A(n_460),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_468),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_394),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_493),
.A2(n_373),
.B1(n_435),
.B2(n_418),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_452),
.B(n_387),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_472),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_394),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_492),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_394),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_502),
.B(n_418),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_476),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_505),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_483),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_482),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_478),
.A2(n_436),
.B1(n_418),
.B2(n_392),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_SL g552 ( 
.A(n_447),
.B(n_388),
.C(n_389),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_SL g553 ( 
.A(n_442),
.B(n_390),
.C(n_393),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_465),
.B(n_427),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_478),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_480),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_SL g559 ( 
.A(n_447),
.B(n_11),
.C(n_12),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_459),
.B(n_418),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_443),
.B(n_367),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_500),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_478),
.B(n_418),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_489),
.Y(n_564)
);

OR2x4_ASAP7_75t_L g565 ( 
.A(n_475),
.B(n_367),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_445),
.B(n_380),
.Y(n_569)
);

NOR3xp33_ASAP7_75t_SL g570 ( 
.A(n_490),
.B(n_11),
.C(n_12),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_495),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_444),
.A2(n_406),
.B1(n_421),
.B2(n_380),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

NOR3xp33_ASAP7_75t_SL g574 ( 
.A(n_477),
.B(n_14),
.C(n_15),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_518),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_445),
.B(n_380),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_442),
.B(n_380),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_473),
.B(n_392),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_458),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_499),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_499),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_464),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_536),
.B(n_448),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_572),
.A2(n_516),
.B(n_515),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_536),
.B(n_463),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_496),
.B(n_486),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_543),
.A2(n_444),
.B(n_446),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_534),
.B(n_463),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_561),
.A2(n_497),
.B(n_507),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_549),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_533),
.B(n_446),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_543),
.A2(n_487),
.B(n_509),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_538),
.A2(n_503),
.B(n_504),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_546),
.B(n_455),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_572),
.A2(n_501),
.B(n_523),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_560),
.B(n_461),
.Y(n_599)
);

AO31x2_ASAP7_75t_L g600 ( 
.A1(n_571),
.A2(n_521),
.A3(n_519),
.B(n_523),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_471),
.Y(n_601)
);

NOR2xp67_ASAP7_75t_L g602 ( 
.A(n_557),
.B(n_484),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_538),
.A2(n_501),
.B(n_485),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_461),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_577),
.A2(n_422),
.B(n_417),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_564),
.B(n_525),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_529),
.B(n_530),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_537),
.B(n_481),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_532),
.B(n_520),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_535),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_571),
.A2(n_514),
.B(n_494),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_560),
.A2(n_382),
.B(n_514),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_540),
.B(n_466),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_545),
.B(n_466),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_527),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_574),
.B(n_498),
.C(n_506),
.Y(n_619)
);

OAI21x1_ASAP7_75t_SL g620 ( 
.A1(n_575),
.A2(n_512),
.B(n_392),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_553),
.A2(n_508),
.B(n_517),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_545),
.B(n_382),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_542),
.A2(n_382),
.B(n_402),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_548),
.B(n_488),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_547),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_553),
.A2(n_408),
.B(n_422),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_542),
.A2(n_555),
.B(n_578),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_550),
.B(n_392),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_547),
.A2(n_382),
.B(n_402),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_583),
.A2(n_408),
.B(n_405),
.Y(n_631)
);

AO22x2_ASAP7_75t_L g632 ( 
.A1(n_569),
.A2(n_488),
.B1(n_392),
.B2(n_18),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_576),
.A2(n_417),
.B(n_419),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_554),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_583),
.A2(n_419),
.B(n_402),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_528),
.B(n_14),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_531),
.A2(n_419),
.B1(n_402),
.B2(n_423),
.Y(n_637)
);

AOI21xp33_ASAP7_75t_L g638 ( 
.A1(n_562),
.A2(n_16),
.B(n_18),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_605),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_633),
.A2(n_627),
.B(n_598),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_627),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_613),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_612),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_614),
.A2(n_552),
.B(n_570),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_613),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_624),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_634),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_607),
.Y(n_648)
);

AO21x2_ASAP7_75t_L g649 ( 
.A1(n_596),
.A2(n_552),
.B(n_584),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_601),
.B(n_528),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_624),
.Y(n_651)
);

AO21x2_ASAP7_75t_L g652 ( 
.A1(n_594),
.A2(n_582),
.B(n_580),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_586),
.B(n_556),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_594),
.B(n_547),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_626),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_633),
.A2(n_573),
.B(n_566),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_604),
.B(n_559),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_619),
.A2(n_531),
.B1(n_559),
.B2(n_585),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_589),
.A2(n_570),
.B(n_574),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_632),
.A2(n_558),
.B1(n_563),
.B2(n_531),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_606),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_591),
.A2(n_602),
.B1(n_597),
.B2(n_616),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_588),
.B(n_544),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_610),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_608),
.A2(n_568),
.B1(n_581),
.B2(n_563),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_599),
.B(n_531),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_635),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_611),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_590),
.A2(n_580),
.B(n_531),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_599),
.A2(n_563),
.B(n_558),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_593),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_595),
.A2(n_631),
.B(n_603),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_629),
.Y(n_673)
);

AO32x2_ASAP7_75t_L g674 ( 
.A1(n_600),
.A2(n_551),
.A3(n_565),
.B1(n_568),
.B2(n_524),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_632),
.A2(n_565),
.B1(n_524),
.B2(n_535),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_632),
.B(n_617),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_636),
.A2(n_526),
.B1(n_535),
.B2(n_524),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_419),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_615),
.A2(n_423),
.B(n_109),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_622),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_603),
.A2(n_423),
.B(n_108),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_621),
.B(n_59),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_592),
.A2(n_423),
.B(n_110),
.Y(n_684)
);

AO21x2_ASAP7_75t_L g685 ( 
.A1(n_589),
.A2(n_107),
.B(n_176),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_600),
.B(n_61),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_655),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_642),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_681),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_642),
.B(n_626),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_683),
.A2(n_620),
.B1(n_618),
.B2(n_609),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_648),
.A2(n_637),
.B1(n_617),
.B2(n_638),
.Y(n_692)
);

BUFx12f_ASAP7_75t_L g693 ( 
.A(n_642),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_657),
.A2(n_628),
.B1(n_622),
.B2(n_593),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_640),
.A2(n_587),
.B(n_623),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_658),
.A2(n_626),
.B1(n_600),
.B2(n_630),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_640),
.A2(n_600),
.B(n_626),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_671),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_645),
.B(n_62),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_658),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_645),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_645),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_646),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_653),
.Y(n_704)
);

OAI21xp33_ASAP7_75t_L g705 ( 
.A1(n_653),
.A2(n_19),
.B(n_20),
.Y(n_705)
);

NAND2x1p5_ASAP7_75t_L g706 ( 
.A(n_661),
.B(n_63),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_661),
.B(n_22),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_643),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_643),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_647),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_647),
.Y(n_711)
);

BUFx12f_ASAP7_75t_L g712 ( 
.A(n_655),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

INVx5_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_657),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_648),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_717)
);

CKINVDCx8_ASAP7_75t_R g718 ( 
.A(n_659),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_676),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_670),
.B(n_64),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_665),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_668),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_663),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_676),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_644),
.A2(n_32),
.B1(n_33),
.B2(n_65),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_670),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_676),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_644),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_664),
.B(n_76),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_662),
.B(n_77),
.Y(n_732)
);

AOI221xp5_ASAP7_75t_L g733 ( 
.A1(n_683),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_660),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_679),
.A2(n_90),
.B(n_96),
.C(n_98),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_682),
.A2(n_100),
.B(n_102),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_676),
.A2(n_103),
.B1(n_111),
.B2(n_113),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_663),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_659),
.B(n_114),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_675),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_675),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_644),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_SL g743 ( 
.A1(n_700),
.A2(n_644),
.B1(n_676),
.B2(n_679),
.Y(n_743)
);

OAI21xp33_ASAP7_75t_L g744 ( 
.A1(n_705),
.A2(n_686),
.B(n_677),
.Y(n_744)
);

AOI221xp5_ASAP7_75t_L g745 ( 
.A1(n_716),
.A2(n_686),
.B1(n_673),
.B2(n_666),
.C(n_669),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_709),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_704),
.B(n_659),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_720),
.A2(n_649),
.B1(n_673),
.B2(n_652),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_712),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_727),
.A2(n_669),
.B1(n_654),
.B2(n_649),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_710),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_726),
.A2(n_649),
.B1(n_652),
.B2(n_680),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_SL g753 ( 
.A1(n_722),
.A2(n_737),
.B1(n_729),
.B2(n_721),
.C(n_733),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_731),
.B(n_654),
.Y(n_754)
);

OAI21xp33_ASAP7_75t_L g755 ( 
.A1(n_694),
.A2(n_680),
.B(n_654),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_711),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_728),
.B(n_652),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_727),
.A2(n_721),
.B1(n_742),
.B2(n_730),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_717),
.A2(n_685),
.B1(n_641),
.B2(n_639),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_717),
.A2(n_685),
.B1(n_641),
.B2(n_639),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_725),
.B(n_674),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_708),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_714),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_721),
.A2(n_685),
.B1(n_682),
.B2(n_684),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_730),
.A2(n_641),
.B1(n_639),
.B2(n_678),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_735),
.A2(n_684),
.B(n_674),
.C(n_656),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_687),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_698),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_742),
.A2(n_674),
.B1(n_672),
.B2(n_667),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_713),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_740),
.A2(n_672),
.B(n_656),
.C(n_667),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_741),
.A2(n_667),
.B1(n_674),
.B2(n_137),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_695),
.A2(n_674),
.B(n_136),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_691),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_699),
.A2(n_734),
.B1(n_702),
.B2(n_692),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_738),
.B(n_140),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_701),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_692),
.A2(n_185),
.B1(n_148),
.B2(n_153),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_724),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_687),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_732),
.A2(n_707),
.B(n_706),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_689),
.A2(n_147),
.B1(n_154),
.B2(n_157),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_693),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_715),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_719),
.Y(n_785)
);

CKINVDCx6p67_ASAP7_75t_R g786 ( 
.A(n_715),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_697),
.A2(n_159),
.B(n_160),
.Y(n_787)
);

BUFx12f_ASAP7_75t_SL g788 ( 
.A(n_699),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_688),
.A2(n_718),
.B1(n_723),
.B2(n_696),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_761),
.B(n_739),
.Y(n_790)
);

AO21x2_ASAP7_75t_L g791 ( 
.A1(n_766),
.A2(n_736),
.B(n_703),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_746),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_751),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_747),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_756),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_757),
.B(n_779),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_757),
.B(n_706),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_772),
.A2(n_690),
.B(n_714),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_770),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_785),
.B(n_714),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_762),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_773),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_750),
.B(n_714),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_789),
.B(n_760),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_787),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_759),
.B(n_690),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_769),
.B(n_161),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_SL g808 ( 
.A1(n_758),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_759),
.A2(n_167),
.B(n_169),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_767),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_767),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_780),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_763),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_780),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_754),
.B(n_170),
.Y(n_816)
);

AO21x1_ASAP7_75t_L g817 ( 
.A1(n_772),
.A2(n_171),
.B(n_172),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_771),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_760),
.B(n_174),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_763),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_743),
.B(n_764),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_755),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_794),
.B(n_754),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_794),
.B(n_765),
.Y(n_824)
);

INVx8_ASAP7_75t_L g825 ( 
.A(n_813),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_792),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_821),
.A2(n_744),
.B1(n_778),
.B2(n_753),
.C(n_781),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_822),
.B(n_778),
.C(n_782),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_808),
.A2(n_775),
.B1(n_782),
.B2(n_745),
.Y(n_829)
);

OAI33xp33_ASAP7_75t_L g830 ( 
.A1(n_815),
.A2(n_776),
.A3(n_777),
.B1(n_786),
.B2(n_784),
.B3(n_752),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_808),
.A2(n_774),
.B1(n_788),
.B2(n_752),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_822),
.B(n_748),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_796),
.B(n_748),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_811),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_817),
.A2(n_783),
.B1(n_765),
.B2(n_749),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_811),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_792),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_820),
.B(n_749),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_793),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_790),
.B(n_763),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_820),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_793),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_795),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_796),
.B(n_763),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_801),
.B(n_768),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_841),
.B(n_820),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_841),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_836),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_823),
.B(n_821),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_837),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_837),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_840),
.B(n_812),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_833),
.B(n_815),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_842),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_842),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_833),
.B(n_790),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_843),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_843),
.Y(n_858)
);

NOR4xp25_ASAP7_75t_SL g859 ( 
.A(n_834),
.B(n_818),
.C(n_814),
.D(n_812),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_840),
.B(n_810),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_849),
.B(n_823),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_849),
.B(n_834),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_853),
.B(n_838),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_856),
.B(n_838),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_856),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_852),
.B(n_838),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_853),
.B(n_844),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_852),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_848),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_850),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_850),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_869),
.B(n_827),
.C(n_835),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_862),
.B(n_809),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_866),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_866),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_867),
.B(n_816),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_862),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_SL g879 ( 
.A1(n_868),
.A2(n_845),
.B(n_847),
.C(n_828),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_864),
.B(n_865),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_871),
.B(n_854),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_864),
.B(n_860),
.Y(n_882)
);

OAI32xp33_ASAP7_75t_L g883 ( 
.A1(n_873),
.A2(n_821),
.A3(n_863),
.B1(n_804),
.B2(n_861),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_872),
.A2(n_873),
.B(n_875),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_878),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_881),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_882),
.B(n_852),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_885),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_884),
.B(n_877),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_886),
.A2(n_879),
.B1(n_877),
.B2(n_817),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_888),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_889),
.Y(n_892)
);

NAND4xp25_ASAP7_75t_L g893 ( 
.A(n_890),
.B(n_883),
.C(n_829),
.D(n_831),
.Y(n_893)
);

XOR2xp5_ASAP7_75t_L g894 ( 
.A(n_889),
.B(n_832),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_892),
.B(n_880),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_SL g896 ( 
.A1(n_891),
.A2(n_893),
.B(n_881),
.C(n_894),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_892),
.B(n_807),
.C(n_819),
.Y(n_897)
);

NAND4xp25_ASAP7_75t_L g898 ( 
.A(n_892),
.B(n_874),
.C(n_816),
.D(n_887),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_SL g899 ( 
.A(n_892),
.B(n_876),
.C(n_859),
.Y(n_899)
);

A2O1A1O1Ixp25_ASAP7_75t_L g900 ( 
.A1(n_892),
.A2(n_818),
.B(n_854),
.C(n_855),
.D(n_798),
.Y(n_900)
);

NAND4xp25_ASAP7_75t_L g901 ( 
.A(n_892),
.B(n_887),
.C(n_807),
.D(n_798),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_892),
.B(n_807),
.C(n_819),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_900),
.A2(n_819),
.B(n_809),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_895),
.B(n_175),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_896),
.B(n_809),
.C(n_804),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_899),
.A2(n_867),
.B(n_847),
.Y(n_906)
);

AND4x1_ASAP7_75t_L g907 ( 
.A(n_897),
.B(n_830),
.C(n_803),
.D(n_797),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_902),
.A2(n_809),
.B1(n_803),
.B2(n_797),
.Y(n_908)
);

OAI221xp5_ASAP7_75t_SL g909 ( 
.A1(n_901),
.A2(n_847),
.B1(n_806),
.B2(n_824),
.C(n_813),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_905),
.A2(n_898),
.B1(n_809),
.B2(n_847),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_R g911 ( 
.A(n_904),
.B(n_813),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_906),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_903),
.B(n_855),
.Y(n_913)
);

NOR2x1_ASAP7_75t_SL g914 ( 
.A(n_909),
.B(n_858),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_907),
.Y(n_915)
);

AOI221xp5_ASAP7_75t_L g916 ( 
.A1(n_908),
.A2(n_824),
.B1(n_860),
.B2(n_852),
.C(n_802),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_R g917 ( 
.A(n_904),
.B(n_813),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_912),
.B(n_860),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_911),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_914),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_913),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_915),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_910),
.B(n_860),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_917),
.B(n_858),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_916),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_912),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_911),
.B(n_846),
.Y(n_927)
);

AND4x1_ASAP7_75t_L g928 ( 
.A(n_922),
.B(n_814),
.C(n_810),
.D(n_800),
.Y(n_928)
);

NAND4xp25_ASAP7_75t_L g929 ( 
.A(n_925),
.B(n_926),
.C(n_920),
.D(n_921),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_919),
.B(n_846),
.Y(n_930)
);

OA22x2_ASAP7_75t_L g931 ( 
.A1(n_918),
.A2(n_846),
.B1(n_851),
.B2(n_857),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_924),
.B(n_805),
.C(n_839),
.Y(n_932)
);

NOR2x1p5_ASAP7_75t_L g933 ( 
.A(n_918),
.B(n_846),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_923),
.A2(n_825),
.B1(n_805),
.B2(n_802),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_927),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_923),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_935),
.B(n_857),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_936),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_933),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_929),
.Y(n_940)
);

XNOR2x1_ASAP7_75t_L g941 ( 
.A(n_931),
.B(n_806),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_930),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_938),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_942),
.A2(n_934),
.B1(n_932),
.B2(n_928),
.Y(n_944)
);

OR4x1_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_826),
.C(n_795),
.D(n_825),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_943),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_944),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_946),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_947),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_948),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_949),
.A2(n_939),
.B(n_937),
.Y(n_951)
);

OAI22xp33_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_945),
.B1(n_941),
.B2(n_851),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_SL g953 ( 
.A1(n_952),
.A2(n_951),
.B1(n_825),
.B2(n_805),
.Y(n_953)
);

OAI221xp5_ASAP7_75t_R g954 ( 
.A1(n_953),
.A2(n_825),
.B1(n_805),
.B2(n_800),
.C(n_791),
.Y(n_954)
);

AOI211xp5_ASAP7_75t_L g955 ( 
.A1(n_954),
.A2(n_801),
.B(n_799),
.C(n_790),
.Y(n_955)
);


endmodule