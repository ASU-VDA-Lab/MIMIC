module fake_netlist_5_1349_n_1516 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_389, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_397, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_400, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_395, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_402, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_66, n_177, n_60, n_403, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_391, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1516);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_389;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_397;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_400;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_395;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_402;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_403;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_391;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1516;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_418;
wire n_968;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_268),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_175),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_208),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_106),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_253),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_200),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_375),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_146),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_250),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_178),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_222),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_365),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_298),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_59),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_374),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_75),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_71),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_380),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_95),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_53),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_258),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_50),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_171),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_143),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_332),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_65),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_266),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_129),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_131),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_201),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_181),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_19),
.B(n_71),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_362),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_261),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_229),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_230),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_38),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_260),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_237),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_254),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_59),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_104),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_337),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_182),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_321),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_401),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_397),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_255),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_264),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_303),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_346),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_101),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_345),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_339),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_180),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_389),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_141),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_85),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_47),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_241),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_154),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_77),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_225),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_350),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_99),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_79),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_103),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_69),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_347),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_377),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_274),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_314),
.B(n_236),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_66),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_5),
.Y(n_483)
);

BUFx2_ASAP7_75t_SL g484 ( 
.A(n_376),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_348),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_244),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_147),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_73),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_184),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_372),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_312),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_76),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_162),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_68),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_12),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_395),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_104),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_115),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_243),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_198),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_16),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_209),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_309),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_68),
.B(n_125),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_126),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_80),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_40),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_83),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_238),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_176),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_356),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_58),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_152),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_308),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_277),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_70),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_7),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_116),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_95),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_381),
.B(n_134),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_276),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_67),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_203),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_8),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_63),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_108),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_353),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_100),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_249),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_292),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_213),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_355),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_257),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_132),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_91),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_159),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_359),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_204),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_311),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_306),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_270),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_338),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_100),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_382),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_174),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_307),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_343),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_49),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_402),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_28),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_283),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_73),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_114),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_262),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_177),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_25),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_173),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_317),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_214),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_235),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_265),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_119),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_188),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_89),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_16),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_148),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_13),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_37),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_195),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_294),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_98),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_289),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_305),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_263),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_330),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_313),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_109),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_151),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_90),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_150),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_18),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_56),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_392),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_340),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_288),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_135),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_144),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_107),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_366),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_44),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_272),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_301),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_24),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_296),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_115),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_393),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_316),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_149),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_433),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_461),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_433),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_433),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_489),
.A2(n_136),
.B(n_133),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_448),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_476),
.B(n_0),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_523),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_448),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_467),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_446),
.Y(n_616)
);

OA21x2_ASAP7_75t_L g617 ( 
.A1(n_421),
.A2(n_0),
.B(n_1),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_467),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_448),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_471),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_471),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_487),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_505),
.B(n_1),
.Y(n_623)
);

OAI22x1_ASAP7_75t_R g624 ( 
.A1(n_507),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_624)
);

CKINVDCx11_ASAP7_75t_R g625 ( 
.A(n_501),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_471),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_471),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_583),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_501),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_503),
.B(n_2),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_505),
.B(n_3),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_451),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_422),
.A2(n_4),
.B(n_5),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_583),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_583),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_519),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_408),
.B(n_6),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_503),
.B(n_570),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

BUFx12f_ASAP7_75t_L g643 ( 
.A(n_544),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_9),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_483),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_428),
.B(n_9),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_494),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_489),
.B(n_10),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_487),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_551),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_409),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_488),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_423),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_654)
);

NOR2x1_ASAP7_75t_L g655 ( 
.A(n_481),
.B(n_521),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_510),
.B(n_137),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_428),
.B(n_11),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_470),
.B(n_13),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_492),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_497),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_510),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_14),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_498),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_508),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_510),
.B(n_138),
.Y(n_665)
);

CKINVDCx6p67_ASAP7_75t_R g666 ( 
.A(n_544),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_443),
.A2(n_140),
.B(n_139),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_525),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_510),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_454),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_557),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_566),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_469),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_572),
.A2(n_582),
.B(n_578),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_594),
.Y(n_676)
);

XNOR2x2_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_15),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_454),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_587),
.B(n_18),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_490),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_405),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_575),
.Y(n_682)
);

OA21x2_ASAP7_75t_L g683 ( 
.A1(n_411),
.A2(n_20),
.B(n_21),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_575),
.Y(n_684)
);

BUFx8_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_670),
.B(n_533),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_631),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_601),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_646),
.A2(n_419),
.B1(n_425),
.B2(n_424),
.Y(n_689)
);

INVx8_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_618),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_635),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_601),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_641),
.B(n_552),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_603),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_607),
.Y(n_697)
);

INVxp67_ASAP7_75t_R g698 ( 
.A(n_624),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_635),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_636),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_603),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_678),
.B(n_552),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_655),
.B(n_514),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_604),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_604),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

BUFx6f_ASAP7_75t_SL g707 ( 
.A(n_630),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_675),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_605),
.Y(n_709)
);

AOI21x1_ASAP7_75t_L g710 ( 
.A1(n_681),
.A2(n_414),
.B(n_413),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_608),
.B(n_522),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_602),
.A2(n_679),
.B1(n_658),
.B2(n_652),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_657),
.B(n_662),
.Y(n_713)
);

CKINVDCx11_ASAP7_75t_R g714 ( 
.A(n_625),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_607),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_614),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_610),
.B(n_649),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_615),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_621),
.A2(n_434),
.B(n_429),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_621),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_607),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_626),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_647),
.B(n_542),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_627),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_627),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_628),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_652),
.B(n_408),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_645),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_647),
.B(n_576),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_602),
.B(n_531),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_609),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_675),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_609),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_727),
.B(n_648),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_689),
.B(n_674),
.C(n_654),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_714),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_733),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_713),
.B(n_717),
.C(n_708),
.Y(n_739)
);

OA21x2_ASAP7_75t_L g740 ( 
.A1(n_719),
.A2(n_606),
.B(n_667),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_733),
.A2(n_644),
.B1(n_630),
.B2(n_683),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_713),
.A2(n_644),
.B1(n_683),
.B2(n_617),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_691),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_697),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_692),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_700),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_731),
.B(n_613),
.Y(n_748)
);

BUFx5_ASAP7_75t_L g749 ( 
.A(n_716),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_706),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_717),
.A2(n_695),
.B1(n_683),
.B2(n_617),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_693),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_712),
.A2(n_418),
.B1(n_447),
.B2(n_439),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_702),
.B(n_629),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_697),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_711),
.A2(n_632),
.B(n_623),
.C(n_640),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_629),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_723),
.B(n_643),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_730),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_707),
.A2(n_462),
.B1(n_502),
.B2(n_485),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_707),
.B(n_680),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_732),
.B(n_684),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_693),
.B(n_643),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_714),
.B(n_632),
.C(n_623),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_707),
.B(n_600),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_732),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_699),
.B(n_666),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_687),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_699),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_729),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_734),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_734),
.B(n_684),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_710),
.B(n_406),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_729),
.B(n_611),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_709),
.B(n_612),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_718),
.B(n_611),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_710),
.B(n_407),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_688),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_720),
.B(n_625),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_697),
.B(n_640),
.Y(n_781)
);

BUFx5_ASAP7_75t_L g782 ( 
.A(n_716),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_698),
.A2(n_504),
.B1(n_438),
.B2(n_427),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_722),
.A2(n_410),
.B1(n_595),
.B2(n_588),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_688),
.B(n_612),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_694),
.B(n_685),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_696),
.B(n_638),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_696),
.B(n_645),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_728),
.B(n_616),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_728),
.B(n_616),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_715),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_715),
.B(n_412),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_701),
.B(n_685),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_715),
.B(n_415),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_722),
.B(n_656),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_457),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_704),
.B(n_656),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_705),
.B(n_416),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_698),
.A2(n_639),
.B1(n_431),
.B2(n_468),
.Y(n_799)
);

BUFx12f_ASAP7_75t_L g800 ( 
.A(n_737),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_735),
.B(n_633),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_745),
.B(n_651),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_788),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_753),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_759),
.B(n_651),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_789),
.B(n_653),
.Y(n_806)
);

CKINVDCx8_ASAP7_75t_R g807 ( 
.A(n_754),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_738),
.A2(n_690),
.B(n_687),
.Y(n_808)
);

A2O1A1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_739),
.A2(n_410),
.B(n_436),
.C(n_435),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_775),
.B(n_633),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_738),
.A2(n_690),
.B(n_687),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_739),
.A2(n_420),
.B1(n_430),
.B2(n_417),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_756),
.A2(n_673),
.B(n_660),
.C(n_663),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_741),
.A2(n_437),
.B1(n_442),
.B2(n_441),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_748),
.B(n_450),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_761),
.B(n_474),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_752),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_751),
.A2(n_719),
.B(n_634),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_742),
.A2(n_725),
.B(n_724),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_757),
.B(n_432),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_781),
.A2(n_726),
.B(n_725),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_784),
.A2(n_444),
.B1(n_449),
.B2(n_445),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_785),
.A2(n_776),
.B(n_798),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_761),
.B(n_440),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_744),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_797),
.A2(n_634),
.B(n_617),
.Y(n_826)
);

AOI21xp33_ASAP7_75t_L g827 ( 
.A1(n_783),
.A2(n_634),
.B(n_477),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_790),
.B(n_659),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_736),
.A2(n_453),
.B1(n_456),
.B2(n_452),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_770),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_777),
.B(n_672),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_771),
.B(n_459),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_766),
.B(n_475),
.Y(n_833)
);

INVx11_ASAP7_75t_L g834 ( 
.A(n_768),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_743),
.B(n_746),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_769),
.A2(n_622),
.B(n_619),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_760),
.B(n_482),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_747),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_780),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_792),
.A2(n_642),
.B(n_622),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_750),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_794),
.A2(n_650),
.B(n_642),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_787),
.B(n_676),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_786),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_758),
.B(n_495),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_763),
.A2(n_661),
.B(n_650),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_740),
.A2(n_665),
.B(n_656),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_767),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_793),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_765),
.B(n_656),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_773),
.A2(n_661),
.B(n_650),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_796),
.B(n_779),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_772),
.B(n_664),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_762),
.A2(n_458),
.B1(n_460),
.B2(n_455),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_749),
.B(n_472),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_749),
.B(n_473),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_795),
.B(n_463),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_744),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_749),
.B(n_491),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_749),
.B(n_493),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_791),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_749),
.B(n_782),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_799),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_782),
.B(n_496),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_782),
.B(n_499),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_764),
.B(n_464),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_755),
.B(n_664),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_782),
.B(n_509),
.Y(n_869)
);

OAI321xp33_ASAP7_75t_L g870 ( 
.A1(n_799),
.A2(n_513),
.A3(n_532),
.B1(n_540),
.B2(n_534),
.C(n_520),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_791),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_791),
.A2(n_561),
.B1(n_564),
.B2(n_548),
.Y(n_872)
);

OA22x2_ASAP7_75t_L g873 ( 
.A1(n_799),
.A2(n_677),
.B1(n_506),
.B2(n_516),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_752),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_738),
.B(n_567),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_738),
.A2(n_571),
.B(n_577),
.C(n_574),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_738),
.B(n_579),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_788),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_788),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_788),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_789),
.B(n_668),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_775),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_759),
.B(n_465),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_738),
.B(n_581),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_735),
.B(n_517),
.C(n_512),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_738),
.B(n_586),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_789),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_738),
.B(n_590),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_735),
.B(n_527),
.C(n_526),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_738),
.B(n_597),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_738),
.B(n_665),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_738),
.A2(n_665),
.B(n_478),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_748),
.B(n_536),
.C(n_529),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_735),
.B(n_668),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_789),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_738),
.A2(n_665),
.B(n_479),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_745),
.B(n_484),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_759),
.B(n_466),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_739),
.A2(n_486),
.B1(n_500),
.B2(n_480),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_744),
.Y(n_900)
);

OAI21x1_ASAP7_75t_SL g901 ( 
.A1(n_813),
.A2(n_671),
.B(n_142),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_894),
.B(n_511),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_818),
.A2(n_682),
.B(n_669),
.Y(n_903)
);

AND2x6_ASAP7_75t_L g904 ( 
.A(n_891),
.B(n_575),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_819),
.A2(n_524),
.B(n_515),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_815),
.A2(n_530),
.B1(n_535),
.B2(n_528),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_882),
.Y(n_907)
);

OAI21x1_ASAP7_75t_SL g908 ( 
.A1(n_875),
.A2(n_671),
.B(n_145),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_826),
.A2(n_538),
.B(n_537),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_807),
.B(n_549),
.Y(n_910)
);

AO31x2_ASAP7_75t_L g911 ( 
.A1(n_809),
.A2(n_599),
.A3(n_24),
.B(n_22),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_816),
.A2(n_541),
.B(n_543),
.C(n_539),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_801),
.B(n_553),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_853),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_814),
.A2(n_546),
.B1(n_547),
.B2(n_545),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_847),
.A2(n_555),
.B(n_550),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_839),
.B(n_554),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_829),
.A2(n_558),
.B(n_559),
.C(n_556),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_863),
.A2(n_682),
.B(n_669),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_878),
.B(n_562),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_877),
.A2(n_584),
.B(n_573),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_810),
.B(n_565),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_887),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_880),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_805),
.B(n_569),
.C(n_568),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_823),
.A2(n_896),
.B(n_892),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_802),
.B(n_589),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_803),
.B(n_585),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_858),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_821),
.A2(n_155),
.B(n_153),
.Y(n_930)
);

INVx6_ASAP7_75t_SL g931 ( 
.A(n_897),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_879),
.B(n_592),
.Y(n_932)
);

AOI21xp33_ASAP7_75t_L g933 ( 
.A1(n_837),
.A2(n_591),
.B(n_593),
.Y(n_933)
);

OA22x2_ASAP7_75t_L g934 ( 
.A1(n_804),
.A2(n_598),
.B1(n_25),
.B2(n_22),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_SL g935 ( 
.A1(n_825),
.A2(n_599),
.B(n_157),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_884),
.A2(n_158),
.B(n_156),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_886),
.A2(n_161),
.B(n_160),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_888),
.A2(n_164),
.B(n_163),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_817),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_808),
.A2(n_404),
.B(n_166),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_811),
.A2(n_403),
.B(n_167),
.Y(n_941)
);

NOR4xp25_ASAP7_75t_L g942 ( 
.A(n_870),
.B(n_27),
.C(n_23),
.D(n_26),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_890),
.A2(n_168),
.B(n_165),
.Y(n_943)
);

AO32x2_ASAP7_75t_L g944 ( 
.A1(n_822),
.A2(n_28),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_835),
.A2(n_170),
.B(n_169),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_L g946 ( 
.A(n_833),
.B(n_29),
.C(n_30),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_881),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_895),
.B(n_30),
.Y(n_948)
);

BUFx4_ASAP7_75t_SL g949 ( 
.A(n_897),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_844),
.B(n_172),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_830),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_874),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_881),
.B(n_31),
.Y(n_953)
);

AO31x2_ASAP7_75t_L g954 ( 
.A1(n_855),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_800),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_806),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_856),
.A2(n_861),
.B(n_860),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_834),
.B(n_33),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_865),
.A2(n_183),
.B(n_179),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_864),
.A2(n_186),
.B1(n_187),
.B2(n_185),
.Y(n_960)
);

OA22x2_ASAP7_75t_L g961 ( 
.A1(n_824),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_831),
.B(n_189),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_838),
.B(n_841),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_885),
.B(n_34),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_889),
.B(n_35),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_806),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_828),
.B(n_36),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_858),
.Y(n_968)
);

BUFx4f_ASAP7_75t_SL g969 ( 
.A(n_883),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_876),
.A2(n_191),
.B(n_190),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_850),
.A2(n_193),
.B1(n_194),
.B2(n_192),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_866),
.A2(n_197),
.B(n_196),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_828),
.B(n_37),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_827),
.A2(n_845),
.B(n_893),
.C(n_812),
.Y(n_974)
);

AO31x2_ASAP7_75t_L g975 ( 
.A1(n_869),
.A2(n_40),
.A3(n_38),
.B(n_39),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_849),
.B(n_199),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_848),
.Y(n_977)
);

AO22x2_ASAP7_75t_L g978 ( 
.A1(n_873),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_836),
.A2(n_205),
.B(n_202),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_899),
.A2(n_207),
.B1(n_210),
.B2(n_206),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_820),
.B(n_41),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_843),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_857),
.A2(n_212),
.B(n_211),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_832),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_898),
.B(n_867),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_859),
.B(n_215),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_859),
.A2(n_217),
.B(n_216),
.Y(n_987)
);

AND2x6_ASAP7_75t_L g988 ( 
.A(n_900),
.B(n_218),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_862),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_862),
.B(n_871),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_862),
.B(n_42),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_854),
.B(n_43),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_871),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_871),
.B(n_43),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_900),
.A2(n_220),
.B1(n_221),
.B2(n_219),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_872),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_900),
.B(n_44),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_840),
.B(n_45),
.Y(n_998)
);

OA22x2_ASAP7_75t_L g999 ( 
.A1(n_842),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_846),
.A2(n_399),
.B(n_224),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_851),
.B(n_223),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_858),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_818),
.A2(n_227),
.B(n_226),
.Y(n_1003)
);

AOI221x1_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_271),
.B1(n_398),
.B2(n_396),
.C(n_394),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_894),
.B(n_48),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_810),
.Y(n_1006)
);

AOI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_815),
.A2(n_48),
.B(n_49),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_809),
.A2(n_52),
.A3(n_50),
.B(n_51),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_882),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_SL g1010 ( 
.A1(n_813),
.A2(n_231),
.B(n_228),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_894),
.B(n_51),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_52),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_818),
.A2(n_233),
.B(n_232),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_815),
.A2(n_53),
.B(n_54),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_839),
.B(n_234),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_868),
.Y(n_1016)
);

AO22x2_ASAP7_75t_L g1017 ( 
.A1(n_829),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_R g1018 ( 
.A(n_800),
.B(n_55),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_815),
.A2(n_60),
.B(n_57),
.C(n_58),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_894),
.B(n_57),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_810),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_894),
.B(n_60),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_894),
.B(n_61),
.Y(n_1023)
);

INVx3_ASAP7_75t_SL g1024 ( 
.A(n_897),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_894),
.B(n_61),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_815),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_801),
.B(n_62),
.Y(n_1027)
);

OA22x2_ASAP7_75t_L g1028 ( 
.A1(n_804),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_1028)
);

AOI211x1_ASAP7_75t_L g1029 ( 
.A1(n_829),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_881),
.B(n_239),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_878),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_815),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_801),
.B(n_72),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_810),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_882),
.B(n_240),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_887),
.B(n_242),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_894),
.B(n_74),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_810),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_801),
.B(n_76),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_818),
.A2(n_246),
.B(n_245),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_810),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_894),
.B(n_77),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_818),
.A2(n_248),
.B(n_247),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_818),
.A2(n_252),
.B(n_251),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_810),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_801),
.B(n_78),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_SL g1047 ( 
.A1(n_813),
.A2(n_259),
.B(n_256),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_801),
.B(n_80),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_974),
.A2(n_299),
.B(n_390),
.C(n_388),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_984),
.B(n_81),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_926),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_1052)
);

INVx6_ASAP7_75t_L g1053 ( 
.A(n_955),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1006),
.B(n_82),
.Y(n_1054)
);

AO32x2_ASAP7_75t_L g1055 ( 
.A1(n_942),
.A2(n_84),
.A3(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_923),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_939),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_957),
.A2(n_84),
.A3(n_86),
.B(n_87),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_951),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_269),
.B(n_267),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_949),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_907),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1034),
.A2(n_310),
.B1(n_387),
.B2(n_385),
.Y(n_1063)
);

AND2x4_ASAP7_75t_SL g1064 ( 
.A(n_929),
.B(n_968),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_931),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_989),
.B(n_273),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1041),
.B(n_88),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1045),
.B(n_88),
.Y(n_1068)
);

INVx4_ASAP7_75t_SL g1069 ( 
.A(n_988),
.Y(n_1069)
);

OAI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_1021),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.C(n_92),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_1043),
.A2(n_318),
.B(n_384),
.C(n_383),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_992),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_927),
.A2(n_315),
.B1(n_379),
.B2(n_378),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_917),
.A2(n_93),
.B(n_94),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_964),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_931),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1038),
.B(n_96),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_SL g1078 ( 
.A1(n_969),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_929),
.Y(n_1079)
);

AOI222xp33_ASAP7_75t_L g1080 ( 
.A1(n_1027),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.C1(n_106),
.C2(n_107),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1016),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_970),
.A2(n_320),
.B(n_373),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_910),
.B(n_102),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_965),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_913),
.B(n_110),
.Y(n_1085)
);

AO21x2_ASAP7_75t_L g1086 ( 
.A1(n_909),
.A2(n_319),
.B(n_370),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1014),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_994),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_981),
.A2(n_933),
.B1(n_1007),
.B2(n_1030),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_1004),
.A2(n_111),
.A3(n_112),
.B(n_113),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_947),
.A2(n_322),
.B1(n_369),
.B2(n_368),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_1024),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_902),
.B(n_113),
.Y(n_1093)
);

OAI22x1_ASAP7_75t_L g1094 ( 
.A1(n_996),
.A2(n_958),
.B1(n_1046),
.B2(n_1039),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_930),
.A2(n_323),
.B(n_367),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1005),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_1009),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_948),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_940),
.A2(n_304),
.B(n_364),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_967),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1033),
.B(n_120),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1040),
.A2(n_302),
.B(n_363),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_963),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_941),
.A2(n_300),
.B(n_361),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_978),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.C(n_123),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_922),
.Y(n_1106)
);

INVx6_ASAP7_75t_L g1107 ( 
.A(n_1030),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_966),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1048),
.B(n_121),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_1010),
.A2(n_297),
.B(n_360),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_956),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1011),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1044),
.A2(n_324),
.B(n_358),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_919),
.A2(n_295),
.B(n_357),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_906),
.B(n_124),
.C(n_125),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_914),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_905),
.A2(n_293),
.B(n_351),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_929),
.Y(n_1118)
);

CKINVDCx11_ASAP7_75t_R g1119 ( 
.A(n_924),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_979),
.A2(n_291),
.B(n_349),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_L g1121 ( 
.A(n_988),
.B(n_290),
.Y(n_1121)
);

OAI211xp5_ASAP7_75t_L g1122 ( 
.A1(n_973),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1031),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1012),
.A2(n_127),
.B(n_128),
.C(n_129),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1019),
.A2(n_130),
.A3(n_275),
.B(n_278),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_977),
.Y(n_1126)
);

AOI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_928),
.A2(n_130),
.B(n_279),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1000),
.A2(n_280),
.B(n_281),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_982),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1026),
.A2(n_286),
.B(n_287),
.C(n_325),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_953),
.Y(n_1131)
);

BUFx10_ASAP7_75t_L g1132 ( 
.A(n_988),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_925),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_991),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_932),
.B(n_329),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_990),
.A2(n_916),
.B(n_962),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_968),
.Y(n_1137)
);

AO21x2_ASAP7_75t_L g1138 ( 
.A1(n_901),
.A2(n_331),
.B(n_334),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_SL g1139 ( 
.A1(n_908),
.A2(n_335),
.B(n_336),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1020),
.B(n_1022),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_993),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_946),
.A2(n_341),
.B1(n_342),
.B2(n_344),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_SL g1143 ( 
.A(n_1018),
.B(n_391),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_993),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1023),
.A2(n_1042),
.B1(n_1037),
.B2(n_1025),
.Y(n_1146)
);

NAND2x1p5_ASAP7_75t_L g1147 ( 
.A(n_989),
.B(n_993),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_976),
.A2(n_961),
.B1(n_978),
.B2(n_999),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1002),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1015),
.A2(n_920),
.B1(n_916),
.B2(n_1002),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_934),
.A2(n_1028),
.B1(n_985),
.B2(n_1017),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_911),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_998),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_936),
.A2(n_938),
.B(n_937),
.C(n_983),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1017),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_911),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_921),
.B(n_912),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_950),
.A2(n_1035),
.B1(n_980),
.B2(n_915),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_911),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_971),
.A2(n_1036),
.B1(n_1032),
.B2(n_1029),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_988),
.A2(n_960),
.B1(n_1013),
.B2(n_995),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1008),
.Y(n_1162)
);

AND2x4_ASAP7_75t_SL g1163 ( 
.A(n_1001),
.B(n_935),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_1001),
.B(n_944),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_904),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1008),
.B(n_944),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_959),
.A2(n_972),
.B(n_945),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_986),
.A2(n_1013),
.B1(n_943),
.B2(n_987),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_904),
.A2(n_918),
.B(n_1008),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_904),
.B(n_944),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_954),
.B(n_975),
.Y(n_1171)
);

AOI31xp67_ASAP7_75t_L g1172 ( 
.A1(n_954),
.A2(n_975),
.A3(n_778),
.B(n_774),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_975),
.A2(n_738),
.B(n_926),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_923),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_955),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_SL g1176 ( 
.A1(n_1010),
.A2(n_1047),
.B(n_908),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_974),
.A2(n_739),
.B1(n_926),
.B2(n_741),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_984),
.B(n_894),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_926),
.A2(n_957),
.B(n_1003),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_989),
.B(n_907),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_974),
.A2(n_815),
.B(n_816),
.C(n_926),
.Y(n_1181)
);

OAI222xp33_ASAP7_75t_L g1182 ( 
.A1(n_1028),
.A2(n_934),
.B1(n_961),
.B2(n_873),
.C1(n_807),
.C2(n_654),
.Y(n_1182)
);

NAND3x1_ASAP7_75t_L g1183 ( 
.A(n_958),
.B(n_753),
.C(n_736),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_926),
.A2(n_903),
.B(n_1003),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_926),
.A2(n_903),
.B(n_1003),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1088),
.B(n_1100),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1119),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1057),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1059),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1132),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1132),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1053),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1053),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1056),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1062),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1049),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1069),
.B(n_1126),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1106),
.B(n_1054),
.Y(n_1198)
);

BUFx2_ASAP7_75t_SL g1199 ( 
.A(n_1175),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1178),
.B(n_1103),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1067),
.B(n_1103),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1174),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1108),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1105),
.A2(n_1084),
.B1(n_1075),
.B2(n_1072),
.Y(n_1204)
);

CKINVDCx14_ASAP7_75t_R g1205 ( 
.A(n_1061),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1149),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1069),
.B(n_1123),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1083),
.A2(n_1183),
.B1(n_1089),
.B2(n_1080),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1140),
.B(n_1164),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1087),
.A2(n_1074),
.B1(n_1115),
.B2(n_1070),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1097),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1081),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1152),
.A2(n_1159),
.B(n_1171),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1177),
.A2(n_1150),
.B(n_1136),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1137),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1164),
.B(n_1181),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1134),
.B(n_1144),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1137),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1051),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1107),
.B(n_1180),
.Y(n_1221)
);

NAND2x1_ASAP7_75t_L g1222 ( 
.A(n_1141),
.B(n_1145),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1162),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1092),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1131),
.B(n_1153),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1152),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1151),
.B(n_1085),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1098),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1156),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1064),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1164),
.B(n_1146),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1065),
.B(n_1076),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1079),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1107),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1155),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1147),
.Y(n_1237)
);

CKINVDCx9p33_ASAP7_75t_R g1238 ( 
.A(n_1068),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1163),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1169),
.A2(n_1154),
.B(n_1102),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1109),
.B(n_1077),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1170),
.A2(n_1160),
.A3(n_1060),
.B(n_1052),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1117),
.A2(n_1157),
.B(n_1161),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1118),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1165),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1172),
.A2(n_1135),
.B(n_1158),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1125),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1148),
.A2(n_1164),
.B(n_1166),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1096),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1063),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1112),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1094),
.B(n_1179),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1078),
.A2(n_1142),
.B1(n_1082),
.B2(n_1124),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1143),
.B(n_1127),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1058),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_1130),
.B(n_1073),
.C(n_1133),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1184),
.B(n_1185),
.Y(n_1257)
);

AO21x1_ASAP7_75t_SL g1258 ( 
.A1(n_1182),
.A2(n_1129),
.B(n_1055),
.Y(n_1258)
);

AOI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1184),
.A2(n_1185),
.B(n_1176),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1055),
.B(n_1122),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1082),
.B(n_1168),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1058),
.Y(n_1262)
);

INVx8_ASAP7_75t_L g1263 ( 
.A(n_1066),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1058),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1091),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1165),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1090),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1090),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1139),
.Y(n_1269)
);

CKINVDCx14_ASAP7_75t_R g1270 ( 
.A(n_1110),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_L g1271 ( 
.A(n_1114),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1138),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1099),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1128),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1120),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1104),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1050),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1113),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1086),
.B(n_1114),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1095),
.Y(n_1280)
);

AOI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1167),
.A2(n_1173),
.B(n_1177),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1071),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1167),
.A2(n_1033),
.B1(n_1083),
.B2(n_1028),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1230),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1201),
.B(n_1227),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1243),
.A2(n_1248),
.B1(n_1253),
.B2(n_1254),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1198),
.B(n_1218),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1186),
.B(n_1225),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1225),
.B(n_1229),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1223),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1188),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1220),
.B(n_1209),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1189),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1209),
.B(n_1241),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1214),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1200),
.B(n_1194),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1226),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1197),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1203),
.B(n_1213),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1204),
.A2(n_1211),
.B1(n_1258),
.B2(n_1283),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1210),
.B(n_1248),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1194),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1206),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1202),
.B(n_1203),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1239),
.B(n_1234),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1206),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1239),
.B(n_1190),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1190),
.B(n_1191),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1219),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1243),
.A2(n_1253),
.B1(n_1232),
.B2(n_1250),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1206),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1266),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1191),
.B(n_1197),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1210),
.B(n_1283),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1208),
.B(n_1236),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1208),
.B(n_1196),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1207),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1204),
.A2(n_1211),
.B1(n_1251),
.B2(n_1249),
.Y(n_1318)
);

INVx3_ASAP7_75t_SL g1319 ( 
.A(n_1192),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1212),
.B(n_1199),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1212),
.B(n_1244),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1266),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1221),
.B(n_1216),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1265),
.A2(n_1260),
.B1(n_1232),
.B2(n_1217),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1221),
.B(n_1216),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1235),
.B(n_1221),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1235),
.B(n_1237),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1235),
.B(n_1252),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1252),
.B(n_1233),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1259),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1267),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1217),
.B(n_1233),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1247),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1268),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1193),
.B(n_1228),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1255),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1231),
.B(n_1263),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1245),
.B(n_1205),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1245),
.B(n_1205),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1262),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1222),
.B(n_1263),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1187),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1263),
.B(n_1195),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1238),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1269),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1242),
.B(n_1256),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1187),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1242),
.B(n_1256),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1270),
.B(n_1187),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1257),
.B(n_1238),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1257),
.B(n_1264),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1246),
.B(n_1240),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1246),
.B(n_1240),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1304),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1343),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1301),
.B(n_1281),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1337),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1296),
.Y(n_1359)
);

OR2x6_ASAP7_75t_SL g1360 ( 
.A(n_1351),
.B(n_1261),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1305),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1341),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1338),
.B(n_1344),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1301),
.B(n_1278),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1292),
.B(n_1271),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1343),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1288),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1290),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1289),
.B(n_1282),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1294),
.B(n_1277),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1286),
.B(n_1272),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1286),
.B(n_1272),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1287),
.B(n_1261),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1329),
.B(n_1328),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1324),
.B(n_1215),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1346),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1324),
.B(n_1285),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1352),
.B(n_1280),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1323),
.B(n_1273),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1346),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1331),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1299),
.B(n_1279),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1334),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1347),
.B(n_1271),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1297),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1276),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1302),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1295),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1309),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1309),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1318),
.B(n_1275),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_1348),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1364),
.B(n_1353),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1364),
.B(n_1357),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1379),
.Y(n_1397)
);

OAI21xp33_ASAP7_75t_L g1398 ( 
.A1(n_1377),
.A2(n_1300),
.B(n_1310),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1359),
.B(n_1314),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1357),
.B(n_1354),
.Y(n_1400)
);

AND2x4_ASAP7_75t_SL g1401 ( 
.A(n_1376),
.B(n_1325),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1355),
.B(n_1300),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1388),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1390),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1358),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1380),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1358),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1374),
.B(n_1295),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1362),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1362),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1382),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1367),
.B(n_1350),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1383),
.B(n_1391),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1385),
.B(n_1330),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1389),
.B(n_1332),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1385),
.B(n_1333),
.Y(n_1417)
);

NAND2x1_ASAP7_75t_SL g1418 ( 
.A(n_1375),
.B(n_1284),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1382),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1284),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1291),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1377),
.B(n_1321),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1371),
.B(n_1293),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1384),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1409),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1409),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1396),
.B(n_1360),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1418),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1405),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1396),
.B(n_1360),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1407),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1400),
.B(n_1386),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1411),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1419),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1425),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1410),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1421),
.B(n_1381),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1401),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1397),
.B(n_1406),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1421),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1418),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1395),
.B(n_1378),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1398),
.A2(n_1372),
.B1(n_1371),
.B2(n_1365),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1446),
.A2(n_1413),
.B(n_1345),
.C(n_1363),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1446),
.B(n_1403),
.C(n_1399),
.Y(n_1448)
);

NOR4xp25_ASAP7_75t_L g1449 ( 
.A(n_1428),
.B(n_1404),
.C(n_1369),
.D(n_1402),
.Y(n_1449)
);

AND2x2_ASAP7_75t_SL g1450 ( 
.A(n_1428),
.B(n_1393),
.Y(n_1450)
);

AOI32xp33_ASAP7_75t_L g1451 ( 
.A1(n_1431),
.A2(n_1372),
.A3(n_1424),
.B1(n_1375),
.B2(n_1422),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1429),
.A2(n_1444),
.B(n_1431),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1426),
.Y(n_1453)
);

AOI32xp33_ASAP7_75t_L g1454 ( 
.A1(n_1438),
.A2(n_1424),
.A3(n_1422),
.B1(n_1395),
.B2(n_1420),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1427),
.Y(n_1455)
);

NAND4xp25_ASAP7_75t_L g1456 ( 
.A(n_1443),
.B(n_1370),
.C(n_1414),
.D(n_1423),
.Y(n_1456)
);

OAI211xp5_ASAP7_75t_L g1457 ( 
.A1(n_1439),
.A2(n_1416),
.B(n_1415),
.C(n_1417),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1442),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1430),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1433),
.A2(n_1381),
.B1(n_1376),
.B2(n_1305),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1441),
.A2(n_1348),
.B(n_1366),
.C(n_1356),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1445),
.B(n_1408),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1432),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1447),
.A2(n_1394),
.B(n_1392),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1453),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1455),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1459),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1448),
.B(n_1416),
.C(n_1434),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1433),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1463),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1465),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1469),
.B(n_1454),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1469),
.A2(n_1450),
.B(n_1452),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1468),
.B(n_1448),
.C(n_1460),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1470),
.A2(n_1451),
.B(n_1456),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1475),
.B(n_1356),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1474),
.B(n_1461),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1473),
.B(n_1464),
.C(n_1466),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1472),
.B(n_1467),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1471),
.B(n_1457),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1471),
.B(n_1458),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1472),
.B(n_1462),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1471),
.Y(n_1483)
);

NOR3x1_ASAP7_75t_L g1484 ( 
.A(n_1478),
.B(n_1311),
.C(n_1303),
.Y(n_1484)
);

NOR4xp25_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1320),
.C(n_1335),
.D(n_1315),
.Y(n_1485)
);

NOR3x1_ASAP7_75t_L g1486 ( 
.A(n_1479),
.B(n_1303),
.C(n_1306),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1477),
.B(n_1435),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1482),
.B(n_1366),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1483),
.B(n_1436),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1480),
.B(n_1442),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1481),
.Y(n_1491)
);

NAND4xp75_ASAP7_75t_L g1492 ( 
.A(n_1484),
.B(n_1339),
.C(n_1340),
.D(n_1336),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_L g1493 ( 
.A(n_1488),
.B(n_1312),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1487),
.B(n_1312),
.Y(n_1494)
);

NOR2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1491),
.B(n_1317),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1490),
.B(n_1306),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1493),
.B(n_1485),
.C(n_1489),
.Y(n_1497)
);

XNOR2xp5_ASAP7_75t_L g1498 ( 
.A(n_1495),
.B(n_1326),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1494),
.B(n_1496),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1492),
.B(n_1319),
.Y(n_1500)
);

NAND4xp25_ASAP7_75t_L g1501 ( 
.A(n_1500),
.B(n_1486),
.C(n_1317),
.D(n_1316),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1499),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1497),
.B(n_1322),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1498),
.B(n_1319),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1502),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1503),
.B(n_1327),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1504),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1505),
.A2(n_1501),
.B(n_1307),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1507),
.A2(n_1440),
.B1(n_1437),
.B2(n_1406),
.Y(n_1509)
);

AOI22x1_ASAP7_75t_L g1510 ( 
.A1(n_1506),
.A2(n_1322),
.B1(n_1440),
.B2(n_1298),
.Y(n_1510)
);

AOI22x1_ASAP7_75t_L g1511 ( 
.A1(n_1508),
.A2(n_1506),
.B1(n_1298),
.B2(n_1376),
.Y(n_1511)
);

AOI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1510),
.A2(n_1342),
.B(n_1308),
.Y(n_1512)
);

AO21x1_ASAP7_75t_L g1513 ( 
.A1(n_1512),
.A2(n_1509),
.B(n_1313),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1513),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1514),
.B(n_1511),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1515),
.A2(n_1308),
.B1(n_1307),
.B2(n_1361),
.Y(n_1516)
);


endmodule