module real_aes_8133_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_715, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_715;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g155 ( .A1(n_0), .A2(n_156), .B(n_157), .C(n_161), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_1), .B(n_150), .Y(n_163) );
INVx1_ASAP7_75t_L g408 ( .A(n_2), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_3), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_4), .A2(n_124), .B(n_141), .C(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_5), .A2(n_144), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_6), .A2(n_144), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_7), .B(n_150), .Y(n_490) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_8), .A2(n_116), .B(n_203), .Y(n_202) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_10), .A2(n_124), .B(n_141), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g455 ( .A(n_11), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_12), .B(n_40), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_13), .B(n_160), .Y(n_465) );
INVx1_ASAP7_75t_L g121 ( .A(n_14), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_15), .B(n_135), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_16), .A2(n_136), .B(n_474), .C(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_17), .B(n_150), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_18), .A2(n_65), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_18), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_19), .B(n_193), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_20), .A2(n_124), .B(n_187), .C(n_192), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_21), .A2(n_159), .B(n_211), .C(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_22), .B(n_160), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_23), .B(n_160), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_24), .Y(n_493) );
INVx1_ASAP7_75t_L g505 ( .A(n_25), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_26), .A2(n_124), .B(n_192), .C(n_206), .Y(n_205) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_27), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_28), .Y(n_461) );
INVx1_ASAP7_75t_L g522 ( .A(n_29), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_30), .A2(n_144), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_32), .A2(n_139), .B(n_171), .C(n_172), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_33), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_34), .A2(n_159), .B(n_487), .C(n_489), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_35), .A2(n_103), .B1(n_414), .B2(n_422), .C1(n_424), .C2(n_709), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_35), .A2(n_105), .B1(n_400), .B2(n_401), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_35), .Y(n_400) );
INVxp67_ASAP7_75t_L g523 ( .A(n_36), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_37), .B(n_208), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g485 ( .A(n_38), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_39), .A2(n_124), .B(n_192), .C(n_504), .Y(n_503) );
AOI222xp33_ASAP7_75t_L g425 ( .A1(n_41), .A2(n_426), .B1(n_695), .B2(n_696), .C1(n_702), .C2(n_706), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_42), .A2(n_161), .B(n_453), .C(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_43), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_44), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_45), .B(n_135), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_46), .B(n_144), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_47), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_48), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_49), .A2(n_139), .B(n_171), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g158 ( .A(n_50), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_51), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_51), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_52), .A2(n_83), .B1(n_700), .B2(n_701), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_52), .Y(n_701) );
INVx1_ASAP7_75t_L g233 ( .A(n_53), .Y(n_233) );
INVx1_ASAP7_75t_L g443 ( .A(n_54), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_55), .B(n_144), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_56), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_57), .Y(n_451) );
INVx1_ASAP7_75t_L g142 ( .A(n_58), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_59), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_60), .B(n_150), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_61), .A2(n_131), .B(n_191), .C(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g120 ( .A(n_62), .Y(n_120) );
INVx1_ASAP7_75t_SL g488 ( .A(n_63), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_64), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_65), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_66), .B(n_135), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_67), .B(n_150), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_68), .B(n_136), .Y(n_222) );
INVx1_ASAP7_75t_L g496 ( .A(n_69), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_70), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_71), .B(n_175), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_72), .A2(n_124), .B(n_129), .C(n_139), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_73), .Y(n_247) );
INVx1_ASAP7_75t_L g421 ( .A(n_74), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_75), .A2(n_144), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_76), .B(n_411), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_77), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_78), .A2(n_144), .B(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_79), .A2(n_185), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g472 ( .A(n_80), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_81), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_82), .B(n_174), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_83), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_84), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_85), .A2(n_144), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g475 ( .A(n_86), .Y(n_475) );
INVx2_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
INVx1_ASAP7_75t_L g464 ( .A(n_88), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_89), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_90), .B(n_160), .Y(n_223) );
OR2x2_ASAP7_75t_L g405 ( .A(n_91), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g429 ( .A(n_91), .B(n_407), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_91), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_92), .A2(n_124), .B(n_139), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_93), .B(n_144), .Y(n_169) );
INVx1_ASAP7_75t_L g173 ( .A(n_94), .Y(n_173) );
INVxp67_ASAP7_75t_L g250 ( .A(n_95), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_96), .B(n_116), .Y(n_456) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g218 ( .A(n_98), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_99), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g446 ( .A(n_100), .Y(n_446) );
AND2x2_ASAP7_75t_L g235 ( .A(n_101), .B(n_178), .Y(n_235) );
OAI21xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_402), .B(n_410), .Y(n_103) );
INVx1_ASAP7_75t_L g401 ( .A(n_105), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx2_ASAP7_75t_L g430 ( .A(n_109), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_109), .A2(n_428), .B1(n_704), .B2(n_705), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_343), .Y(n_109) );
AND4x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_283), .C(n_298), .D(n_323), .Y(n_110) );
NOR2xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_256), .Y(n_111) );
OAI21xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_164), .B(n_236), .Y(n_112) );
AND2x2_ASAP7_75t_L g286 ( .A(n_113), .B(n_182), .Y(n_286) );
AND2x2_ASAP7_75t_L g299 ( .A(n_113), .B(n_181), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_113), .B(n_165), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_113), .Y(n_353) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_149), .Y(n_113) );
INVx2_ASAP7_75t_L g270 ( .A(n_114), .Y(n_270) );
BUFx2_ASAP7_75t_L g297 ( .A(n_114), .Y(n_297) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_122), .B(n_147), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_115), .B(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_115), .B(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_115), .A2(n_217), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_115), .B(n_468), .Y(n_467) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_115), .A2(n_492), .B(n_498), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_115), .B(n_508), .Y(n_507) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_116), .A2(n_204), .B(n_205), .Y(n_203) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_116), .Y(n_244) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g226 ( .A(n_117), .Y(n_226) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_118), .B(n_119), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_143), .Y(n_122) );
INVx5_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
BUFx3_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
INVx1_ASAP7_75t_L g212 ( .A(n_126), .Y(n_212) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_128), .Y(n_133) );
INVx3_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
AND2x2_ASAP7_75t_L g145 ( .A(n_128), .B(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
INVx1_ASAP7_75t_L g208 ( .A(n_128), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_134), .C(n_137), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_132), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_132), .B(n_475), .Y(n_474) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_132), .A2(n_135), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
INVx2_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_135), .B(n_250), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_135), .A2(n_190), .B(n_505), .C(n_506), .Y(n_504) );
INVx5_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_136), .B(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g489 ( .A(n_138), .Y(n_489) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g152 ( .A1(n_140), .A2(n_153), .B(n_154), .C(n_155), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_140), .A2(n_154), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g442 ( .A1(n_140), .A2(n_154), .B(n_443), .C(n_444), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_SL g450 ( .A1(n_140), .A2(n_154), .B(n_451), .C(n_452), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_SL g471 ( .A1(n_140), .A2(n_154), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_140), .A2(n_154), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_140), .A2(n_154), .B(n_519), .C(n_520), .Y(n_518) );
INVx4_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g144 ( .A(n_141), .B(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_141), .B(n_145), .Y(n_219) );
BUFx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx1_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
AND2x2_ASAP7_75t_L g237 ( .A(n_149), .B(n_182), .Y(n_237) );
INVx2_ASAP7_75t_L g253 ( .A(n_149), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_149), .B(n_181), .Y(n_262) );
AND2x2_ASAP7_75t_L g341 ( .A(n_149), .B(n_270), .Y(n_341) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_163), .Y(n_149) );
INVx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_159), .B(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g453 ( .A(n_160), .Y(n_453) );
INVx2_ASAP7_75t_L g466 ( .A(n_161), .Y(n_466) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx1_ASAP7_75t_L g476 ( .A(n_162), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_198), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_165), .B(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g394 ( .A(n_165), .Y(n_394) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_181), .Y(n_165) );
AND2x2_ASAP7_75t_L g252 ( .A(n_166), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g266 ( .A(n_166), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_166), .Y(n_295) );
OR2x2_ASAP7_75t_L g327 ( .A(n_166), .B(n_269), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_166), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g368 ( .A(n_166), .B(n_337), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_166), .B(n_237), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_166), .B(n_297), .Y(n_393) );
AND2x2_ASAP7_75t_L g399 ( .A(n_166), .B(n_286), .Y(n_399) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx2_ASAP7_75t_L g259 ( .A(n_167), .Y(n_259) );
AND2x2_ASAP7_75t_L g289 ( .A(n_167), .B(n_269), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_167), .B(n_282), .Y(n_322) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_182), .Y(n_342) );
AND2x2_ASAP7_75t_L g376 ( .A(n_167), .B(n_242), .Y(n_376) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_179), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_178), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_176), .C(n_177), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_174), .A2(n_177), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp5_ASAP7_75t_L g463 ( .A1(n_174), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_174), .A2(n_466), .B(n_496), .C(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_178), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_178), .A2(n_230), .B(n_231), .Y(n_229) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_178), .A2(n_449), .B(n_456), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_178), .A2(n_219), .B(n_502), .C(n_503), .Y(n_501) );
AND2x4_ASAP7_75t_L g282 ( .A(n_181), .B(n_253), .Y(n_282) );
AND2x2_ASAP7_75t_L g293 ( .A(n_181), .B(n_289), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_181), .B(n_269), .Y(n_332) );
INVx2_ASAP7_75t_L g347 ( .A(n_181), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_181), .B(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_181), .B(n_341), .Y(n_389) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_182), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g337 ( .A(n_182), .B(n_253), .Y(n_337) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_195), .Y(n_182) );
AOI21xp5_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_186), .B(n_193), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_191), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_194), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_197), .A2(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x2_ASAP7_75t_L g260 ( .A(n_200), .B(n_243), .Y(n_260) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_201), .B(n_216), .Y(n_240) );
OR2x2_ASAP7_75t_L g273 ( .A(n_201), .B(n_243), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_201), .B(n_243), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_201), .B(n_242), .Y(n_305) );
AND2x2_ASAP7_75t_L g357 ( .A(n_201), .B(n_215), .Y(n_357) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_202), .B(n_227), .Y(n_265) );
AND2x2_ASAP7_75t_L g301 ( .A(n_202), .B(n_216), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_210), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_210), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_213), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g291 ( .A(n_214), .B(n_273), .Y(n_291) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_227), .Y(n_214) );
OAI322xp33_ASAP7_75t_L g256 ( .A1(n_215), .A2(n_257), .A3(n_261), .B1(n_263), .B2(n_266), .C1(n_271), .C2(n_279), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_215), .B(n_242), .Y(n_264) );
OR2x2_ASAP7_75t_L g274 ( .A(n_215), .B(n_228), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_215), .B(n_228), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_215), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_215), .B(n_243), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_215), .B(n_372), .Y(n_371) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_216), .B(n_260), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_219), .A2(n_461), .B(n_462), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_219), .A2(n_493), .B(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g516 ( .A(n_226), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_227), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_227), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g316 ( .A(n_227), .B(n_243), .Y(n_316) );
AOI211xp5_ASAP7_75t_SL g344 ( .A1(n_227), .A2(n_345), .B(n_348), .C(n_360), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_227), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g382 ( .A(n_227), .B(n_357), .Y(n_382) );
INVx5_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g310 ( .A(n_228), .B(n_243), .Y(n_310) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_228), .Y(n_319) );
AND2x2_ASAP7_75t_L g359 ( .A(n_228), .B(n_357), .Y(n_359) );
AND2x2_ASAP7_75t_SL g390 ( .A(n_228), .B(n_260), .Y(n_390) );
AND2x2_ASAP7_75t_L g397 ( .A(n_228), .B(n_356), .Y(n_397) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B1(n_252), .B2(n_254), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_237), .B(n_259), .Y(n_307) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g255 ( .A(n_240), .Y(n_255) );
OR2x2_ASAP7_75t_L g315 ( .A(n_240), .B(n_316), .Y(n_315) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_240), .A2(n_364), .B1(n_366), .B2(n_367), .C(n_369), .Y(n_363) );
INVx2_ASAP7_75t_L g302 ( .A(n_241), .Y(n_302) );
AND2x2_ASAP7_75t_L g275 ( .A(n_242), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g365 ( .A(n_242), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_242), .B(n_357), .Y(n_378) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g320 ( .A(n_243), .Y(n_320) );
AND2x2_ASAP7_75t_L g356 ( .A(n_243), .B(n_357), .Y(n_356) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_244), .A2(n_441), .B(n_447), .Y(n_440) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_244), .A2(n_470), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_244), .A2(n_483), .B(n_490), .Y(n_482) );
AND2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_297), .Y(n_358) );
AND2x2_ASAP7_75t_L g268 ( .A(n_253), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_253), .B(n_326), .Y(n_325) );
NOR2xp33_ASAP7_75t_SL g339 ( .A(n_255), .B(n_302), .Y(n_339) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g345 ( .A(n_258), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OR2x2_ASAP7_75t_L g331 ( .A(n_259), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g396 ( .A(n_259), .B(n_341), .Y(n_396) );
INVx2_ASAP7_75t_L g329 ( .A(n_260), .Y(n_329) );
NAND4xp25_ASAP7_75t_SL g392 ( .A(n_261), .B(n_393), .C(n_394), .D(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_262), .B(n_326), .Y(n_361) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx1_ASAP7_75t_SL g398 ( .A(n_265), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_SL g360 ( .A1(n_266), .A2(n_329), .B(n_333), .C(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g355 ( .A(n_268), .B(n_347), .Y(n_355) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_270), .Y(n_313) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_275), .C(n_277), .Y(n_271) );
AND2x2_ASAP7_75t_L g292 ( .A(n_272), .B(n_276), .Y(n_292) );
OAI322xp33_ASAP7_75t_SL g330 ( .A1(n_272), .A2(n_331), .A3(n_333), .B1(n_334), .B2(n_338), .C1(n_339), .C2(n_340), .Y(n_330) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g352 ( .A(n_274), .B(n_278), .Y(n_352) );
INVx1_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
INVx1_ASAP7_75t_SL g351 ( .A(n_278), .Y(n_351) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AOI222xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_290), .B1(n_292), .B2(n_293), .C1(n_294), .C2(n_715), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_285), .A2(n_347), .A3(n_352), .B1(n_374), .B2(n_375), .C1(n_377), .C2(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_300), .B1(n_324), .B2(n_328), .C(n_330), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OAI222xp33_ASAP7_75t_L g303 ( .A1(n_291), .A2(n_304), .B1(n_306), .B2(n_307), .C1(n_308), .C2(n_311), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_293), .A2(n_300), .B1(n_370), .B2(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .C(n_314), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g379 ( .A1(n_300), .A2(n_337), .B(n_380), .C(n_383), .Y(n_379) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_301), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g372 ( .A(n_305), .Y(n_372) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_312), .B(n_337), .Y(n_366) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_321), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_315), .A2(n_384), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_383) );
INVxp33_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_326), .B(n_337), .Y(n_377) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g388 ( .A(n_341), .B(n_347), .Y(n_388) );
AND4x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_362), .C(n_379), .D(n_391), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_350), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_359), .Y(n_354) );
INVx1_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
INVx1_ASAP7_75t_SL g374 ( .A(n_359), .Y(n_374) );
NOR2xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_375), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_382), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_397), .B1(n_398), .B2(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g413 ( .A(n_405), .Y(n_413) );
INVx1_ASAP7_75t_SL g713 ( .A(n_405), .Y(n_713) );
NOR2x2_ASAP7_75t_L g708 ( .A(n_406), .B(n_433), .Y(n_708) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g432 ( .A(n_407), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OA21x2_ASAP7_75t_L g423 ( .A1(n_413), .A2(n_418), .B(n_419), .Y(n_423) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g711 ( .A(n_418), .B(n_420), .Y(n_711) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_431), .B2(n_434), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx6_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g704 ( .A(n_432), .Y(n_704) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g705 ( .A(n_435), .Y(n_705) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_621), .Y(n_435) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_437), .B(n_563), .C(n_593), .D(n_603), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_478), .B(n_526), .C(n_553), .Y(n_437) );
OAI222xp33_ASAP7_75t_L g648 ( .A1(n_438), .A2(n_568), .B1(n_649), .B2(n_650), .C1(n_651), .C2(n_652), .Y(n_648) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_457), .Y(n_438) );
AOI33xp33_ASAP7_75t_L g574 ( .A1(n_439), .A2(n_561), .A3(n_562), .B1(n_575), .B2(n_580), .B3(n_582), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g631 ( .A1(n_439), .A2(n_632), .B(n_634), .C(n_636), .Y(n_631) );
OR2x2_ASAP7_75t_L g647 ( .A(n_439), .B(n_633), .Y(n_647) );
INVx1_ASAP7_75t_L g680 ( .A(n_439), .Y(n_680) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_448), .Y(n_439) );
INVx2_ASAP7_75t_L g557 ( .A(n_440), .Y(n_557) );
AND2x2_ASAP7_75t_L g573 ( .A(n_440), .B(n_469), .Y(n_573) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_440), .Y(n_608) );
AND2x2_ASAP7_75t_L g637 ( .A(n_440), .B(n_448), .Y(n_637) );
INVx2_ASAP7_75t_L g537 ( .A(n_448), .Y(n_537) );
BUFx3_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_448), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g556 ( .A(n_448), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_448), .B(n_458), .Y(n_585) );
AND2x2_ASAP7_75t_L g654 ( .A(n_448), .B(n_588), .Y(n_654) );
INVx2_ASAP7_75t_SL g548 ( .A(n_457), .Y(n_548) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_469), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_458), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g590 ( .A(n_458), .Y(n_590) );
AND2x2_ASAP7_75t_L g601 ( .A(n_458), .B(n_557), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_458), .B(n_586), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_458), .B(n_588), .Y(n_633) );
AND2x2_ASAP7_75t_L g692 ( .A(n_458), .B(n_637), .Y(n_692) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g562 ( .A(n_459), .B(n_469), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_459), .B(n_573), .Y(n_572) );
BUFx3_ASAP7_75t_L g594 ( .A(n_459), .Y(n_594) );
AND3x2_ASAP7_75t_L g653 ( .A(n_459), .B(n_654), .C(n_655), .Y(n_653) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_469), .Y(n_544) );
INVx1_ASAP7_75t_SL g588 ( .A(n_469), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_469), .B(n_537), .C(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_509), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_479), .A2(n_572), .B(n_624), .C(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_481), .B(n_500), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_481), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g640 ( .A(n_481), .Y(n_640) );
AND2x2_ASAP7_75t_L g661 ( .A(n_481), .B(n_511), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_481), .B(n_570), .Y(n_689) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
AND2x2_ASAP7_75t_L g534 ( .A(n_482), .B(n_525), .Y(n_534) );
INVx2_ASAP7_75t_L g541 ( .A(n_482), .Y(n_541) );
AND2x2_ASAP7_75t_L g561 ( .A(n_482), .B(n_511), .Y(n_561) );
AND2x2_ASAP7_75t_L g611 ( .A(n_482), .B(n_500), .Y(n_611) );
INVx1_ASAP7_75t_L g615 ( .A(n_482), .Y(n_615) );
INVx2_ASAP7_75t_SL g525 ( .A(n_491), .Y(n_525) );
BUFx2_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
AND2x2_ASAP7_75t_L g678 ( .A(n_491), .B(n_500), .Y(n_678) );
INVx3_ASAP7_75t_SL g511 ( .A(n_500), .Y(n_511) );
AND2x2_ASAP7_75t_L g533 ( .A(n_500), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g540 ( .A(n_500), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g570 ( .A(n_500), .B(n_530), .Y(n_570) );
OR2x2_ASAP7_75t_L g579 ( .A(n_500), .B(n_525), .Y(n_579) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_500), .Y(n_597) );
AND2x2_ASAP7_75t_L g602 ( .A(n_500), .B(n_555), .Y(n_602) );
AND2x2_ASAP7_75t_L g630 ( .A(n_500), .B(n_513), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_500), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g668 ( .A(n_500), .B(n_512), .Y(n_668) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g592 ( .A(n_511), .B(n_541), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_511), .B(n_534), .Y(n_620) );
AND2x2_ASAP7_75t_L g638 ( .A(n_511), .B(n_555), .Y(n_638) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .Y(n_512) );
AND2x2_ASAP7_75t_L g539 ( .A(n_513), .B(n_525), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_513), .B(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g577 ( .A(n_513), .Y(n_577) );
OR2x2_ASAP7_75t_L g625 ( .A(n_513), .B(n_545), .Y(n_625) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_517), .B(n_524), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_515), .A2(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g531 ( .A(n_517), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_524), .Y(n_532) );
AND2x2_ASAP7_75t_L g560 ( .A(n_525), .B(n_530), .Y(n_560) );
INVx1_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
AND2x2_ASAP7_75t_L g663 ( .A(n_525), .B(n_541), .Y(n_663) );
AOI222xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_535), .B1(n_538), .B2(n_542), .C1(n_546), .C2(n_549), .Y(n_526) );
INVx1_ASAP7_75t_L g658 ( .A(n_527), .Y(n_658) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AND2x2_ASAP7_75t_L g554 ( .A(n_528), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g565 ( .A(n_528), .B(n_534), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_528), .B(n_556), .Y(n_581) );
OAI222xp33_ASAP7_75t_L g603 ( .A1(n_528), .A2(n_604), .B1(n_609), .B2(n_610), .C1(n_618), .C2(n_620), .Y(n_603) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g591 ( .A(n_530), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_530), .B(n_611), .Y(n_651) );
AND2x2_ASAP7_75t_L g662 ( .A(n_530), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_533), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_535), .B(n_586), .Y(n_649) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_537), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx3_ASAP7_75t_L g552 ( .A(n_540), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_540), .A2(n_643), .B(n_646), .C(n_648), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_540), .B(n_577), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_540), .B(n_560), .Y(n_682) );
AND2x2_ASAP7_75t_L g555 ( .A(n_541), .B(n_551), .Y(n_555) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_545), .B(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g634 ( .A(n_545), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g673 ( .A(n_545), .B(n_573), .Y(n_673) );
INVx1_ASAP7_75t_L g685 ( .A(n_545), .Y(n_685) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_548), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g666 ( .A(n_551), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_556), .B(n_558), .C(n_562), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_554), .A2(n_584), .B1(n_599), .B2(n_602), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_555), .B(n_569), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_555), .B(n_577), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_556), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g619 ( .A(n_556), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_556), .B(n_606), .Y(n_626) );
INVx2_ASAP7_75t_L g587 ( .A(n_557), .Y(n_587) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NOR4xp25_ASAP7_75t_L g564 ( .A(n_561), .B(n_565), .C(n_566), .D(n_569), .Y(n_564) );
INVx1_ASAP7_75t_SL g635 ( .A(n_562), .Y(n_635) );
AND2x2_ASAP7_75t_L g679 ( .A(n_562), .B(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g563 ( .A1(n_564), .A2(n_571), .B(n_574), .C(n_583), .Y(n_563) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_570), .B(n_640), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_572), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
INVx1_ASAP7_75t_SL g645 ( .A(n_573), .Y(n_645) );
AND2x2_ASAP7_75t_L g684 ( .A(n_573), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_577), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_581), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_582), .B(n_607), .Y(n_667) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_589), .B(n_591), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g659 ( .A(n_586), .Y(n_659) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g687 ( .A(n_587), .Y(n_687) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_598), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g606 ( .A(n_594), .Y(n_606) );
OR2x2_ASAP7_75t_L g644 ( .A(n_594), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g639 ( .A1(n_597), .A2(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_601), .A2(n_628), .B1(n_631), .B2(n_638), .C(n_639), .Y(n_627) );
INVx1_ASAP7_75t_SL g671 ( .A(n_602), .Y(n_671) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OR2x2_ASAP7_75t_L g618 ( .A(n_606), .B(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_L g655 ( .A(n_608), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_615), .B2(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g650 ( .A(n_611), .Y(n_650) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_614), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_656), .C(n_669), .D(n_681), .Y(n_621) );
NAND3xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_627), .C(n_642), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_625), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_632), .B(n_637), .Y(n_641) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI221xp5_ASAP7_75t_SL g669 ( .A1(n_644), .A2(n_670), .B1(n_671), .B2(n_672), .C(n_674), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_646), .A2(n_661), .B(n_662), .C(n_664), .Y(n_660) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_647), .A2(n_665), .B1(n_667), .B2(n_668), .Y(n_664) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B(n_659), .C(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g675 ( .A(n_668), .Y(n_675) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B1(n_686), .B2(n_688), .C(n_690), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx3_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
endmodule