module real_jpeg_6091_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_0),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_0),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_0),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_0),
.B(n_117),
.Y(n_188)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_2),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_135),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_2),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_2),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_2),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_2),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_3),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_246),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_4),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_4),
.Y(n_382)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_6),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_6),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

BUFx5_ASAP7_75t_L g408 ( 
.A(n_7),
.Y(n_408)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_8),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_9),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_9),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_9),
.B(n_129),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_9),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_9),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_9),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_9),
.B(n_385),
.Y(n_384)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_11),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_12),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_12),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_12),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_12),
.B(n_222),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_12),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_13),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_13),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_13),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_13),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_14),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_14),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_14),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_14),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_14),
.B(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_207),
.B1(n_452),
.B2(n_453),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_18),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_206),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_177),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_21),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.C(n_145),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_22),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.C(n_90),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_23),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.C(n_54),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_24),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_28),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_27),
.A2(n_28),
.B1(n_346),
.B2(n_347),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_30),
.C(n_36),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_28),
.B(n_154),
.C(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_28),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_30),
.A2(n_35),
.B1(n_232),
.B2(n_233),
.Y(n_318)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_33),
.Y(n_405)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g349 ( 
.A(n_34),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_36),
.A2(n_40),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_38),
.Y(n_317)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_39),
.Y(n_141)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_39),
.Y(n_263)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_39),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_41),
.B(n_54),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.C(n_50),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_42),
.B(n_50),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_44),
.Y(n_219)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_45),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_46),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_50),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_50),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_52),
.Y(n_361)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_53),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_55),
.Y(n_152)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_66),
.C(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_65),
.Y(n_354)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_71),
.B(n_90),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.C(n_86),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_73),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.C(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_74),
.A2(n_75),
.B1(n_81),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_75),
.B(n_110),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_75),
.B(n_110),
.Y(n_355)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_77),
.Y(n_274)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_77),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_78),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_78),
.Y(n_238)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_116),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_80),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_81),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_83),
.B(n_86),
.Y(n_295)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_99),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_97),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_97),
.A2(n_99),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_99),
.B(n_169),
.C(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_101),
.B(n_145),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_119),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_102),
.B(n_120),
.C(n_132),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_103),
.A2(n_104),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_103),
.A2(n_104),
.B1(n_227),
.B2(n_305),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_104),
.B(n_110),
.C(n_115),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_104),
.B(n_226),
.C(n_227),
.Y(n_225)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_118),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_110),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_121),
.C(n_127),
.Y(n_120)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_126),
.Y(n_309)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_131),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_138),
.B2(n_144),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_134),
.B(n_139),
.C(n_143),
.Y(n_193)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_165),
.B2(n_166),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_167),
.C(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_148),
.B(n_151),
.Y(n_330)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_153),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_154),
.A2(n_163),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_154),
.B(n_257),
.C(n_261),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_158),
.Y(n_398)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_191),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_184),
.B1(n_216),
.B2(n_220),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_184),
.B(n_216),
.C(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_207),
.Y(n_453)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_335),
.B(n_338),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_325),
.B(n_334),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_296),
.B(n_324),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_210),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_285),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_211),
.B(n_285),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_255),
.C(n_279),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_212),
.B(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_236),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_213),
.B(n_237),
.C(n_242),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_225),
.C(n_230),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_214),
.B(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_225),
.A2(n_230),
.B1(n_231),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_225),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_226),
.B(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_242),
.Y(n_455)
);

FAx1_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.CI(n_252),
.CON(n_242),
.SN(n_242)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_247),
.C(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.C(n_267),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_265),
.B1(n_266),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_258),
.B(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_258),
.B(n_398),
.Y(n_418)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.C(n_275),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_268),
.A2(n_269),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_270),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_440)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_273),
.Y(n_385)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_322),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_297),
.B(n_322),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.C(n_319),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_298),
.A2(n_299),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_302),
.B(n_319),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_318),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_303),
.B(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_306),
.B(n_318),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.C(n_313),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_314),
.B(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_326),
.B(n_335),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_336),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_328),
.B(n_336),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_331),
.CI(n_333),
.CON(n_328),
.SN(n_328)
);

OAI31xp33_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_448),
.A3(n_449),
.B(n_451),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_442),
.B(n_447),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_429),
.B(n_441),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_387),
.B(n_428),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_373),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_373),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_356),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_344),
.B(n_357),
.C(n_370),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_351),
.C(n_355),
.Y(n_437)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx8_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_370),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.C(n_367),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_358),
.B(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_362),
.A2(n_363),
.B1(n_367),
.B2(n_368),
.Y(n_375)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.C(n_386),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_377),
.B1(n_386),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_383),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_379),
.B1(n_383),
.B2(n_384),
.Y(n_399)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_422),
.B(n_427),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_409),
.B(n_421),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_400),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_400),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_399),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_396),
.C(n_399),
.Y(n_423)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_406),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_401),
.A2(n_402),
.B1(n_406),
.B2(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_417),
.B(n_420),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_414),
.Y(n_410)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_419),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_424),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_431),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_436),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_437),
.C(n_438),
.Y(n_446)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_446),
.Y(n_447)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_444),
.Y(n_445)
);


endmodule