module fake_jpeg_28924_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_26),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_56),
.Y(n_115)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_58),
.B(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_86),
.Y(n_111)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_32),
.Y(n_77)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_87),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_89),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_51),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_40),
.B(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_14),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_97),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_24),
.B(n_51),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_18),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_96),
.Y(n_139)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_110),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_139),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_42),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_25),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

CKINVDCx6p67_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_102),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_39),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_36),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_158),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_39),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_46),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_70),
.B(n_28),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_163),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_170),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_77),
.B1(n_64),
.B2(n_61),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_172),
.B1(n_213),
.B2(n_223),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_85),
.B1(n_100),
.B2(n_73),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_174),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_13),
.B(n_14),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_177),
.B(n_194),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_66),
.B(n_54),
.C(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_178),
.B(n_179),
.Y(n_244)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

CKINVDCx12_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_67),
.B1(n_101),
.B2(n_81),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_189),
.A2(n_196),
.B1(n_155),
.B2(n_121),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_191),
.Y(n_273)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_136),
.B(n_105),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_134),
.A2(n_63),
.B1(n_91),
.B2(n_69),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_116),
.A2(n_76),
.B1(n_92),
.B2(n_82),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_215),
.B1(n_224),
.B2(n_125),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_47),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_216),
.Y(n_227)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_127),
.B(n_0),
.C(n_1),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_116),
.B(n_78),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_218),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_108),
.A2(n_79),
.B(n_75),
.C(n_93),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_212),
.A2(n_219),
.B(n_151),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_151),
.A2(n_28),
.B1(n_47),
.B2(n_46),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_126),
.A2(n_53),
.B1(n_45),
.B2(n_38),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_220),
.B1(n_222),
.B2(n_226),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_138),
.B(n_45),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_117),
.A2(n_45),
.B1(n_32),
.B2(n_38),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_34),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_126),
.A2(n_38),
.B1(n_32),
.B2(n_50),
.Y(n_224)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_109),
.B1(n_141),
.B2(n_165),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_228),
.B(n_230),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_129),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_231),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_135),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_109),
.B(n_110),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_237),
.A2(n_203),
.B(n_185),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_224),
.B1(n_218),
.B2(n_178),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_249),
.B1(n_254),
.B2(n_258),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_179),
.A2(n_155),
.B1(n_120),
.B2(n_121),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_159),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_250),
.B(n_268),
.C(n_204),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_165),
.B1(n_157),
.B2(n_117),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_196),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_216),
.A2(n_113),
.B1(n_164),
.B2(n_140),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_261),
.A2(n_269),
.B(n_171),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_176),
.B(n_162),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_234),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_189),
.A2(n_113),
.B1(n_164),
.B2(n_47),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_267),
.A2(n_272),
.B1(n_203),
.B2(n_214),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_153),
.C(n_140),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_172),
.A2(n_153),
.B1(n_197),
.B2(n_208),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_168),
.A2(n_47),
.B1(n_46),
.B2(n_28),
.Y(n_272)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_238),
.B1(n_260),
.B2(n_233),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_275),
.A2(n_262),
.B1(n_235),
.B2(n_251),
.Y(n_349)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_212),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_278),
.B(n_280),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_174),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_281),
.B(n_284),
.Y(n_334)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_282),
.Y(n_322)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_312),
.B(n_237),
.Y(n_315)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_183),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_290),
.B(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_292),
.Y(n_340)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_184),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_229),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_313),
.B1(n_262),
.B2(n_241),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_214),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_298),
.A2(n_305),
.B(n_227),
.C(n_213),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_232),
.B(n_225),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_299),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_258),
.B(n_230),
.Y(n_323)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_271),
.Y(n_302)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_247),
.B(n_46),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_307),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_214),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_242),
.B(n_1),
.Y(n_307)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_308),
.Y(n_321)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_311),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_310),
.B(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_345),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_323),
.A2(n_329),
.B(n_343),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_247),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_327),
.B(n_346),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_268),
.C(n_232),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_332),
.C(n_336),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_242),
.C(n_265),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_279),
.A2(n_254),
.B1(n_239),
.B2(n_267),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_306),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_248),
.B(n_235),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_255),
.B(n_241),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_248),
.C(n_271),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_281),
.B(n_255),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_276),
.C(n_285),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_348),
.B(n_302),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_279),
.B1(n_287),
.B2(n_295),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_353),
.B1(n_371),
.B2(n_377),
.Y(n_393)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_374),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_318),
.B(n_294),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_358),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_323),
.A2(n_306),
.B1(n_287),
.B2(n_289),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_307),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_354),
.B(n_355),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_293),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_357),
.A2(n_329),
.B1(n_326),
.B2(n_317),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_360),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_321),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_368),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_338),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_363),
.B(n_373),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_316),
.A2(n_300),
.B1(n_288),
.B2(n_296),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_364),
.A2(n_333),
.B(n_330),
.Y(n_407)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_334),
.B(n_292),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_328),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_291),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_372),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_297),
.B1(n_278),
.B2(n_305),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_341),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_283),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_341),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_375),
.A2(n_319),
.B1(n_324),
.B2(n_344),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_347),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_326),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_315),
.A2(n_311),
.B1(n_301),
.B2(n_313),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_304),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_381),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_265),
.C(n_264),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_264),
.C(n_236),
.Y(n_410)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_333),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_387),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_346),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_384),
.A2(n_378),
.B(n_380),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_336),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_329),
.B(n_335),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_404),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_368),
.B(n_337),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_390),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_329),
.C(n_344),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_395),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_329),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_220),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_351),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_401),
.A2(n_407),
.B(n_411),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_319),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_403),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_282),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_358),
.A2(n_324),
.B1(n_317),
.B2(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_379),
.C(n_375),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_362),
.A2(n_274),
.B(n_308),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_304),
.B1(n_309),
.B2(n_286),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_412),
.A2(n_361),
.B1(n_372),
.B2(n_374),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_414),
.A2(n_423),
.B(n_1),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g415 ( 
.A(n_396),
.B(n_362),
.CI(n_377),
.CON(n_415),
.SN(n_415)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_431),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_427),
.C(n_433),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_422),
.B1(n_424),
.B2(n_432),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_362),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_437),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_393),
.A2(n_352),
.B1(n_375),
.B2(n_365),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_391),
.A2(n_365),
.B(n_361),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_350),
.B1(n_370),
.B2(n_381),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_410),
.C(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_398),
.Y(n_428)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_382),
.B(n_367),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_430),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_360),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_170),
.B1(n_190),
.B2(n_217),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_246),
.C(n_245),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_434),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_386),
.B(n_401),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_409),
.A2(n_351),
.B1(n_245),
.B2(n_236),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_408),
.B1(n_406),
.B2(n_400),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_246),
.C(n_220),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_400),
.C(n_408),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_399),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_446),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_431),
.Y(n_443)
);

INVx13_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_419),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_425),
.A2(n_391),
.B1(n_399),
.B2(n_412),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_452),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_389),
.Y(n_450)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_453),
.C(n_454),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_390),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_404),
.C(n_388),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_407),
.C(n_402),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_455),
.A2(n_413),
.B1(n_438),
.B2(n_433),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_426),
.A2(n_384),
.B1(n_406),
.B2(n_405),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_415),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_417),
.B(n_389),
.C(n_41),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_421),
.C(n_415),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_459),
.A2(n_420),
.B(n_432),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_423),
.B(n_414),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_461),
.A2(n_2),
.B(n_3),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_425),
.B1(n_429),
.B2(n_420),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_463),
.A2(n_445),
.B1(n_449),
.B2(n_444),
.Y(n_484)
);

AO22x1_ASAP7_75t_L g466 ( 
.A1(n_450),
.A2(n_443),
.B1(n_448),
.B2(n_428),
.Y(n_466)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_466),
.B(n_2),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_437),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_470),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_468),
.B(n_469),
.Y(n_487)
);

AOI221xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_418),
.B1(n_413),
.B2(n_422),
.C(n_424),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_2),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_473),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_439),
.B(n_456),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_456),
.CI(n_453),
.CON(n_476),
.SN(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_476),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_463),
.A2(n_459),
.B1(n_447),
.B2(n_454),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_480),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_440),
.Y(n_478)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_472),
.CI(n_468),
.CON(n_479),
.SN(n_479)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_475),
.Y(n_498)
);

MAJx2_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_458),
.C(n_442),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_442),
.C(n_451),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_482),
.B(n_484),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_485),
.B(n_486),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_41),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g493 ( 
.A1(n_488),
.A2(n_469),
.B(n_466),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_475),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_34),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_464),
.C(n_470),
.Y(n_496)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_502),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_501),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_465),
.B(n_466),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_499),
.A2(n_477),
.B1(n_489),
.B2(n_479),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_460),
.C(n_465),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_481),
.A2(n_460),
.B(n_475),
.Y(n_502)
);

FAx1_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_483),
.CI(n_476),
.CON(n_503),
.SN(n_503)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_509),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_497),
.A2(n_485),
.B1(n_489),
.B2(n_483),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_505),
.B(n_498),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_480),
.C(n_490),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_504),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_511),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_507),
.A2(n_494),
.B(n_502),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_513),
.C(n_5),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_495),
.C(n_491),
.Y(n_513)
);

A2O1A1O1Ixp25_ASAP7_75t_L g517 ( 
.A1(n_515),
.A2(n_508),
.B(n_503),
.C(n_7),
.D(n_9),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g519 ( 
.A1(n_517),
.A2(n_514),
.B(n_7),
.Y(n_519)
);

AO21x1_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_6),
.B(n_7),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_519),
.B(n_520),
.Y(n_521)
);

AOI322xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_516),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_9),
.C2(n_41),
.Y(n_522)
);

OAI31xp33_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_11),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_41),
.Y(n_525)
);


endmodule