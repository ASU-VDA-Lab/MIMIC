module fake_jpeg_24764_n_41 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_41);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

HAxp5_ASAP7_75t_SL g20 ( 
.A(n_13),
.B(n_17),
.CON(n_20),
.SN(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_14),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_5),
.B1(n_16),
.B2(n_15),
.Y(n_25)
);

AOI22x1_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_2),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.C(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_32),
.B1(n_35),
.B2(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_27),
.B1(n_3),
.B2(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_3),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_4),
.C(n_6),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_12),
.B(n_18),
.Y(n_41)
);


endmodule