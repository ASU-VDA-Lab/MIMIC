module fake_jpeg_25302_n_273 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_33),
.B1(n_35),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_33),
.B1(n_35),
.B2(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_27),
.B1(n_32),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_62),
.B1(n_65),
.B2(n_28),
.Y(n_82)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_26),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_67),
.A2(n_69),
.B(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_0),
.B(n_2),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_27),
.A3(n_26),
.B1(n_19),
.B2(n_34),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_71),
.A2(n_91),
.B1(n_97),
.B2(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_85),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_12),
.B(n_13),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_83),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_0),
.Y(n_80)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_88),
.CI(n_90),
.CON(n_110),
.SN(n_110)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_82),
.A2(n_99),
.B1(n_16),
.B2(n_14),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_86),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_28),
.C(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_3),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_21),
.C(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_4),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_5),
.C(n_6),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_7),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_12),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_49),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_8),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_11),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_80),
.Y(n_133)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_113),
.Y(n_151)
);

OAI22x1_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_48),
.B1(n_45),
.B2(n_46),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_121),
.B1(n_91),
.B2(n_102),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_101),
.B1(n_77),
.B2(n_87),
.Y(n_152)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_87),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_14),
.B1(n_15),
.B2(n_82),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_95),
.B1(n_77),
.B2(n_76),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_143),
.B1(n_152),
.B2(n_154),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_74),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_137),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_88),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_104),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_67),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_148),
.C(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_79),
.C(n_83),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_92),
.B(n_94),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_94),
.B1(n_127),
.B2(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_152),
.B1(n_154),
.B2(n_147),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_121),
.B1(n_105),
.B2(n_123),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_185),
.B1(n_135),
.B2(n_118),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_110),
.C(n_115),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_184),
.C(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_179),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_159),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_140),
.B(n_151),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_110),
.C(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_189),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_196),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_193),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_195),
.C(n_200),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_205),
.C(n_174),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_133),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_145),
.B(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_137),
.C(n_145),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_186),
.A2(n_141),
.B1(n_153),
.B2(n_127),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_174),
.B1(n_170),
.B2(n_180),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_140),
.B1(n_120),
.B2(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_107),
.B1(n_117),
.B2(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_171),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_216),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_168),
.B(n_187),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_221),
.B(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_214),
.B1(n_224),
.B2(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_193),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_167),
.B1(n_165),
.B2(n_162),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_219),
.A2(n_222),
.B1(n_198),
.B2(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_168),
.B1(n_173),
.B2(n_176),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_161),
.B(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_200),
.C(n_198),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_234),
.C(n_237),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_201),
.B(n_190),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_229),
.B(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_164),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_238),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_191),
.C(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_210),
.B1(n_205),
.B2(n_163),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_216),
.C(n_219),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_208),
.B(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_179),
.B1(n_182),
.B2(n_163),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_239),
.A2(n_212),
.B1(n_215),
.B2(n_217),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_233),
.B1(n_236),
.B2(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_239),
.B1(n_237),
.B2(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_210),
.C(n_117),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_226),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_241),
.B(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_256),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_227),
.B(n_231),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_246),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_227),
.B1(n_232),
.B2(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_242),
.C(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_261),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_242),
.C(n_244),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_255),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_251),
.CI(n_249),
.CON(n_264),
.SN(n_264)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_268),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_263),
.B(n_265),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_252),
.B1(n_244),
.B2(n_223),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_264),
.C(n_113),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_126),
.B(n_269),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_126),
.Y(n_273)
);


endmodule