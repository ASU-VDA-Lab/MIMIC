module fake_jpeg_15109_n_120 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_5),
.B(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_2),
.B(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_26),
.Y(n_27)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_17),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AO22x2_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_6),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_22),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_15),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_20),
.B1(n_19),
.B2(n_40),
.Y(n_65)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_7),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_54),
.B1(n_9),
.B2(n_11),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_9),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_14),
.B(n_24),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_11),
.B(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_21),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_30),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_64),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_14),
.C(n_24),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_71),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_71),
.B(n_75),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_19),
.B(n_10),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_13),
.B1(n_60),
.B2(n_54),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_63),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_48),
.C(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_94),
.C(n_79),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_R g104 ( 
.A(n_92),
.B(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_64),
.C(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.C(n_103),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_65),
.B1(n_75),
.B2(n_69),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_104),
.B1(n_73),
.B2(n_66),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_81),
.C(n_93),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_104),
.B(n_96),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_86),
.C(n_83),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_70),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_70),
.A3(n_66),
.B1(n_61),
.B2(n_45),
.C1(n_59),
.C2(n_58),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_78),
.C(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_102),
.B1(n_98),
.B2(n_103),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_66),
.B(n_99),
.C(n_84),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_50),
.A3(n_56),
.B1(n_58),
.B2(n_113),
.C1(n_112),
.C2(n_114),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_105),
.B(n_45),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.C(n_114),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);


endmodule