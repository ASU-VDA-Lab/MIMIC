module fake_netlist_6_2279_n_1028 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1028);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1028;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_261;
wire n_527;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_89),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_99),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_101),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_29),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_66),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_106),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_44),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_122),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_20),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_68),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_56),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_224),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_87),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_100),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_166),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_119),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_86),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_144),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_41),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_125),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_65),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_194),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_3),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_197),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_10),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_156),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_93),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_150),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_17),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_96),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_14),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_84),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_5),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_108),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_80),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_189),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_217),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_1),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_141),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_226),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_103),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_179),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_25),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_24),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_196),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_116),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_27),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_72),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_147),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_195),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_160),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_176),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_152),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_161),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_168),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_102),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_17),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_182),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_129),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_146),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_155),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_35),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_33),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_127),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_153),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_149),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_131),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_178),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_30),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_256),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_228),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_233),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_245),
.B(n_0),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_229),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_243),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_307),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_231),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_232),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_318),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_235),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_238),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_239),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_241),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_246),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_262),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_271),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_272),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_240),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_250),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_251),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_282),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_245),
.B(n_1),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_230),
.B(n_2),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_242),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_265),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_253),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_230),
.B(n_304),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_247),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_289),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_290),
.B(n_2),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_304),
.B(n_3),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_248),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_295),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_302),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_249),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_258),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_308),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_255),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_233),
.B(n_4),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_261),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_263),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_266),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_267),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_268),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_270),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_325),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_254),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_327),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_274),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_335),
.B(n_285),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_337),
.B(n_278),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_341),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_280),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_310),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_284),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_350),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_355),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_365),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_288),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_362),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_348),
.B(n_296),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_297),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_344),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_324),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_428),
.B(n_254),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_428),
.B(n_433),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_352),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_396),
.B(n_428),
.Y(n_446)
);

OAI22xp33_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_323),
.B1(n_252),
.B2(n_257),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

INVx4_ASAP7_75t_SL g450 ( 
.A(n_385),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_353),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_395),
.A2(n_370),
.B1(n_357),
.B2(n_353),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_396),
.B(n_244),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_357),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_254),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

BUFx8_ASAP7_75t_SL g459 ( 
.A(n_413),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_404),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_425),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_370),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_414),
.B(n_373),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_428),
.B(n_254),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_396),
.B(n_259),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_384),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_395),
.A2(n_373),
.B1(n_322),
.B2(n_234),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_410),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_384),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_396),
.B(n_273),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_395),
.A2(n_434),
.B1(n_426),
.B2(n_420),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_420),
.B(n_277),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_279),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_393),
.B(n_298),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_393),
.B(n_281),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g489 ( 
.A(n_429),
.B(n_305),
.Y(n_489)
);

AND2x2_ASAP7_75t_SL g490 ( 
.A(n_434),
.B(n_311),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_435),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_436),
.B(n_416),
.C(n_421),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_389),
.B(n_283),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_388),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_429),
.B(n_399),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

OAI22x1_ASAP7_75t_L g504 ( 
.A1(n_437),
.A2(n_312),
.B1(n_319),
.B2(n_313),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_435),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_403),
.B(n_233),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_435),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_401),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_411),
.B(n_233),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_418),
.B(n_286),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_416),
.B(n_287),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_476),
.A2(n_434),
.B1(n_436),
.B2(n_437),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_446),
.B(n_431),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_449),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_431),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_465),
.B(n_438),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_424),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_430),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_419),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_444),
.B(n_432),
.Y(n_526)
);

AO22x2_ASAP7_75t_L g527 ( 
.A1(n_453),
.A2(n_439),
.B1(n_438),
.B2(n_432),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_461),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_464),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_493),
.A2(n_439),
.B1(n_430),
.B2(n_412),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_401),
.Y(n_533)
);

AO22x2_ASAP7_75t_L g534 ( 
.A1(n_455),
.A2(n_381),
.B1(n_387),
.B2(n_390),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_496),
.Y(n_536)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_511),
.Y(n_537)
);

BUFx8_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

OAI221xp5_ASAP7_75t_L g539 ( 
.A1(n_483),
.A2(n_390),
.B1(n_387),
.B2(n_391),
.C(n_406),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_391),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_467),
.A2(n_381),
.B1(n_6),
.B2(n_7),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_454),
.B(n_385),
.Y(n_543)
);

BUFx8_ASAP7_75t_L g544 ( 
.A(n_510),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_477),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_469),
.A2(n_381),
.B1(n_6),
.B2(n_7),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_475),
.B(n_427),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_479),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_505),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_443),
.A2(n_320),
.B1(n_317),
.B2(n_385),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_478),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_502),
.A2(n_385),
.B1(n_292),
.B2(n_316),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_473),
.B(n_385),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

BUFx8_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_463),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_460),
.B(n_385),
.Y(n_557)
);

OAI221xp5_ASAP7_75t_L g558 ( 
.A1(n_486),
.A2(n_398),
.B1(n_406),
.B2(n_405),
.C(n_400),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_463),
.B(n_413),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_482),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_442),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_422),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_490),
.A2(n_385),
.B1(n_315),
.B2(n_293),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_400),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_515),
.B(n_400),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_492),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_484),
.B(n_422),
.Y(n_568)
);

OAI221xp5_ASAP7_75t_L g569 ( 
.A1(n_486),
.A2(n_405),
.B1(n_398),
.B2(n_408),
.C(n_321),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_470),
.B(n_408),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_445),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_515),
.B(n_408),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_447),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_576)
);

AO22x2_ASAP7_75t_L g577 ( 
.A1(n_447),
.A2(n_441),
.B1(n_471),
.B2(n_512),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_509),
.B(n_299),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_441),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_488),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_471),
.A2(n_507),
.B1(n_512),
.B2(n_490),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_301),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_485),
.B(n_303),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_501),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_501),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_470),
.B(n_31),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_507),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_516),
.B(n_306),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_514),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_500),
.A2(n_314),
.B1(n_309),
.B2(n_276),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_504),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_489),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_489),
.B(n_19),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_498),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_459),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_499),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_554),
.B(n_500),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_522),
.B(n_480),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_533),
.B(n_500),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_526),
.B(n_466),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_524),
.B(n_513),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_548),
.B(n_499),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_568),
.B(n_583),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_530),
.B(n_450),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_518),
.B(n_472),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_550),
.B(n_458),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_562),
.B(n_458),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_SL g613 ( 
.A(n_559),
.B(n_458),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_582),
.B(n_458),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_547),
.B(n_462),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_595),
.B(n_462),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_590),
.B(n_462),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_SL g618 ( 
.A(n_521),
.B(n_462),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_519),
.B(n_472),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_523),
.B(n_528),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_531),
.B(n_481),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_535),
.B(n_481),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_536),
.B(n_497),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_542),
.B(n_497),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_525),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_529),
.B(n_451),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_578),
.B(n_545),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_564),
.B(n_451),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_SL g629 ( 
.A(n_551),
.B(n_456),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_532),
.B(n_456),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_532),
.B(n_457),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_592),
.B(n_233),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_520),
.B(n_233),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_552),
.B(n_276),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_596),
.B(n_276),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_560),
.B(n_276),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_567),
.B(n_19),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_570),
.B(n_32),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_540),
.B(n_276),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_572),
.B(n_276),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_571),
.B(n_20),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_543),
.B(n_21),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_593),
.B(n_36),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_597),
.B(n_37),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_577),
.B(n_21),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_601),
.B(n_38),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_598),
.B(n_39),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_566),
.B(n_40),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_577),
.B(n_22),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_575),
.B(n_42),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_553),
.B(n_45),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g652 ( 
.A(n_565),
.B(n_23),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_SL g653 ( 
.A(n_557),
.B(n_23),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_574),
.B(n_46),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_539),
.B(n_25),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_580),
.B(n_47),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_584),
.B(n_48),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_585),
.B(n_50),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_586),
.B(n_51),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_588),
.B(n_52),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_587),
.B(n_53),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_SL g662 ( 
.A(n_517),
.B(n_26),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_538),
.B(n_54),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_544),
.B(n_59),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_517),
.B(n_26),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_561),
.B(n_60),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_563),
.B(n_62),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_608),
.A2(n_581),
.B1(n_534),
.B2(n_527),
.Y(n_668)
);

AO31x2_ASAP7_75t_L g669 ( 
.A1(n_645),
.A2(n_573),
.A3(n_591),
.B(n_581),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_605),
.B(n_527),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_603),
.B(n_534),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_610),
.A2(n_558),
.B(n_569),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_638),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_638),
.B(n_541),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_619),
.A2(n_589),
.B(n_579),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_541),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_604),
.A2(n_589),
.B(n_579),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_627),
.A2(n_546),
.B1(n_576),
.B2(n_594),
.Y(n_678)
);

OA22x2_ASAP7_75t_L g679 ( 
.A1(n_649),
.A2(n_600),
.B1(n_576),
.B2(n_546),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_630),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_655),
.A2(n_594),
.B(n_556),
.C(n_549),
.Y(n_681)
);

OA22x2_ASAP7_75t_L g682 ( 
.A1(n_663),
.A2(n_556),
.B1(n_549),
.B2(n_537),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_623),
.A2(n_143),
.B(n_225),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_626),
.B(n_602),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_614),
.A2(n_142),
.B(n_223),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_632),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_641),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_628),
.A2(n_140),
.B(n_222),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_SL g690 ( 
.A(n_615),
.B(n_555),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_607),
.B(n_63),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_611),
.A2(n_139),
.B(n_218),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_620),
.B(n_64),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_634),
.A2(n_138),
.B(n_216),
.Y(n_694)
);

NAND3x1_ASAP7_75t_L g695 ( 
.A(n_631),
.B(n_27),
.C(n_28),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_617),
.A2(n_145),
.B(n_215),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_633),
.A2(n_137),
.B(n_214),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_625),
.Y(n_698)
);

O2A1O1Ixp5_ASAP7_75t_L g699 ( 
.A1(n_635),
.A2(n_135),
.B(n_213),
.C(n_67),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_613),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_612),
.A2(n_134),
.B1(n_211),
.B2(n_69),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_651),
.A2(n_148),
.B(n_210),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_609),
.A2(n_133),
.B1(n_209),
.B2(n_71),
.Y(n_703)
);

CKINVDCx11_ASAP7_75t_R g704 ( 
.A(n_664),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_616),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_662),
.B(n_74),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_643),
.A2(n_151),
.B(n_208),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_621),
.B(n_28),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_618),
.B(n_75),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_648),
.A2(n_154),
.B(n_76),
.Y(n_710)
);

AO31x2_ASAP7_75t_L g711 ( 
.A1(n_665),
.A2(n_30),
.A3(n_77),
.B(n_78),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_637),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_624),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_640),
.A2(n_639),
.B(n_650),
.Y(n_715)
);

AO22x2_ASAP7_75t_L g716 ( 
.A1(n_661),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_716)
);

INVx8_ASAP7_75t_L g717 ( 
.A(n_652),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_642),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_629),
.B(n_85),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_667),
.A2(n_88),
.B(n_90),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_712),
.B(n_636),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_671),
.A2(n_667),
.B(n_644),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_680),
.B(n_653),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_689),
.A2(n_683),
.B(n_715),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_702),
.A2(n_657),
.B(n_660),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_673),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_698),
.B(n_646),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_673),
.Y(n_728)
);

AO21x2_ASAP7_75t_L g729 ( 
.A1(n_677),
.A2(n_692),
.B(n_672),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_670),
.Y(n_730)
);

AOI21x1_ASAP7_75t_L g731 ( 
.A1(n_709),
.A2(n_659),
.B(n_658),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_717),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_714),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_681),
.A2(n_656),
.B(n_654),
.C(n_647),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_685),
.A2(n_666),
.B(n_92),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_704),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_705),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_674),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_738)
);

OA21x2_ASAP7_75t_L g739 ( 
.A1(n_675),
.A2(n_97),
.B(n_98),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_720),
.A2(n_104),
.B(n_105),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_688),
.B(n_107),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_674),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_742)
);

CKINVDCx14_ASAP7_75t_R g743 ( 
.A(n_690),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_686),
.B(n_113),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_713),
.B(n_114),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_688),
.B(n_115),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_694),
.A2(n_117),
.B(n_118),
.Y(n_747)
);

AOI21x1_ASAP7_75t_L g748 ( 
.A1(n_668),
.A2(n_120),
.B(n_121),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_679),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_669),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_SL g751 ( 
.A1(n_676),
.A2(n_128),
.B(n_130),
.C(n_157),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_719),
.A2(n_158),
.B(n_159),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_710),
.A2(n_162),
.B(n_163),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_717),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_713),
.B(n_164),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_696),
.A2(n_167),
.B(n_171),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_682),
.Y(n_757)
);

OAI21x1_ASAP7_75t_SL g758 ( 
.A1(n_707),
.A2(n_172),
.B(n_173),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_669),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_669),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_687),
.Y(n_761)
);

AOI222xp33_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_175),
.B1(n_177),
.B2(n_180),
.C1(n_181),
.C2(n_183),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_706),
.Y(n_763)
);

OAI21x1_ASAP7_75t_SL g764 ( 
.A1(n_684),
.A2(n_184),
.B(n_185),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_708),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_699),
.A2(n_186),
.B(n_187),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_706),
.A2(n_188),
.B1(n_190),
.B2(n_192),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_700),
.B(n_193),
.Y(n_768)
);

AO21x1_ASAP7_75t_L g769 ( 
.A1(n_691),
.A2(n_198),
.B(n_199),
.Y(n_769)
);

OAI21x1_ASAP7_75t_SL g770 ( 
.A1(n_700),
.A2(n_200),
.B(n_201),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_693),
.A2(n_202),
.B(n_203),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_761),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_750),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_726),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_760),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_765),
.B(n_678),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_759),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_761),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_739),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_729),
.A2(n_716),
.B(n_697),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_739),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_729),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_711),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_724),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_737),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_726),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_723),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_721),
.B(n_718),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_748),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_752),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_749),
.B(n_716),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_747),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_763),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_740),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_751),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_751),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_768),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_733),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_768),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_756),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_754),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_768),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_744),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_744),
.Y(n_804)
);

OA21x2_ASAP7_75t_L g805 ( 
.A1(n_722),
.A2(n_701),
.B(n_703),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_747),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_757),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_747),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_721),
.B(n_695),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_753),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_728),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_744),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_766),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_771),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_771),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_763),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_736),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_764),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_728),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_725),
.A2(n_711),
.B(n_206),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_735),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_758),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_731),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_745),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_769),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_787),
.B(n_746),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_817),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_824),
.B(n_754),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_R g829 ( 
.A(n_809),
.B(n_741),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_793),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_R g831 ( 
.A(n_774),
.B(n_743),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_807),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_787),
.B(n_749),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_R g834 ( 
.A(n_788),
.B(n_745),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_793),
.B(n_732),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_801),
.B(n_745),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_801),
.B(n_755),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_773),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_793),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_R g840 ( 
.A(n_774),
.B(n_743),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_824),
.B(n_755),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_786),
.B(n_755),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_773),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_793),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_793),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_816),
.B(n_727),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_776),
.B(n_742),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_798),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_816),
.B(n_762),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_816),
.B(n_711),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_785),
.B(n_742),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_R g852 ( 
.A(n_797),
.B(n_204),
.Y(n_852)
);

CKINVDCx11_ASAP7_75t_R g853 ( 
.A(n_816),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_R g854 ( 
.A(n_786),
.B(n_207),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_816),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_797),
.B(n_734),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_799),
.B(n_770),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_799),
.B(n_802),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_811),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_819),
.B(n_785),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_819),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_R g862 ( 
.A(n_802),
.B(n_220),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_772),
.B(n_767),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_772),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_R g865 ( 
.A(n_783),
.B(n_738),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_778),
.Y(n_866)
);

NAND2xp33_ASAP7_75t_R g867 ( 
.A(n_791),
.B(n_767),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_803),
.B(n_734),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_775),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_803),
.B(n_738),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_783),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_848),
.B(n_778),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_838),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_860),
.B(n_791),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_843),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_869),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_849),
.A2(n_812),
.B1(n_804),
.B2(n_818),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_871),
.B(n_775),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_863),
.B(n_782),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_845),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_864),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_858),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_858),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_866),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_826),
.B(n_812),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_868),
.Y(n_886)
);

AOI222xp33_ASAP7_75t_L g887 ( 
.A1(n_847),
.A2(n_795),
.B1(n_796),
.B2(n_818),
.C1(n_825),
.C2(n_804),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_868),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_827),
.B(n_822),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_856),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_870),
.B(n_782),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_870),
.B(n_782),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_850),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_861),
.B(n_777),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_844),
.B(n_784),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_851),
.B(n_808),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_857),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_857),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_865),
.B(n_777),
.Y(n_899)
);

AOI222xp33_ASAP7_75t_L g900 ( 
.A1(n_833),
.A2(n_796),
.B1(n_795),
.B2(n_825),
.C1(n_806),
.C2(n_808),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_832),
.B(n_823),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_859),
.Y(n_902)
);

AND2x4_ASAP7_75t_SL g903 ( 
.A(n_855),
.B(n_822),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_828),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_879),
.B(n_806),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_873),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_886),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_884),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_898),
.B(n_784),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_881),
.B(n_823),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_873),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_898),
.B(n_784),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_875),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_875),
.Y(n_914)
);

AND4x1_ASAP7_75t_L g915 ( 
.A(n_900),
.B(n_852),
.C(n_780),
.D(n_829),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_897),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_876),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_877),
.B(n_846),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_886),
.A2(n_805),
.B1(n_841),
.B2(n_862),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_884),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_888),
.A2(n_805),
.B1(n_828),
.B2(n_837),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_879),
.B(n_792),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_891),
.B(n_792),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_896),
.B(n_792),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_891),
.B(n_815),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_907),
.B(n_896),
.Y(n_926)
);

AND2x4_ASAP7_75t_SL g927 ( 
.A(n_925),
.B(n_899),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_916),
.B(n_893),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_906),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_916),
.B(n_893),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_918),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_909),
.B(n_912),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_911),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_911),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_924),
.B(n_874),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_905),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_892),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_913),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_913),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_932),
.Y(n_941)
);

INVxp33_ASAP7_75t_SL g942 ( 
.A(n_928),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_926),
.B(n_931),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_934),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_931),
.A2(n_867),
.B1(n_834),
.B2(n_915),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_933),
.B(n_914),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_928),
.B(n_840),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_SL g948 ( 
.A(n_930),
.B(n_831),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_941),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_944),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_946),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_948),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_938),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_945),
.B(n_915),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_942),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_947),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_954),
.A2(n_956),
.B(n_952),
.C(n_955),
.Y(n_957)
);

OAI221xp5_ASAP7_75t_L g958 ( 
.A1(n_956),
.A2(n_920),
.B1(n_908),
.B2(n_889),
.C(n_919),
.Y(n_958)
);

AOI322xp5_ASAP7_75t_L g959 ( 
.A1(n_954),
.A2(n_937),
.A3(n_930),
.B1(n_902),
.B2(n_938),
.C1(n_921),
.C2(n_899),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_953),
.B(n_927),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_949),
.B(n_880),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_960),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_957),
.B(n_950),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_958),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_962),
.Y(n_966)
);

INVxp33_ASAP7_75t_L g967 ( 
.A(n_964),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_963),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_965),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_962),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_966),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_959),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_967),
.B(n_951),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_970),
.Y(n_974)
);

NAND4xp75_ASAP7_75t_L g975 ( 
.A(n_969),
.B(n_853),
.C(n_897),
.D(n_878),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_SL g976 ( 
.A(n_968),
.B(n_854),
.C(n_842),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_967),
.B(n_900),
.C(n_901),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_968),
.Y(n_978)
);

OAI21x1_ASAP7_75t_SL g979 ( 
.A1(n_973),
.A2(n_971),
.B(n_972),
.Y(n_979)
);

OAI211xp5_ASAP7_75t_SL g980 ( 
.A1(n_978),
.A2(n_887),
.B(n_888),
.C(n_910),
.Y(n_980)
);

OAI211xp5_ASAP7_75t_SL g981 ( 
.A1(n_974),
.A2(n_936),
.B(n_885),
.C(n_890),
.Y(n_981)
);

AOI221xp5_ASAP7_75t_SL g982 ( 
.A1(n_975),
.A2(n_878),
.B1(n_940),
.B2(n_939),
.C(n_935),
.Y(n_982)
);

AOI221xp5_ASAP7_75t_L g983 ( 
.A1(n_977),
.A2(n_880),
.B1(n_927),
.B2(n_929),
.C(n_872),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_976),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_973),
.B(n_839),
.Y(n_985)
);

AOI222xp33_ASAP7_75t_L g986 ( 
.A1(n_972),
.A2(n_903),
.B1(n_836),
.B2(n_890),
.C1(n_794),
.C2(n_933),
.Y(n_986)
);

NAND4xp75_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_895),
.C(n_805),
.D(n_894),
.Y(n_987)
);

NOR2x1p5_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_883),
.Y(n_988)
);

XNOR2xp5_ASAP7_75t_L g989 ( 
.A(n_984),
.B(n_835),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_929),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_986),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_983),
.A2(n_835),
.B1(n_933),
.B2(n_903),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_980),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_981),
.B(n_895),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_991),
.B(n_830),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_914),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_989),
.B(n_882),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_992),
.B(n_912),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_993),
.B(n_882),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_990),
.B(n_917),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_987),
.B(n_994),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_SL g1002 ( 
.A(n_988),
.B(n_917),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_876),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_999),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_996),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_998),
.A2(n_912),
.B1(n_909),
.B2(n_883),
.Y(n_1007)
);

OAI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_1000),
.A2(n_805),
.B1(n_790),
.B2(n_794),
.C(n_789),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1002),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1001),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1009),
.Y(n_1011)
);

AND2x2_ASAP7_75t_SL g1012 ( 
.A(n_1006),
.B(n_909),
.Y(n_1012)
);

NOR4xp25_ASAP7_75t_SL g1013 ( 
.A(n_1010),
.B(n_790),
.C(n_815),
.D(n_779),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_1004),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_1005),
.B(n_1003),
.Y(n_1015)
);

AO22x2_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_1008),
.B1(n_1007),
.B2(n_904),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_820),
.B(n_894),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1013),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_1018),
.A2(n_925),
.B1(n_904),
.B2(n_810),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1017),
.A2(n_810),
.B1(n_924),
.B2(n_821),
.Y(n_1020)
);

OAI322xp33_ASAP7_75t_L g1021 ( 
.A1(n_1019),
.A2(n_1015),
.A3(n_1016),
.B1(n_789),
.B2(n_821),
.C1(n_813),
.C2(n_800),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_1020),
.A2(n_789),
.B(n_814),
.C(n_800),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1021),
.A2(n_814),
.B(n_810),
.C(n_813),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_1022),
.A2(n_820),
.B(n_810),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1024),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_1025),
.A2(n_779),
.B1(n_781),
.B2(n_784),
.C(n_922),
.Y(n_1027)
);

AOI211xp5_ASAP7_75t_L g1028 ( 
.A1(n_1027),
.A2(n_1026),
.B(n_922),
.C(n_923),
.Y(n_1028)
);


endmodule