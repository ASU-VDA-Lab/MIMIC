module fake_ibex_74_n_1166 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_132, n_174, n_210, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1166);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_132;
input n_174;
input n_210;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1166;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1148;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1134;
wire n_727;
wire n_1138;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_698;
wire n_498;
wire n_375;
wire n_280;
wire n_317;
wire n_340;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1140;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_711;
wire n_497;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_732;
wire n_673;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_1057;
wire n_325;
wire n_301;
wire n_617;
wire n_496;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_1075;
wire n_1136;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_1020;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_1070;
wire n_454;
wire n_980;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1028;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_234;
wire n_300;
wire n_1151;
wire n_1135;
wire n_1146;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1062;
wire n_847;
wire n_830;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_630;
wire n_354;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_1158;
wire n_745;
wire n_329;
wire n_1149;
wire n_447;
wire n_940;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_1160;
wire n_615;
wire n_512;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1118;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_899;
wire n_843;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_700;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_741;
wire n_430;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_977;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_1150;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_921;
wire n_890;
wire n_912;
wire n_1058;
wire n_1105;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_1000;
wire n_394;
wire n_984;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_67),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_62),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_28),
.B(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_68),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_76),
.B(n_153),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_96),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_31),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_102),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_14),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_18),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_97),
.Y(n_230)
);

BUFx2_ASAP7_75t_SL g231 ( 
.A(n_186),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_112),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_61),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_20),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx12_ASAP7_75t_R g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_125),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_55),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_74),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_182),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_7),
.B(n_108),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_91),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_94),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_99),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_18),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_60),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_106),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_163),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_117),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_124),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_159),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_32),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_41),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_84),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_146),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_134),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_72),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_23),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_36),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_42),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_82),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_196),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_107),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_121),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_203),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_160),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_187),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_87),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_122),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_56),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_147),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_195),
.B(n_138),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_133),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_120),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_79),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_63),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_30),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_183),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_179),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_9),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_101),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_119),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_129),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_175),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_152),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_197),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_144),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_3),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_29),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_151),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_154),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_198),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_11),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_25),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_189),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_110),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_169),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_21),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_199),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_53),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_54),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_149),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_83),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_31),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_77),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_173),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_43),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_8),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_69),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_130),
.B(n_0),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_57),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_135),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_51),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_98),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_24),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_70),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_34),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_65),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_85),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_168),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_166),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_78),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_100),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_126),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_44),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_22),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_208),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_127),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_41),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_118),
.B(n_164),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_140),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_205),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_17),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_58),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_150),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_177),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_229),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_279),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_229),
.B(n_1),
.Y(n_376)
);

OAI22x1_ASAP7_75t_R g377 ( 
.A1(n_241),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_299),
.B(n_4),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_233),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g380 ( 
.A1(n_255),
.A2(n_89),
.B(n_211),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_5),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_233),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_227),
.Y(n_383)
);

BUFx8_ASAP7_75t_SL g384 ( 
.A(n_241),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_240),
.B(n_6),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_250),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_299),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_294),
.B(n_228),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_287),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_233),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_237),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_327),
.B(n_6),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_294),
.B(n_7),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_304),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_8),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_240),
.B(n_9),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_237),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_236),
.B(n_10),
.Y(n_401)
);

INVxp33_ASAP7_75t_SL g402 ( 
.A(n_287),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_270),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_240),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_310),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_310),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_257),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_237),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_307),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_261),
.B(n_12),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_281),
.B(n_13),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_281),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_263),
.B(n_13),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_281),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_237),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_250),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_266),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_293),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_310),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_293),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_275),
.B(n_15),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_293),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_282),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_331),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_310),
.Y(n_427)
);

OAI22x1_ASAP7_75t_R g428 ( 
.A1(n_270),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_293),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_215),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_338),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_255),
.Y(n_433)
);

BUFx12f_ASAP7_75t_L g434 ( 
.A(n_243),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_265),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_267),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

BUFx8_ASAP7_75t_L g438 ( 
.A(n_213),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_273),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_273),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_265),
.A2(n_104),
.B(n_210),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_297),
.B(n_283),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_283),
.B(n_64),
.Y(n_443)
);

BUFx8_ASAP7_75t_SL g444 ( 
.A(n_311),
.Y(n_444)
);

AOI22x1_ASAP7_75t_SL g445 ( 
.A1(n_311),
.A2(n_215),
.B1(n_223),
.B2(n_216),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_300),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_216),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_306),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_297),
.B(n_32),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_223),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_306),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_235),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_218),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_316),
.B(n_351),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_286),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_316),
.B(n_37),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_224),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_351),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_230),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_286),
.B(n_40),
.Y(n_464)
);

AO22x1_ASAP7_75t_L g465 ( 
.A1(n_284),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_326),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_296),
.B(n_46),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_234),
.B(n_48),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_231),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_285),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_246),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_296),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_247),
.B(n_48),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_323),
.B(n_49),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_323),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g476 ( 
.A(n_308),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_235),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_320),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_248),
.B(n_249),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_251),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_339),
.Y(n_481)
);

CKINVDCx6p67_ASAP7_75t_R g482 ( 
.A(n_238),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_439),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

AO22x2_ASAP7_75t_L g486 ( 
.A1(n_430),
.A2(n_225),
.B1(n_305),
.B2(n_371),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_391),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_442),
.B(n_212),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_383),
.B(n_226),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_404),
.B(n_318),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_482),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_252),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g499 ( 
.A1(n_460),
.A2(n_256),
.B(n_253),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_398),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_415),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_376),
.Y(n_504)
);

OA22x2_ASAP7_75t_L g505 ( 
.A1(n_375),
.A2(n_321),
.B1(n_328),
.B2(n_332),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_376),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_459),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_413),
.B(n_365),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_378),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_426),
.A2(n_383),
.B1(n_402),
.B2(n_430),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_443),
.B(n_220),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_472),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_415),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_406),
.B(n_335),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_379),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_464),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_467),
.B(n_259),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_403),
.B(n_217),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_387),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g528 ( 
.A1(n_460),
.A2(n_262),
.B(n_260),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_424),
.B(n_344),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_389),
.Y(n_531)
);

AND3x2_ASAP7_75t_L g532 ( 
.A(n_424),
.B(n_245),
.C(n_264),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_443),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_481),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_390),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_451),
.B(n_239),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_449),
.B(n_345),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_467),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_415),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_481),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_386),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_402),
.A2(n_319),
.B1(n_244),
.B2(n_368),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_457),
.B(n_268),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_379),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_461),
.B(n_269),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_374),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_382),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_382),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_392),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_386),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_392),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_436),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_397),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_480),
.B(n_474),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_469),
.B(n_369),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_410),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_448),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_448),
.B(n_369),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_443),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_385),
.B(n_302),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_478),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_478),
.B(n_373),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_417),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_393),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_393),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_405),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_381),
.A2(n_239),
.B1(n_368),
.B2(n_244),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_435),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_434),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_405),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

CKINVDCx6p67_ASAP7_75t_R g575 ( 
.A(n_476),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_348),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_450),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_388),
.B(n_350),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_407),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_458),
.B(n_274),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_458),
.B(n_276),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_407),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_407),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_479),
.B(n_277),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_431),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_388),
.B(n_353),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_420),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_462),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_479),
.B(n_280),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_399),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_380),
.A2(n_289),
.B(n_288),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_432),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_420),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_463),
.B(n_471),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_412),
.B(n_363),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_408),
.B(n_295),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_384),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_418),
.B(n_214),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_420),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_425),
.B(n_221),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_427),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_427),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_468),
.B(n_303),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_475),
.B(n_301),
.Y(n_606)
);

AOI21x1_ASAP7_75t_L g607 ( 
.A1(n_441),
.A2(n_313),
.B(n_309),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_314),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_427),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_429),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_447),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_475),
.B(n_317),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_429),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_455),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_429),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_421),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_475),
.B(n_222),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_475),
.B(n_325),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_473),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_411),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_423),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_394),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_411),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_422),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_400),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_422),
.Y(n_629)
);

CKINVDCx6p67_ASAP7_75t_R g630 ( 
.A(n_401),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_444),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_542),
.B(n_381),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_477),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_618),
.B(n_622),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_541),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_623),
.B(n_333),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_626),
.B(n_340),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_627),
.B(n_438),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_438),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_585),
.B(n_346),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_578),
.B(n_347),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_502),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_587),
.B(n_352),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_355),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_560),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_590),
.B(n_358),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_591),
.B(n_466),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_503),
.B(n_219),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_502),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_563),
.B(n_449),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_488),
.B(n_452),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_490),
.B(n_232),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_557),
.B(n_242),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_515),
.B(n_465),
.C(n_364),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

O2A1O1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_513),
.A2(n_454),
.B(n_452),
.C(n_319),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_564),
.Y(n_661)
);

OAI21xp33_ASAP7_75t_L g662 ( 
.A1(n_516),
.A2(n_312),
.B(n_254),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_602),
.B(n_258),
.Y(n_663)
);

INVxp33_ASAP7_75t_L g664 ( 
.A(n_520),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_566),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_551),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_519),
.B(n_372),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_515),
.B(n_454),
.C(n_367),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_630),
.B(n_303),
.Y(n_670)
);

BUFx5_ASAP7_75t_L g671 ( 
.A(n_597),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_543),
.Y(n_672)
);

BUFx5_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_612),
.B(n_271),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_554),
.Y(n_675)
);

BUFx6f_ASAP7_75t_SL g676 ( 
.A(n_555),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_615),
.B(n_278),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_617),
.B(n_290),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_538),
.B(n_291),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_538),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_292),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_565),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_574),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_577),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_504),
.B(n_298),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_521),
.B(n_360),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_533),
.B(n_315),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_507),
.A2(n_360),
.B1(n_409),
.B2(n_416),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_556),
.B(n_493),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_510),
.A2(n_419),
.B1(n_322),
.B2(n_356),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_529),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_539),
.B(n_576),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_586),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_556),
.B(n_324),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_527),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_511),
.B(n_329),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_531),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_562),
.A2(n_349),
.B1(n_336),
.B2(n_337),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_330),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_566),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_535),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_565),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_605),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_553),
.B(n_343),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_484),
.B(n_354),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_485),
.B(n_359),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_594),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_571),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_500),
.B(n_377),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_489),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_489),
.Y(n_713)
);

AO221x1_ASAP7_75t_L g714 ( 
.A1(n_486),
.A2(n_445),
.B1(n_428),
.B2(n_444),
.C(n_53),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_597),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_66),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_555),
.B(n_50),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_495),
.B(n_51),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_589),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_589),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_597),
.B(n_137),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_555),
.B(n_52),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_562),
.B(n_52),
.C(n_54),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_494),
.B(n_525),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_558),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_605),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_572),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_584),
.B(n_88),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_584),
.B(n_90),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_509),
.B(n_92),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_608),
.B(n_93),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_537),
.A2(n_105),
.B1(n_111),
.B2(n_115),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_532),
.Y(n_735)
);

AND2x6_ASAP7_75t_SL g736 ( 
.A(n_537),
.B(n_123),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_570),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_483),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_483),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_487),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_599),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_575),
.B(n_128),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_634),
.A2(n_581),
.B(n_580),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_632),
.B(n_580),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_632),
.A2(n_581),
.B(n_613),
.Y(n_745)
);

CKINVDCx10_ASAP7_75t_R g746 ( 
.A(n_676),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_679),
.A2(n_621),
.B(n_606),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_657),
.A2(n_598),
.B(n_544),
.C(n_546),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_660),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_635),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_677),
.A2(n_546),
.B(n_620),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_677),
.A2(n_596),
.B(n_540),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_664),
.B(n_536),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_669),
.B(n_537),
.Y(n_754)
);

BUFx2_ASAP7_75t_SL g755 ( 
.A(n_676),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_678),
.A2(n_596),
.B(n_540),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_659),
.A2(n_690),
.B(n_711),
.C(n_704),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_681),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_731),
.A2(n_592),
.B(n_607),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_712),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_636),
.B(n_486),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_637),
.A2(n_526),
.B(n_631),
.C(n_624),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_643),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_637),
.A2(n_526),
.B(n_624),
.C(n_619),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_712),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_696),
.B(n_698),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_702),
.B(n_499),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_668),
.A2(n_505),
.B1(n_526),
.B2(n_528),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_645),
.B(n_505),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_651),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_687),
.B(n_619),
.Y(n_773)
);

NAND2x1_ASAP7_75t_L g774 ( 
.A(n_713),
.B(n_658),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_686),
.A2(n_517),
.B(n_534),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_638),
.B(n_492),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_686),
.A2(n_518),
.B(n_534),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_647),
.A2(n_644),
.B(n_642),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_642),
.A2(n_517),
.B(n_530),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_737),
.A2(n_625),
.B(n_514),
.C(n_530),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_657),
.A2(n_512),
.B(n_508),
.C(n_506),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

CKINVDCx10_ASAP7_75t_R g783 ( 
.A(n_741),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_640),
.B(n_496),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_496),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_649),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_729),
.Y(n_787)
);

OAI21xp33_ASAP7_75t_L g788 ( 
.A1(n_654),
.A2(n_625),
.B(n_497),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_684),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_646),
.A2(n_501),
.B(n_498),
.C(n_628),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_706),
.A2(n_498),
.B(n_573),
.Y(n_791)
);

AO21x1_ASAP7_75t_L g792 ( 
.A1(n_716),
.A2(n_610),
.B(n_614),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_727),
.B(n_136),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_639),
.B(n_141),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_661),
.A2(n_628),
.B(n_614),
.C(n_611),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_685),
.B(n_628),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_668),
.A2(n_733),
.B(n_730),
.C(n_725),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_694),
.B(n_142),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_707),
.B(n_143),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_652),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_633),
.B(n_726),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_726),
.B(n_145),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_699),
.B(n_148),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_693),
.A2(n_548),
.B(n_609),
.C(n_604),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_689),
.A2(n_549),
.B1(n_604),
.B2(n_603),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_666),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_674),
.A2(n_545),
.B(n_550),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_720),
.A2(n_545),
.B(n_603),
.C(n_601),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_705),
.B(n_156),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_641),
.B(n_616),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_683),
.Y(n_812)
);

AND2x2_ASAP7_75t_SL g813 ( 
.A(n_670),
.B(n_158),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_653),
.B(n_162),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_710),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_648),
.A2(n_552),
.B1(n_601),
.B2(n_595),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_663),
.B(n_165),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_703),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_719),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_722),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_718),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_648),
.B(n_170),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_700),
.A2(n_656),
.B(n_697),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_721),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_655),
.A2(n_567),
.B(n_568),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_735),
.A2(n_567),
.B(n_595),
.C(n_593),
.Y(n_826)
);

NOR2x2_ASAP7_75t_L g827 ( 
.A(n_672),
.B(n_171),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_665),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_682),
.A2(n_568),
.B(n_569),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_742),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_723),
.A2(n_588),
.B(n_583),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_714),
.A2(n_579),
.B1(n_583),
.B2(n_582),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_708),
.A2(n_695),
.B(n_688),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_701),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_732),
.A2(n_180),
.B(n_181),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_789),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_792),
.A2(n_740),
.A3(n_739),
.B(n_738),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_787),
.B(n_662),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_754),
.B(n_717),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_813),
.B(n_724),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_761),
.B(n_734),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_782),
.Y(n_842)
);

OA22x2_ASAP7_75t_L g843 ( 
.A1(n_755),
.A2(n_822),
.B1(n_770),
.B2(n_771),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_778),
.B(n_715),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_753),
.B(n_650),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_801),
.B(n_667),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_823),
.A2(n_691),
.B(n_728),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_778),
.B(n_736),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_744),
.B(n_715),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_769),
.A2(n_751),
.B(n_768),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_783),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_773),
.B(n_715),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_745),
.A2(n_748),
.B(n_743),
.Y(n_853)
);

AO31x2_ASAP7_75t_L g854 ( 
.A1(n_831),
.A2(n_715),
.A3(n_673),
.B(n_671),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_757),
.B(n_830),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_762),
.A2(n_673),
.B(n_671),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_749),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_761),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_761),
.B(n_201),
.Y(n_859)
);

AOI21xp33_ASAP7_75t_L g860 ( 
.A1(n_780),
.A2(n_616),
.B(n_522),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_814),
.A2(n_817),
.B(n_794),
.C(n_809),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_766),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_766),
.B(n_767),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_747),
.A2(n_752),
.B(n_756),
.Y(n_864)
);

AO31x2_ASAP7_75t_L g865 ( 
.A1(n_835),
.A2(n_808),
.A3(n_804),
.B(n_781),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_763),
.A2(n_790),
.B(n_795),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_767),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_827),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_776),
.A2(n_802),
.B(n_788),
.C(n_833),
.Y(n_869)
);

AOI211x1_ASAP7_75t_L g870 ( 
.A1(n_784),
.A2(n_785),
.B(n_803),
.C(n_779),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_815),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_816),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_758),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_759),
.B(n_764),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_746),
.B(n_800),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_828),
.B(n_834),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_772),
.B(n_821),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_750),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_824),
.B(n_819),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_796),
.Y(n_880)
);

OAI22x1_ASAP7_75t_L g881 ( 
.A1(n_783),
.A2(n_746),
.B1(n_832),
.B2(n_811),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_793),
.B(n_774),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_825),
.A2(n_775),
.B(n_777),
.Y(n_883)
);

AOI21xp33_ASAP7_75t_L g884 ( 
.A1(n_826),
.A2(n_799),
.B(n_798),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_820),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_832),
.A2(n_805),
.B(n_786),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_829),
.A2(n_791),
.B(n_807),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_806),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_806),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_L g890 ( 
.A1(n_810),
.A2(n_792),
.B(n_831),
.C(n_797),
.Y(n_890)
);

INVx8_ASAP7_75t_L g891 ( 
.A(n_812),
.Y(n_891)
);

BUFx5_ASAP7_75t_L g892 ( 
.A(n_818),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_778),
.A2(n_823),
.B(n_765),
.C(n_743),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_761),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_782),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_761),
.B(n_766),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_797),
.A2(n_760),
.B(n_792),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_789),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_787),
.B(n_653),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_778),
.B(n_634),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_761),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_778),
.B(n_634),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_787),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_778),
.B(n_634),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_782),
.Y(n_905)
);

BUFx12f_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_797),
.A2(n_745),
.B(n_748),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_787),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_761),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_634),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_760),
.A2(n_515),
.B(n_561),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_797),
.A2(n_760),
.B(n_792),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_778),
.B(n_634),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_761),
.B(n_727),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_782),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_787),
.B(n_692),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_778),
.B(n_634),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_782),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_778),
.B(n_634),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_797),
.A2(n_745),
.B(n_748),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_778),
.B(n_634),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_787),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_692),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_782),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_761),
.B(n_727),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_778),
.B(n_634),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_797),
.A2(n_745),
.B(n_748),
.Y(n_928)
);

OAI22x1_ASAP7_75t_L g929 ( 
.A1(n_787),
.A2(n_543),
.B1(n_570),
.B2(n_477),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_787),
.B(n_692),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_778),
.B(n_634),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_903),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_872),
.Y(n_934)
);

CKINVDCx16_ASAP7_75t_R g935 ( 
.A(n_868),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_899),
.B(n_840),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_908),
.B(n_923),
.Y(n_937)
);

BUFx4f_ASAP7_75t_SL g938 ( 
.A(n_894),
.Y(n_938)
);

INVx6_ASAP7_75t_L g939 ( 
.A(n_909),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_916),
.B(n_924),
.Y(n_940)
);

AO21x2_ASAP7_75t_L g941 ( 
.A1(n_907),
.A2(n_928),
.B(n_921),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_909),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_861),
.A2(n_893),
.B(n_884),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_884),
.A2(n_847),
.B(n_850),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_902),
.A2(n_927),
.B(n_904),
.C(n_931),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_929),
.A2(n_855),
.B1(n_846),
.B2(n_845),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_930),
.Y(n_947)
);

BUFx2_ASAP7_75t_SL g948 ( 
.A(n_909),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_842),
.Y(n_949)
);

CKINVDCx6p67_ASAP7_75t_R g950 ( 
.A(n_901),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_898),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_883),
.A2(n_887),
.B(n_869),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_875),
.B(n_881),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_839),
.A2(n_838),
.B1(n_880),
.B2(n_841),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_866),
.A2(n_853),
.B(n_844),
.Y(n_955)
);

OAI21x1_ASAP7_75t_SL g956 ( 
.A1(n_900),
.A2(n_913),
.B(n_920),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_895),
.B(n_905),
.Y(n_957)
);

OAI21x1_ASAP7_75t_SL g958 ( 
.A1(n_910),
.A2(n_922),
.B(n_917),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_857),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_915),
.B(n_918),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_925),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_874),
.B(n_877),
.Y(n_962)
);

OA21x2_ASAP7_75t_L g963 ( 
.A1(n_890),
.A2(n_864),
.B(n_853),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_871),
.B(n_873),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_879),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_863),
.B(n_843),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_885),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_866),
.A2(n_886),
.B1(n_852),
.B2(n_878),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_862),
.B(n_867),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_851),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_886),
.B(n_870),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_876),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_891),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_891),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_862),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_876),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_896),
.B(n_867),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_860),
.A2(n_912),
.B(n_897),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_858),
.B(n_870),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_914),
.B(n_926),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_912),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_859),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_849),
.B(n_889),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_860),
.A2(n_856),
.B(n_911),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_888),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_892),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_854),
.A2(n_837),
.B(n_892),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_854),
.A2(n_837),
.B(n_865),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_882),
.A2(n_888),
.B1(n_889),
.B2(n_865),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_882),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_899),
.B(n_737),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_899),
.B(n_634),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_903),
.Y(n_993)
);

OR3x4_ASAP7_75t_SL g994 ( 
.A(n_868),
.B(n_737),
.C(n_746),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_848),
.A2(n_657),
.B(n_668),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_906),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_899),
.B(n_634),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_836),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_940),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_962),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_962),
.B(n_941),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_979),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_941),
.B(n_949),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_985),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_956),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_958),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_991),
.A2(n_936),
.B1(n_954),
.B2(n_946),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_949),
.B(n_959),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_959),
.Y(n_1009)
);

BUFx2_ASAP7_75t_SL g1010 ( 
.A(n_932),
.Y(n_1010)
);

OR2x2_ASAP7_75t_SL g1011 ( 
.A(n_935),
.B(n_939),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_992),
.B(n_997),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_965),
.B(n_947),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_985),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_SL g1015 ( 
.A1(n_953),
.A2(n_948),
.B1(n_933),
.B2(n_993),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_937),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_938),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_998),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_932),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_932),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_932),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_934),
.Y(n_1022)
);

AO21x1_ASAP7_75t_SL g1023 ( 
.A1(n_989),
.A2(n_983),
.B(n_968),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_964),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_967),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_939),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_957),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_SL g1028 ( 
.A1(n_953),
.A2(n_936),
.B1(n_982),
.B2(n_969),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_960),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_961),
.B(n_951),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_986),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_986),
.B(n_975),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_939),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_944),
.A2(n_952),
.B(n_943),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_942),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_942),
.Y(n_1036)
);

OAI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_953),
.A2(n_982),
.B1(n_975),
.B2(n_938),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_996),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_963),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_963),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_963),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_SL g1042 ( 
.A(n_970),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1003),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_1007),
.A2(n_966),
.B(n_995),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1031),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1001),
.B(n_981),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1022),
.Y(n_1047)
);

OA211x2_ASAP7_75t_L g1048 ( 
.A1(n_1011),
.A2(n_999),
.B(n_1010),
.C(n_969),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1001),
.B(n_1002),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1027),
.B(n_945),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1005),
.B(n_987),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1008),
.B(n_978),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1009),
.B(n_978),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1009),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1028),
.A2(n_966),
.B1(n_961),
.B2(n_955),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1034),
.B(n_988),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1000),
.A2(n_972),
.B1(n_976),
.B2(n_971),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1023),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1018),
.B(n_945),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1016),
.B(n_990),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1025),
.B(n_984),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1044),
.B(n_1038),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1047),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1044),
.A2(n_1037),
.B1(n_1014),
.B2(n_1015),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_1058),
.A2(n_1011),
.B1(n_1014),
.B2(n_1019),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1060),
.B(n_1042),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_1047),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_1049),
.B(n_1034),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1049),
.B(n_1034),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1054),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_1045),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1045),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1060),
.B(n_1004),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1049),
.B(n_1039),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1046),
.B(n_1052),
.Y(n_1075)
);

OAI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_1055),
.A2(n_1012),
.B1(n_1010),
.B2(n_1029),
.C(n_1027),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1046),
.B(n_1039),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1050),
.B(n_1029),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1046),
.B(n_1040),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1052),
.B(n_1040),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1050),
.B(n_1024),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1061),
.B(n_1041),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_1056),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1072),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1070),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1075),
.B(n_1056),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1063),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1075),
.B(n_1056),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1080),
.B(n_1051),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1069),
.B(n_1053),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1066),
.B(n_1019),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1069),
.B(n_1059),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1071),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1076),
.A2(n_1055),
.B1(n_1048),
.B2(n_1058),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1070),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1068),
.B(n_1043),
.Y(n_1096)
);

AND2x4_ASAP7_75t_SL g1097 ( 
.A(n_1063),
.B(n_1045),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1086),
.B(n_1077),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_1096),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1092),
.B(n_1062),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_1097),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1085),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1085),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1086),
.B(n_1079),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_1090),
.B(n_1098),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1088),
.B(n_1098),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1095),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1089),
.B(n_1082),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1088),
.B(n_1079),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1104),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1103),
.Y(n_1112)
);

XOR2x2_ASAP7_75t_L g1113 ( 
.A(n_1106),
.B(n_1065),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1106),
.B(n_1090),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1107),
.B(n_1083),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1104),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1108),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1100),
.B(n_1092),
.Y(n_1118)
);

AOI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1101),
.A2(n_1076),
.B(n_1064),
.Y(n_1119)
);

OAI32xp33_ASAP7_75t_L g1120 ( 
.A1(n_1102),
.A2(n_1094),
.A3(n_1064),
.B1(n_1087),
.B2(n_1067),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1107),
.B(n_1083),
.Y(n_1121)
);

OAI32xp33_ASAP7_75t_L g1122 ( 
.A1(n_1102),
.A2(n_1087),
.A3(n_1067),
.B1(n_1093),
.B2(n_1084),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1099),
.B(n_1096),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1123),
.B(n_1099),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1113),
.A2(n_1109),
.B1(n_1065),
.B2(n_1089),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1113),
.A2(n_1109),
.B1(n_1089),
.B2(n_1073),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1111),
.Y(n_1128)
);

OAI32xp33_ASAP7_75t_L g1129 ( 
.A1(n_1114),
.A2(n_1110),
.A3(n_1105),
.B1(n_1091),
.B2(n_1021),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_1120),
.B1(n_1119),
.B2(n_1122),
.C(n_1118),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1124),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_L g1132 ( 
.A(n_1126),
.B(n_1115),
.Y(n_1132)
);

OAI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_1127),
.A2(n_1121),
.B(n_1115),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1125),
.A2(n_1121),
.B1(n_1109),
.B2(n_1105),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1128),
.B(n_1117),
.C(n_1116),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1124),
.B(n_1110),
.Y(n_1136)
);

OAI211xp5_ASAP7_75t_L g1137 ( 
.A1(n_1130),
.A2(n_1020),
.B(n_994),
.C(n_1017),
.Y(n_1137)
);

NOR3xp33_ASAP7_75t_L g1138 ( 
.A(n_1132),
.B(n_1020),
.C(n_994),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_1135),
.B(n_1131),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1134),
.B(n_1109),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1136),
.Y(n_1141)
);

NAND4xp25_ASAP7_75t_L g1142 ( 
.A(n_1133),
.B(n_1048),
.C(n_1017),
.D(n_1057),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1141),
.B(n_1112),
.Y(n_1143)
);

NAND5xp2_ASAP7_75t_L g1144 ( 
.A(n_1137),
.B(n_1057),
.C(n_1032),
.D(n_1006),
.E(n_1024),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1140),
.B(n_1093),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1142),
.A2(n_1112),
.B(n_1013),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1017),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_1108),
.Y(n_1149)
);

NOR2x1_ASAP7_75t_SL g1150 ( 
.A(n_1143),
.B(n_974),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_1144),
.B(n_974),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1147),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1152),
.Y(n_1153)
);

NAND4xp75_ASAP7_75t_L g1154 ( 
.A(n_1151),
.B(n_1026),
.C(n_1033),
.D(n_980),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1154),
.A2(n_1148),
.B1(n_1149),
.B2(n_1150),
.Y(n_1155)
);

XNOR2x1_ASAP7_75t_L g1156 ( 
.A(n_1153),
.B(n_1149),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1156),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_1078),
.B1(n_1081),
.B2(n_1093),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1157),
.A2(n_950),
.B1(n_1036),
.B2(n_1035),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1159),
.A2(n_1158),
.B1(n_1026),
.B2(n_1033),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1159),
.Y(n_1161)
);

OA22x2_ASAP7_75t_L g1162 ( 
.A1(n_1161),
.A2(n_1097),
.B1(n_1025),
.B2(n_977),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1162),
.B(n_1160),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1163),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_1164),
.B(n_973),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_1030),
.B(n_973),
.Y(n_1166)
);


endmodule