module fake_jpeg_23604_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_45),
.C(n_30),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_1),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_51),
.B1(n_59),
.B2(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_74),
.B1(n_16),
.B2(n_3),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_30),
.B2(n_21),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_64),
.B1(n_55),
.B2(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_42),
.B1(n_24),
.B2(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_20),
.B1(n_29),
.B2(n_22),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_22),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_16),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_83),
.B1(n_50),
.B2(n_67),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_91),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_47),
.B1(n_73),
.B2(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_2),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_35),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_48),
.B(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_16),
.C(n_4),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_95),
.C(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_4),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_8),
.Y(n_109)
);

NAND2x1_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_6),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_6),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_7),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_57),
.B(n_8),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_9),
.Y(n_121)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_120),
.B1(n_95),
.B2(n_80),
.Y(n_141)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_118),
.B1(n_96),
.B2(n_95),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_47),
.B1(n_72),
.B2(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_89),
.A2(n_77),
.B1(n_82),
.B2(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_84),
.Y(n_126)
);

NOR4xp25_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_85),
.C(n_92),
.D(n_78),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_138),
.B1(n_110),
.B2(n_103),
.C(n_112),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_131),
.B1(n_141),
.B2(n_118),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_82),
.B1(n_87),
.B2(n_100),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_111),
.C(n_105),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_110),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_100),
.B(n_80),
.Y(n_138)
);

BUFx12f_ASAP7_75t_SL g139 ( 
.A(n_122),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_109),
.C(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_114),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_114),
.B(n_116),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_144),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_148),
.C(n_155),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_111),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_150),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_165),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_152),
.B(n_14),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_129),
.B1(n_127),
.B2(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_143),
.B1(n_142),
.B2(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_135),
.C(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_161),
.C(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_170),
.C(n_172),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_123),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_123),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_157),
.C(n_166),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_11),
.B(n_159),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_178),
.Y(n_184)
);

AOI31xp33_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_125),
.A3(n_167),
.B(n_171),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_165),
.B1(n_158),
.B2(n_156),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_132),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_174),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_169),
.A2(n_125),
.B(n_136),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_181),
.A2(n_168),
.B(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_180),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_179),
.C(n_176),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_184),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule