module fake_jpeg_3107_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx12f_ASAP7_75t_SL g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_0),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_76),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_55),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_98),
.B1(n_52),
.B2(n_68),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_76),
.B1(n_56),
.B2(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_114),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_65),
.B1(n_64),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_116),
.B1(n_70),
.B2(n_60),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_67),
.C(n_60),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_100),
.C(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_66),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_68),
.B1(n_71),
.B2(n_58),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_90),
.B1(n_56),
.B2(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_126),
.B1(n_12),
.B2(n_14),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_108),
.B1(n_9),
.B2(n_10),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_70),
.B1(n_72),
.B2(n_68),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_3),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_4),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_58),
.C(n_33),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_12),
.C(n_14),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_7),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_5),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_34),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_149),
.C(n_161),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_8),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_145),
.B(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_50),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_16),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_37),
.B1(n_47),
.B2(n_46),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_15),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_181),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_135),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_184),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_138),
.B(n_20),
.Y(n_182)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_182),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_153),
.B1(n_163),
.B2(n_168),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_159),
.B(n_151),
.C(n_156),
.D(n_152),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_183),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_147),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_170),
.Y(n_194)
);

OA21x2_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_146),
.B(n_161),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.C(n_27),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_184),
.C(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_200),
.B1(n_175),
.B2(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_169),
.C(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_190),
.B1(n_176),
.B2(n_178),
.Y(n_203)
);

FAx1_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_192),
.CI(n_170),
.CON(n_204),
.SN(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_197),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_201),
.B(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_205),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_204),
.C(n_35),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_209),
.B(n_29),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_39),
.Y(n_211)
);

OAI311xp33_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_41),
.A3(n_42),
.B1(n_43),
.C1(n_44),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_45),
.Y(n_213)
);


endmodule