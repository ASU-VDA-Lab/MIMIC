module fake_jpeg_29259_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_4),
.B(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_18),
.B1(n_9),
.B2(n_10),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_28),
.B1(n_16),
.B2(n_6),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_14),
.C(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_24),
.B1(n_9),
.B2(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_6),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_30),
.B1(n_29),
.B2(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B(n_33),
.Y(n_36)
);

AOI321xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_10),
.A3(n_13),
.B1(n_35),
.B2(n_29),
.C(n_30),
.Y(n_37)
);


endmodule