module fake_ariane_938_n_1705 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1705);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1705;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_64),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_18),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_5),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_84),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_52),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_22),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_19),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_5),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_19),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_57),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_9),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_62),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_43),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_50),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_45),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_47),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_66),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_56),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_61),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_20),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_97),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_14),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_43),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_103),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_117),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_30),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_59),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_58),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_24),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_42),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_76),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_44),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_22),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_136),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_7),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_69),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_31),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_77),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_26),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_92),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_134),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_98),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_113),
.Y(n_249)
);

INVx4_ASAP7_75t_R g250 ( 
.A(n_53),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_10),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_49),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_67),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_55),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_109),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_23),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_91),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_54),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_96),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_31),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_143),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_89),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_26),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_124),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_138),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_63),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_73),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_106),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_41),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_3),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_6),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_68),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_126),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_51),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_72),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_133),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_14),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_75),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_25),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_209),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_172),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_155),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_209),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_227),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_152),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_239),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_276),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_152),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_224),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_224),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_267),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_287),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_287),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_224),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_200),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_236),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_150),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_203),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_211),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_150),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_241),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_156),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_163),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_163),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_157),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_258),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_161),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_161),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_161),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_268),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_170),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_170),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_170),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_159),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_149),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_257),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_221),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_273),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_173),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_185),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_188),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_189),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_190),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_154),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_191),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_194),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_204),
.B(n_199),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_154),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_183),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_313),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_303),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_171),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_171),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_313),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_231),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_266),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_314),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_305),
.A2(n_186),
.B1(n_180),
.B2(n_238),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_340),
.A2(n_186),
.B1(n_180),
.B2(n_238),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_177),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_348),
.B(n_159),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_314),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_351),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_207),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_320),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_308),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_310),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_316),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_325),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_328),
.B(n_214),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_326),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_315),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_299),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_296),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_332),
.B(n_301),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_312),
.B(n_348),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_297),
.B(n_262),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_324),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_361),
.B(n_177),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_355),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_354),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_352),
.B(n_354),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_341),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_352),
.B(n_216),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_371),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_305),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_302),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_383),
.B(n_183),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_307),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_373),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_371),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_302),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_183),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_382),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_433),
.B(n_342),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_421),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_371),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_307),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_346),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_165),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_374),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_350),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_380),
.B(n_160),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_389),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_378),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_380),
.B(n_424),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_423),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_369),
.A2(n_368),
.B1(n_323),
.B2(n_321),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_383),
.B(n_362),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_369),
.A2(n_367),
.B1(n_365),
.B2(n_364),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_372),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_432),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_407),
.B(n_363),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_380),
.B(n_424),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_SL g490 ( 
.A1(n_436),
.A2(n_365),
.B(n_364),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

AND2x4_ASAP7_75t_SL g494 ( 
.A(n_380),
.B(n_165),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_384),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_397),
.B(n_160),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_372),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_372),
.B(n_182),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_397),
.B(n_298),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_369),
.A2(n_333),
.B1(n_329),
.B2(n_330),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_397),
.B(n_331),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_432),
.B(n_334),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_394),
.Y(n_512)
);

INVx6_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_372),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_436),
.B(n_335),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_394),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_381),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_417),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_435),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_386),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_399),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_431),
.B(n_336),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_400),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_429),
.B(n_265),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_375),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_402),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_431),
.B(n_162),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_381),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_413),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_431),
.B(n_337),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_381),
.B(n_339),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_372),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_431),
.B(n_162),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_420),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_369),
.A2(n_345),
.B1(n_344),
.B2(n_343),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_422),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_420),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_426),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_420),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_381),
.B(n_426),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_426),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_386),
.B(n_166),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_415),
.Y(n_555)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_419),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_372),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_372),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_385),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_390),
.B(n_198),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_403),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_393),
.B(n_164),
.C(n_169),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_412),
.Y(n_563)
);

AND3x2_ASAP7_75t_L g564 ( 
.A(n_395),
.B(n_217),
.C(n_178),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_379),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_410),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_430),
.B(n_166),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_L g569 ( 
.A(n_395),
.B(n_182),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_411),
.B(n_327),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_421),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_380),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_437),
.B(n_167),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_425),
.B(n_167),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_370),
.Y(n_575)
);

AND2x2_ASAP7_75t_SL g576 ( 
.A(n_424),
.B(n_223),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_406),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_425),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_370),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_561),
.B(n_265),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_184),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_552),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_441),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_514),
.B(n_279),
.Y(n_587)
);

O2A1O1Ixp33_ASAP7_75t_L g588 ( 
.A1(n_490),
.A2(n_439),
.B(n_453),
.C(n_447),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_499),
.B(n_576),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_441),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_561),
.B(n_327),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_488),
.B(n_279),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_450),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_499),
.B(n_281),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_470),
.B(n_281),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_453),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_499),
.B(n_242),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_456),
.B(n_445),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_464),
.A2(n_576),
.B1(n_545),
.B2(n_483),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_555),
.B(n_193),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_438),
.B(n_210),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_469),
.A2(n_226),
.B(n_292),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_169),
.C(n_157),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_569),
.A2(n_153),
.B1(n_254),
.B2(n_164),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_566),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_438),
.B(n_578),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_578),
.B(n_215),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_545),
.B(n_219),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_524),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_545),
.B(n_220),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_510),
.B(n_222),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_514),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_466),
.B(n_158),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_444),
.B(n_230),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_234),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_524),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_480),
.B(n_235),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_240),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_528),
.A2(n_282),
.B1(n_158),
.B2(n_283),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_483),
.B(n_248),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_483),
.B(n_251),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_560),
.B(n_283),
.C(n_284),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_443),
.B(n_252),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_475),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_561),
.B(n_284),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_449),
.A2(n_153),
.B1(n_225),
.B2(n_289),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_523),
.B(n_271),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_557),
.B(n_237),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_530),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_557),
.B(n_244),
.Y(n_636)
);

AND2x4_ASAP7_75t_SL g637 ( 
.A(n_572),
.B(n_245),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_569),
.B(n_501),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_443),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_449),
.A2(n_254),
.B1(n_288),
.B2(n_259),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_572),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_492),
.B(n_285),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_454),
.B(n_293),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_475),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_L g645 ( 
.A(n_449),
.B(n_182),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_449),
.A2(n_280),
.B1(n_255),
.B2(n_182),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_476),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_463),
.B(n_1),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_4),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_530),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_534),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_566),
.B(n_7),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_448),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_558),
.B(n_182),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_534),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_440),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_484),
.A2(n_175),
.B1(n_286),
.B2(n_275),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_449),
.A2(n_174),
.B1(n_274),
.B2(n_270),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_518),
.B(n_151),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_482),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_462),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_457),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_440),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_482),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_536),
.A2(n_291),
.B(n_269),
.C(n_264),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_457),
.A2(n_463),
.B1(n_551),
.B2(n_467),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_494),
.B(n_8),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_520),
.B(n_533),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_518),
.B(n_263),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_481),
.B(n_256),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_520),
.B(n_253),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_497),
.B(n_11),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_457),
.A2(n_182),
.B1(n_249),
.B2(n_247),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_515),
.B(n_549),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_532),
.B(n_541),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_565),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_565),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_457),
.A2(n_485),
.B1(n_558),
.B2(n_505),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_520),
.B(n_533),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_529),
.B(n_568),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_570),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_570),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_SL g684 ( 
.A(n_529),
.B(n_233),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_457),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_496),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_496),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_559),
.B(n_205),
.C(n_246),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_515),
.B(n_232),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_179),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_570),
.Y(n_691)
);

BUFx6f_ASAP7_75t_SL g692 ( 
.A(n_568),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_462),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_571),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_574),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_548),
.B(n_181),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_471),
.A2(n_202),
.B1(n_229),
.B2(n_228),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_548),
.B(n_197),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_573),
.B(n_554),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_533),
.B(n_182),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_550),
.B(n_187),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_550),
.B(n_192),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_556),
.A2(n_579),
.B1(n_498),
.B2(n_575),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_504),
.B(n_11),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_498),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_442),
.B(n_208),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_502),
.A2(n_218),
.B1(n_213),
.B2(n_212),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_502),
.A2(n_201),
.B1(n_196),
.B2(n_195),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_458),
.B(n_12),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_503),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_503),
.A2(n_250),
.B(n_48),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_577),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_511),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_511),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_571),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_446),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_486),
.B(n_12),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_512),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_568),
.Y(n_719)
);

OAI21xp33_ASAP7_75t_L g720 ( 
.A1(n_512),
.A2(n_15),
.B(n_16),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_486),
.B(n_537),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_516),
.B(n_17),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_570),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_516),
.A2(n_579),
.B(n_575),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_506),
.B(n_21),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_517),
.B(n_25),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_567),
.B(n_27),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_486),
.B(n_29),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_486),
.B(n_29),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_526),
.B(n_32),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_535),
.B(n_460),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_477),
.B(n_34),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_517),
.Y(n_733)
);

BUFx12f_ASAP7_75t_L g734 ( 
.A(n_715),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_685),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_653),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_599),
.B(n_525),
.Y(n_739)
);

HB1xp67_ASAP7_75t_SL g740 ( 
.A(n_662),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_656),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_599),
.B(n_563),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_586),
.B(n_590),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_597),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_525),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_602),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_604),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_615),
.B(n_622),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_638),
.B(n_609),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_664),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_593),
.B(n_559),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_581),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_613),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_630),
.B(n_644),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_659),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_653),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_661),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_601),
.B(n_563),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_665),
.B(n_527),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_663),
.B(n_489),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_686),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_687),
.B(n_527),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_693),
.A2(n_564),
.B1(n_513),
.B2(n_546),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_705),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_710),
.B(n_542),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_713),
.B(n_542),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_663),
.B(n_487),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_714),
.B(n_540),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_663),
.B(n_487),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_663),
.B(n_486),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_718),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_733),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_583),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_675),
.B(n_540),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_619),
.B(n_547),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_724),
.B(n_543),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_584),
.A2(n_513),
.B1(n_501),
.B2(n_538),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_667),
.B(n_731),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_694),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_610),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_611),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_692),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_633),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_712),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_685),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_652),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_695),
.B(n_543),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_SL g788 ( 
.A(n_684),
.B(n_538),
.C(n_531),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_581),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_638),
.B(n_539),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_719),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_635),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_650),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_580),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_651),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_588),
.A2(n_531),
.B(n_553),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_677),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_589),
.B(n_547),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_654),
.A2(n_544),
.B(n_459),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_584),
.B(n_513),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_581),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_655),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_641),
.B(n_537),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_716),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_585),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_606),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_653),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_653),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_703),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_685),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_589),
.A2(n_493),
.B1(n_446),
.B2(n_522),
.Y(n_812)
);

OR2x2_ASAP7_75t_SL g813 ( 
.A(n_727),
.B(n_553),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_731),
.B(n_679),
.Y(n_814)
);

BUFx4f_ASAP7_75t_L g815 ( 
.A(n_637),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_725),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_730),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_704),
.Y(n_818)
);

OAI22xp33_ASAP7_75t_L g819 ( 
.A1(n_592),
.A2(n_461),
.B1(n_473),
.B2(n_478),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_591),
.B(n_537),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_591),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_639),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_654),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_607),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_639),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_607),
.Y(n_827)
);

NOR2x1_ASAP7_75t_L g828 ( 
.A(n_641),
.B(n_461),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_649),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_692),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_668),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_634),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_679),
.B(n_493),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_681),
.B(n_537),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_596),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_699),
.B(n_461),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_682),
.B(n_537),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_625),
.B(n_683),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_596),
.B(n_448),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_609),
.A2(n_473),
.B1(n_478),
.B2(n_519),
.Y(n_841)
);

AND2x6_ASAP7_75t_L g842 ( 
.A(n_596),
.B(n_448),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_648),
.Y(n_843)
);

OR2x2_ASAP7_75t_SL g844 ( 
.A(n_625),
.B(n_522),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_603),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_723),
.B(n_521),
.Y(n_846)
);

NAND2x1p5_ASAP7_75t_L g847 ( 
.A(n_596),
.B(n_473),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_720),
.A2(n_521),
.B1(n_519),
.B2(n_509),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_620),
.B(n_509),
.Y(n_849)
);

AND2x6_ASAP7_75t_L g850 ( 
.A(n_618),
.B(n_448),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_673),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_726),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_699),
.B(n_478),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_631),
.B(n_448),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_620),
.A2(n_452),
.B1(n_507),
.B2(n_500),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_676),
.B(n_508),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_709),
.A2(n_673),
.B(n_647),
.C(n_595),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_605),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_689),
.B(n_612),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_732),
.B(n_618),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_618),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_636),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_621),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_676),
.B(n_508),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_732),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_608),
.A2(n_507),
.B1(n_500),
.B2(n_495),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_618),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_623),
.Y(n_869)
);

BUFx8_ASAP7_75t_SL g870 ( 
.A(n_614),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_628),
.B(n_495),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_SL g872 ( 
.A1(n_640),
.A2(n_452),
.B1(n_35),
.B2(n_38),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_624),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_690),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_626),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_627),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_680),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_688),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_642),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_616),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_629),
.B(n_643),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_696),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_680),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_669),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_629),
.B(n_452),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_672),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_632),
.B(n_452),
.Y(n_887)
);

INVx6_ASAP7_75t_L g888 ( 
.A(n_717),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_698),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_643),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_701),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_594),
.A2(n_491),
.B(n_479),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_717),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_728),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_608),
.A2(n_491),
.B1(n_479),
.B2(n_474),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_617),
.B(n_474),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_702),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_640),
.B(n_472),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_671),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_646),
.B(n_472),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_658),
.B(n_465),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_707),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_707),
.B(n_465),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_729),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_803),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_881),
.A2(n_729),
.B(n_594),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_890),
.B(n_657),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_815),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_785),
.B(n_700),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_736),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_738),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_815),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_885),
.A2(n_700),
.B(n_598),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_739),
.B(n_646),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_785),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_739),
.A2(n_587),
.B(n_645),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_744),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_708),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_779),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_776),
.A2(n_598),
.B(n_660),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_749),
.A2(n_674),
.B1(n_708),
.B2(n_666),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_751),
.B(n_657),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_866),
.B(n_674),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_776),
.A2(n_670),
.B(n_706),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_866),
.B(n_697),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_785),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_822),
.B(n_721),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_748),
.B(n_711),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_746),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_747),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_753),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_755),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_773),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_SL g934 ( 
.A(n_734),
.B(n_34),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_851),
.B(n_35),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_735),
.Y(n_936)
);

OAI22x1_ASAP7_75t_L g937 ( 
.A1(n_851),
.A2(n_794),
.B1(n_818),
.B2(n_820),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_818),
.A2(n_38),
.B(n_40),
.C(n_41),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_749),
.A2(n_60),
.B1(n_70),
.B2(n_83),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_737),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_774),
.A2(n_88),
.B(n_93),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_780),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_757),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_737),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_814),
.B(n_115),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_735),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_859),
.B(n_128),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_820),
.A2(n_132),
.B1(n_139),
.B2(n_140),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_736),
.B(n_141),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_758),
.A2(n_796),
.B(n_892),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_782),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_780),
.Y(n_952)
);

OAI22x1_ASAP7_75t_L g953 ( 
.A1(n_902),
.A2(n_786),
.B1(n_874),
.B2(n_886),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_787),
.B(n_790),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_SL g955 ( 
.A(n_838),
.B(n_788),
.C(n_858),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_740),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_742),
.A2(n_858),
.B(n_860),
.C(n_843),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_810),
.B(n_775),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_830),
.B(n_845),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_787),
.A2(n_800),
.B(n_790),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_SL g961 ( 
.A1(n_872),
.A2(n_763),
.B1(n_844),
.B2(n_783),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_SL g962 ( 
.A(n_811),
.B(n_904),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_745),
.A2(n_762),
.B(n_759),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_740),
.B(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_882),
.B(n_889),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_880),
.A2(n_879),
.B(n_869),
.C(n_864),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_SL g967 ( 
.A1(n_813),
.A2(n_904),
.B1(n_786),
.B2(n_888),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_743),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_891),
.B(n_754),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_745),
.A2(n_766),
.B(n_765),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_737),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_799),
.A2(n_796),
.B(n_892),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_761),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_764),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_897),
.B(n_875),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_771),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_797),
.B(n_801),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_759),
.A2(n_766),
.B(n_768),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_762),
.A2(n_765),
.B(n_768),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_SL g980 ( 
.A1(n_852),
.A2(n_853),
.B(n_778),
.C(n_816),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_SL g981 ( 
.A1(n_873),
.A2(n_876),
.B(n_817),
.C(n_836),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_772),
.Y(n_982)
);

CKINVDCx10_ASAP7_75t_R g983 ( 
.A(n_904),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_829),
.B(n_831),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_811),
.B(n_804),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_883),
.B(n_854),
.Y(n_986)
);

CKINVDCx16_ASAP7_75t_R g987 ( 
.A(n_878),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_756),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_781),
.B(n_823),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_777),
.A2(n_888),
.B1(n_788),
.B2(n_849),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_840),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_888),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_781),
.B(n_826),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_804),
.B(n_877),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_883),
.B(n_877),
.Y(n_995)
);

O2A1O1Ixp5_ASAP7_75t_L g996 ( 
.A1(n_855),
.A2(n_819),
.B(n_849),
.C(n_876),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_857),
.B(n_865),
.Y(n_997)
);

AO221x1_ASAP7_75t_L g998 ( 
.A1(n_894),
.A2(n_819),
.B1(n_873),
.B2(n_883),
.C(n_899),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_837),
.B(n_884),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_884),
.B(n_846),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_870),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_805),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_806),
.B(n_807),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_893),
.Y(n_1004)
);

NOR2xp67_ASAP7_75t_L g1005 ( 
.A(n_871),
.B(n_865),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_SL g1006 ( 
.A(n_862),
.B(n_868),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_SL g1007 ( 
.A(n_756),
.B(n_808),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_792),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_857),
.B(n_795),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_828),
.B(n_760),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_861),
.B(n_899),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_893),
.Y(n_1012)
);

OAI211xp5_ASAP7_75t_L g1013 ( 
.A1(n_867),
.A2(n_895),
.B(n_903),
.C(n_856),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_793),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_R g1015 ( 
.A(n_808),
.B(n_809),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_894),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_896),
.A2(n_863),
.B(n_901),
.C(n_798),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_802),
.A2(n_798),
.B(n_834),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_741),
.B(n_750),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_784),
.B(n_832),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_802),
.A2(n_833),
.B(n_821),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_808),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_841),
.A2(n_812),
.B(n_848),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_833),
.A2(n_898),
.B1(n_848),
.B2(n_900),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_824),
.B(n_809),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_825),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_809),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_900),
.A2(n_898),
.B(n_769),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_812),
.B(n_827),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_752),
.B(n_789),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_SL g1031 ( 
.A(n_887),
.B(n_868),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_847),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_752),
.B(n_789),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_835),
.B(n_862),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_887),
.B(n_835),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_R g1036 ( 
.A(n_862),
.B(n_839),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_839),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_767),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_767),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_985),
.B(n_770),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_936),
.B(n_946),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_972),
.A2(n_839),
.B(n_842),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_951),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_1024),
.A2(n_887),
.A3(n_842),
.B(n_850),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_969),
.B(n_887),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_950),
.A2(n_842),
.B(n_850),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_965),
.B(n_975),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_960),
.A2(n_842),
.B(n_850),
.Y(n_1048)
);

BUFx4_ASAP7_75t_SL g1049 ( 
.A(n_1001),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_922),
.A2(n_850),
.B(n_923),
.C(n_921),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_SL g1051 ( 
.A1(n_935),
.A2(n_850),
.B(n_918),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_961),
.A2(n_955),
.B1(n_921),
.B2(n_967),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_914),
.A2(n_978),
.B(n_970),
.Y(n_1053)
);

AOI31xp67_ASAP7_75t_L g1054 ( 
.A1(n_928),
.A2(n_945),
.A3(n_986),
.B(n_997),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_911),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1002),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_933),
.B(n_956),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_964),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_R g1059 ( 
.A(n_908),
.B(n_912),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_957),
.A2(n_966),
.B(n_925),
.C(n_979),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_996),
.A2(n_914),
.B(n_920),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1000),
.B(n_987),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_916),
.A2(n_924),
.B(n_980),
.Y(n_1063)
);

AO31x2_ASAP7_75t_L g1064 ( 
.A1(n_1024),
.A2(n_1029),
.A3(n_1026),
.B(n_906),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_990),
.A2(n_954),
.B(n_945),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1037),
.B(n_994),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_952),
.B(n_942),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1023),
.A2(n_981),
.B(n_939),
.C(n_958),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1021),
.A2(n_1017),
.B(n_1013),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_939),
.A2(n_1005),
.B(n_938),
.C(n_959),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1009),
.B(n_999),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1011),
.A2(n_1025),
.B(n_992),
.C(n_941),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_917),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1031),
.A2(n_962),
.B(n_1018),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_992),
.A2(n_968),
.B1(n_993),
.B2(n_989),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_SL g1076 ( 
.A1(n_913),
.A2(n_1035),
.B(n_1006),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_929),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_984),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_999),
.B(n_1004),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1015),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_930),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_909),
.A2(n_1029),
.B(n_1010),
.Y(n_1082)
);

NOR2xp67_ASAP7_75t_SL g1083 ( 
.A(n_1037),
.B(n_919),
.Y(n_1083)
);

AND3x4_ASAP7_75t_L g1084 ( 
.A(n_983),
.B(n_934),
.C(n_994),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_977),
.B(n_1012),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_991),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_931),
.B(n_976),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1038),
.A2(n_1032),
.B(n_995),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_948),
.A2(n_1020),
.B(n_910),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_1037),
.B(n_949),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_985),
.Y(n_1091)
);

INVx5_ASAP7_75t_L g1092 ( 
.A(n_949),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_937),
.A2(n_1003),
.A3(n_1014),
.B(n_1008),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_962),
.B(n_1027),
.Y(n_1094)
);

CKINVDCx11_ASAP7_75t_R g1095 ( 
.A(n_949),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_927),
.A2(n_982),
.B(n_974),
.C(n_973),
.Y(n_1096)
);

AOI211x1_ASAP7_75t_L g1097 ( 
.A1(n_932),
.A2(n_943),
.B(n_948),
.C(n_947),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_1007),
.B(n_915),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1016),
.B(n_1036),
.C(n_1033),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_SL g1100 ( 
.A1(n_927),
.A2(n_1019),
.B(n_998),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1039),
.C(n_1022),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_988),
.Y(n_1102)
);

NAND3x1_ASAP7_75t_L g1103 ( 
.A(n_953),
.B(n_915),
.C(n_926),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_940),
.B(n_944),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_940),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_944),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_926),
.A2(n_971),
.B(n_988),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_971),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_907),
.A2(n_599),
.B1(n_820),
.B2(n_818),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_SL g1111 ( 
.A(n_907),
.B(n_385),
.C(n_375),
.Y(n_1111)
);

AOI221x1_ASAP7_75t_L g1112 ( 
.A1(n_955),
.A2(n_939),
.B1(n_921),
.B2(n_599),
.C(n_961),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_969),
.B(n_599),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_1001),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_969),
.B(n_599),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_950),
.A2(n_924),
.B(n_920),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_985),
.B(n_908),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_1037),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_963),
.A2(n_739),
.B(n_970),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_936),
.B(n_583),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_907),
.B(n_890),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_955),
.B(n_599),
.C(n_922),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_907),
.A2(n_314),
.B1(n_316),
.B2(n_313),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_905),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_963),
.A2(n_739),
.B(n_970),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_936),
.B(n_583),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_969),
.B(n_599),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_963),
.A2(n_739),
.B(n_970),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1024),
.A2(n_825),
.A3(n_827),
.B(n_1029),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_911),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_936),
.B(n_583),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_922),
.A2(n_599),
.B(n_866),
.C(n_881),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1037),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_907),
.A2(n_599),
.B1(n_820),
.B2(n_818),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_969),
.B(n_599),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_969),
.B(n_599),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_933),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_907),
.B(n_599),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_969),
.B(n_599),
.Y(n_1143)
);

AOI31xp67_ASAP7_75t_L g1144 ( 
.A1(n_928),
.A2(n_885),
.A3(n_758),
.B(n_945),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_963),
.A2(n_739),
.B(n_970),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_907),
.A2(n_599),
.B(n_820),
.C(n_818),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_907),
.B(n_890),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_911),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_969),
.B(n_599),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_911),
.Y(n_1150)
);

OAI22x1_ASAP7_75t_L g1151 ( 
.A1(n_907),
.A2(n_314),
.B1(n_316),
.B2(n_313),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_911),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_933),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_905),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_963),
.A2(n_739),
.B(n_970),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_1001),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_933),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1037),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_1001),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_911),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_972),
.A2(n_950),
.B(n_1028),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_969),
.B(n_599),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_907),
.B(n_890),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_951),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_961),
.A2(n_599),
.B1(n_749),
.B2(n_907),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_907),
.B(n_890),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1037),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_933),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1024),
.A2(n_825),
.A3(n_827),
.B(n_1029),
.Y(n_1169)
);

AOI221x1_ASAP7_75t_L g1170 ( 
.A1(n_955),
.A2(n_939),
.B1(n_921),
.B2(n_599),
.C(n_961),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1165),
.A2(n_1052),
.B1(n_1112),
.B2(n_1170),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1087),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1117),
.A2(n_1113),
.B(n_1110),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1141),
.B(n_1079),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1058),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1131),
.A2(n_1139),
.B(n_1135),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1164),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_1121),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1067),
.Y(n_1179)
);

INVx5_ASAP7_75t_SL g1180 ( 
.A(n_1090),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1120),
.A2(n_1155),
.A3(n_1145),
.B(n_1129),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_R g1182 ( 
.A(n_1095),
.B(n_1115),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1161),
.A2(n_1053),
.B(n_1061),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1142),
.A2(n_1137),
.B1(n_1109),
.B2(n_1123),
.C(n_1151),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1046),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1055),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1165),
.A2(n_1052),
.B1(n_1124),
.B2(n_1147),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1114),
.B(n_1116),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1071),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1064),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1128),
.B(n_1138),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_1092),
.B(n_1086),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1064),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1146),
.A2(n_1111),
.B(n_1134),
.C(n_1122),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1051),
.A2(n_1042),
.B(n_1126),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1073),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1140),
.A2(n_1162),
.B1(n_1149),
.B2(n_1143),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1091),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1127),
.B(n_1133),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1119),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1062),
.B(n_1041),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_R g1203 ( 
.A(n_1043),
.B(n_1092),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1064),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_1060),
.A2(n_1070),
.B(n_1166),
.C(n_1163),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1168),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1090),
.B(n_1119),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1153),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1141),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1069),
.A2(n_1074),
.B(n_1048),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1119),
.B(n_1158),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1083),
.B(n_1080),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1069),
.A2(n_1048),
.B(n_1089),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1075),
.A2(n_1157),
.B(n_1050),
.C(n_1072),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1078),
.B(n_1057),
.Y(n_1215)
);

OAI211xp5_ASAP7_75t_L g1216 ( 
.A1(n_1097),
.A2(n_1085),
.B(n_1096),
.C(n_1047),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1076),
.A2(n_1045),
.B(n_1082),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1077),
.A2(n_1148),
.A3(n_1081),
.B(n_1152),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1132),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1105),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1156),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1100),
.A2(n_1088),
.B(n_1103),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1150),
.B(n_1160),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1094),
.A2(n_1101),
.B(n_1099),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1136),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1107),
.A2(n_1158),
.B(n_1098),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1049),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1091),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1156),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_1097),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1108),
.A2(n_1102),
.B(n_1066),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1108),
.A2(n_1040),
.B(n_1104),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1056),
.A2(n_1154),
.B(n_1125),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1044),
.A2(n_1118),
.B(n_1169),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1044),
.A2(n_1169),
.B(n_1130),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1169),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1093),
.A2(n_1106),
.B(n_1167),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1091),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1136),
.B(n_1167),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1105),
.B(n_1059),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1084),
.B(n_1159),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1087),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1164),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1142),
.A2(n_599),
.B(n_1123),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1165),
.B(n_1142),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1142),
.A2(n_310),
.B1(n_308),
.B2(n_303),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1087),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1249)
);

NAND2x1p5_ASAP7_75t_L g1250 ( 
.A(n_1092),
.B(n_1119),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1168),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1165),
.A2(n_1052),
.B1(n_1112),
.B2(n_1170),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1142),
.B(n_1165),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1087),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1168),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1064),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1064),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1092),
.B(n_956),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1142),
.B(n_1114),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1142),
.A2(n_599),
.B(n_1123),
.Y(n_1263)
);

NAND2x1p5_ASAP7_75t_L g1264 ( 
.A(n_1092),
.B(n_1119),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1165),
.A2(n_1052),
.B1(n_1112),
.B2(n_1170),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1164),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1142),
.A2(n_599),
.B(n_1146),
.C(n_1137),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1058),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1068),
.A2(n_1024),
.A3(n_1065),
.B(n_1112),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1119),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1087),
.Y(n_1272)
);

OAI221xp5_ASAP7_75t_L g1273 ( 
.A1(n_1142),
.A2(n_599),
.B1(n_1165),
.B2(n_580),
.C(n_467),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1087),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1064),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1168),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1068),
.A2(n_1024),
.A3(n_1065),
.B(n_1112),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1142),
.A2(n_599),
.B(n_1123),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1142),
.A2(n_1165),
.B(n_599),
.C(n_1123),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1142),
.B(n_1165),
.Y(n_1280)
);

OAI222xp33_ASAP7_75t_L g1281 ( 
.A1(n_1165),
.A2(n_393),
.B1(n_1052),
.B2(n_340),
.C1(n_341),
.C2(n_314),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1164),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1164),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1064),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1092),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1142),
.B(n_1114),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1168),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1063),
.A2(n_1117),
.B(n_1113),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1071),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1064),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1063),
.A2(n_1113),
.B(n_1110),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1087),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1142),
.A2(n_961),
.B1(n_1165),
.B2(n_395),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1087),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1279),
.A2(n_1263),
.B(n_1245),
.C(n_1278),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1253),
.A2(n_1280),
.B1(n_1279),
.B2(n_1273),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1268),
.A2(n_1253),
.B(n_1280),
.C(n_1184),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1192),
.B(n_1207),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1246),
.B(n_1198),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1200),
.B(n_1202),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1246),
.B(n_1179),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1242),
.A2(n_1256),
.B(n_1249),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1293),
.A2(n_1187),
.B1(n_1265),
.B2(n_1252),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_SL g1304 ( 
.A(n_1224),
.B(n_1216),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1171),
.A2(n_1281),
.B(n_1195),
.C(n_1205),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1191),
.B(n_1243),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1206),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1221),
.B(n_1229),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1178),
.B(n_1215),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1218),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1192),
.B(n_1207),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1251),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1293),
.A2(n_1187),
.B1(n_1262),
.B2(n_1286),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1248),
.B(n_1254),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1255),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1276),
.B(n_1209),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1192),
.B(n_1207),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1174),
.B(n_1287),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1272),
.B(n_1274),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_SL g1322 ( 
.A1(n_1188),
.A2(n_1185),
.B(n_1214),
.C(n_1275),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1189),
.B(n_1289),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1223),
.B(n_1186),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1205),
.B(n_1247),
.C(n_1230),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1208),
.B(n_1175),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1197),
.B(n_1219),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1175),
.B(n_1269),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1269),
.B(n_1220),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1227),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1212),
.A2(n_1240),
.B(n_1241),
.C(n_1210),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1233),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1241),
.B(n_1199),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1237),
.Y(n_1338)
);

AOI221xp5_ASAP7_75t_L g1339 ( 
.A1(n_1210),
.A2(n_1282),
.B1(n_1244),
.B2(n_1177),
.C(n_1266),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1199),
.B(n_1238),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1212),
.A2(n_1240),
.B(n_1283),
.C(n_1285),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1283),
.A2(n_1266),
.B1(n_1282),
.B2(n_1177),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1244),
.A2(n_1193),
.B1(n_1180),
.B2(n_1261),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1227),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1285),
.B(n_1238),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1183),
.B(n_1257),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1221),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1203),
.A2(n_1264),
.B(n_1250),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_1229),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1225),
.A2(n_1264),
.B(n_1250),
.C(n_1230),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1180),
.A2(n_1230),
.B1(n_1239),
.B2(n_1228),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1211),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1225),
.A2(n_1190),
.B(n_1257),
.C(n_1259),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1201),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1232),
.B(n_1231),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1190),
.B(n_1194),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1194),
.B(n_1275),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1204),
.B(n_1290),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1201),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1182),
.A2(n_1211),
.B(n_1271),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1204),
.A2(n_1284),
.B(n_1239),
.C(n_1217),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1196),
.A2(n_1181),
.B(n_1213),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1217),
.B(n_1213),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1234),
.B(n_1235),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1291),
.A2(n_1236),
.B(n_1176),
.C(n_1235),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1234),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1176),
.A2(n_1235),
.B(n_1181),
.C(n_1222),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1176),
.A2(n_1181),
.B(n_1222),
.C(n_1196),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1181),
.B(n_1226),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1201),
.B(n_1271),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1258),
.A2(n_1260),
.B(n_1267),
.C(n_1288),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1173),
.A2(n_1279),
.B(n_1170),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1279),
.A2(n_599),
.B(n_1142),
.C(n_1245),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1253),
.A2(n_1142),
.B1(n_1280),
.B2(n_1165),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1242),
.A2(n_1256),
.B(n_1249),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1251),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1336),
.B(n_1329),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1346),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1364),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1363),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1369),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1329),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1330),
.B(n_1335),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1334),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1302),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1302),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1311),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1365),
.A2(n_1367),
.B(n_1372),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1368),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1327),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1344),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1362),
.A2(n_1371),
.B(n_1361),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1299),
.B(n_1319),
.Y(n_1393)
);

NOR2x1_ASAP7_75t_R g1394 ( 
.A(n_1299),
.B(n_1328),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1300),
.B(n_1366),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1301),
.B(n_1355),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1347),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1322),
.A2(n_1374),
.B(n_1338),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1296),
.A2(n_1304),
.A3(n_1357),
.B(n_1358),
.Y(n_1400)
);

OAI221xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1297),
.A2(n_1373),
.B1(n_1305),
.B2(n_1295),
.C(n_1339),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1375),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1376),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1310),
.B(n_1308),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1325),
.A2(n_1356),
.B(n_1358),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1350),
.A2(n_1351),
.B(n_1353),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1315),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1331),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1317),
.B(n_1326),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1315),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1320),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1339),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1298),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1306),
.B(n_1307),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1396),
.B(n_1306),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1407),
.B(n_1307),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1384),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1387),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1396),
.B(n_1323),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1387),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1396),
.B(n_1295),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1379),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1407),
.B(n_1321),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1386),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1396),
.B(n_1337),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1407),
.B(n_1352),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1392),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1387),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1392),
.A2(n_1370),
.B(n_1345),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1401),
.A2(n_1303),
.B1(n_1314),
.B2(n_1354),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1413),
.A2(n_1312),
.B1(n_1318),
.B2(n_1342),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1403),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1386),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1392),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1387),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1399),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1399),
.B(n_1340),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1406),
.B(n_1312),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1413),
.A2(n_1359),
.B1(n_1343),
.B2(n_1318),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1396),
.B(n_1345),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1391),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1392),
.A2(n_1402),
.B(n_1385),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

INVx2_ASAP7_75t_R g1445 ( 
.A(n_1389),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1380),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1378),
.B(n_1333),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1380),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1386),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1395),
.B(n_1349),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1444),
.B(n_1414),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1424),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1450),
.B(n_1409),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1422),
.B(n_1415),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1417),
.B(n_1399),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1442),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1447),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1432),
.A2(n_1440),
.B1(n_1422),
.B2(n_1447),
.C(n_1401),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1424),
.Y(n_1460)
);

AOI322xp5_ASAP7_75t_L g1461 ( 
.A1(n_1432),
.A2(n_1393),
.A3(n_1377),
.B1(n_1415),
.B2(n_1401),
.C1(n_1383),
.C2(n_1381),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1419),
.Y(n_1462)
);

NAND2xp33_ASAP7_75t_R g1463 ( 
.A(n_1430),
.B(n_1413),
.Y(n_1463)
);

OAI33xp33_ASAP7_75t_L g1464 ( 
.A1(n_1431),
.A2(n_1399),
.A3(n_1390),
.B1(n_1408),
.B2(n_1411),
.B3(n_1412),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1428),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1422),
.B(n_1415),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1438),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1431),
.A2(n_1413),
.B1(n_1405),
.B2(n_1398),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1419),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1413),
.C(n_1389),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1421),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1421),
.Y(n_1472)
);

INVxp67_ASAP7_75t_SL g1473 ( 
.A(n_1446),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1429),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1440),
.A2(n_1413),
.B1(n_1389),
.B2(n_1341),
.C(n_1379),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1418),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1428),
.A2(n_1389),
.B1(n_1408),
.B2(n_1411),
.C(n_1412),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1445),
.A2(n_1413),
.B1(n_1405),
.B2(n_1398),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1428),
.B(n_1413),
.C(n_1380),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1418),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1429),
.Y(n_1481)
);

OAI31xp33_ASAP7_75t_L g1482 ( 
.A1(n_1439),
.A2(n_1381),
.A3(n_1377),
.B(n_1400),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1442),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1436),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1439),
.A2(n_1412),
.B1(n_1411),
.B2(n_1408),
.C(n_1378),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1445),
.A2(n_1405),
.B1(n_1398),
.B2(n_1388),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1445),
.A2(n_1405),
.B1(n_1398),
.B2(n_1388),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1428),
.B(n_1403),
.C(n_1382),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1438),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1450),
.A2(n_1388),
.B1(n_1377),
.B2(n_1398),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1403),
.C(n_1382),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1428),
.A2(n_1412),
.B1(n_1408),
.B2(n_1411),
.C(n_1415),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1437),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1418),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1476),
.Y(n_1495)
);

INVx4_ASAP7_75t_SL g1496 ( 
.A(n_1457),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1476),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1462),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1478),
.A2(n_1434),
.B(n_1449),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1469),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_L g1501 ( 
.A(n_1470),
.B(n_1434),
.C(n_1425),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1478),
.A2(n_1487),
.B(n_1486),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1479),
.A2(n_1394),
.B(n_1443),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1457),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1452),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1468),
.A2(n_1433),
.B(n_1448),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1471),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1451),
.Y(n_1508)
);

NOR2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1455),
.B(n_1450),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1486),
.A2(n_1487),
.B(n_1434),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1397),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1454),
.B(n_1426),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1435),
.C(n_1443),
.Y(n_1514)
);

AND2x6_ASAP7_75t_L g1515 ( 
.A(n_1451),
.B(n_1414),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1474),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1456),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_1435),
.C(n_1443),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1481),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1465),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1451),
.B(n_1426),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1493),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1488),
.A2(n_1425),
.B(n_1434),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1484),
.Y(n_1524)
);

INVx4_ASAP7_75t_SL g1525 ( 
.A(n_1453),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1480),
.Y(n_1526)
);

INVx4_ASAP7_75t_SL g1527 ( 
.A(n_1460),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1480),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1458),
.Y(n_1529)
);

NAND3xp33_ASAP7_75t_SL g1530 ( 
.A(n_1482),
.B(n_1439),
.C(n_1417),
.Y(n_1530)
);

AND2x6_ASAP7_75t_L g1531 ( 
.A(n_1459),
.B(n_1414),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1505),
.B(n_1435),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1498),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1500),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1529),
.B(n_1466),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1504),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1531),
.A2(n_1464),
.B1(n_1475),
.B2(n_1388),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1517),
.B(n_1467),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1521),
.B(n_1489),
.Y(n_1540)
);

NAND2x1_ASAP7_75t_SL g1541 ( 
.A(n_1521),
.B(n_1465),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1531),
.B(n_1492),
.Y(n_1542)
);

NOR3xp33_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1485),
.C(n_1477),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_L g1544 ( 
.A(n_1530),
.B(n_1491),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1507),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1463),
.C(n_1503),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1513),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1508),
.B(n_1426),
.Y(n_1552)
);

NAND4xp25_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1463),
.C(n_1461),
.D(n_1465),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1505),
.A2(n_1435),
.B(n_1439),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1519),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1524),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1504),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1527),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1495),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1531),
.B(n_1416),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1512),
.B(n_1525),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1512),
.B(n_1441),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1531),
.B(n_1416),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1416),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1531),
.B(n_1393),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1393),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1496),
.B(n_1393),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1496),
.B(n_1448),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1502),
.A2(n_1388),
.B1(n_1405),
.B2(n_1435),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1495),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1502),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1497),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1497),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1545),
.B(n_1397),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1558),
.B(n_1496),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1545),
.B(n_1397),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1496),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1538),
.B(n_1506),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1535),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1547),
.A2(n_1503),
.B1(n_1520),
.B2(n_1437),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1571),
.B(n_1473),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1550),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1558),
.B(n_1525),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1550),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1551),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1551),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1539),
.B(n_1417),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1544),
.A2(n_1520),
.B1(n_1437),
.B2(n_1435),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1555),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1555),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1539),
.B(n_1438),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1556),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1556),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1533),
.B(n_1446),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1546),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1536),
.B(n_1390),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1534),
.B(n_1391),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1561),
.B(n_1525),
.Y(n_1601)
);

OAI31xp33_ASAP7_75t_L g1602 ( 
.A1(n_1553),
.A2(n_1501),
.A3(n_1510),
.B(n_1526),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1536),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

NAND2x1_ASAP7_75t_L g1605 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1537),
.B(n_1420),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1559),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1578),
.A2(n_1602),
.B1(n_1569),
.B2(n_1542),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1580),
.A2(n_1565),
.B1(n_1560),
.B2(n_1564),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1598),
.B(n_1511),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1548),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1577),
.A2(n_1510),
.B1(n_1532),
.B2(n_1567),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1589),
.A2(n_1435),
.B1(n_1388),
.B2(n_1445),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1603),
.B(n_1540),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1587),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1588),
.B(n_1599),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1590),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1591),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1579),
.B(n_1540),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1598),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1593),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1309),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1601),
.B(n_1549),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1581),
.B(n_1527),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1599),
.B(n_1562),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1607),
.A2(n_1388),
.B1(n_1532),
.B2(n_1405),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1613),
.B(n_1618),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1621),
.Y(n_1635)
);

AOI32xp33_ASAP7_75t_L g1636 ( 
.A1(n_1609),
.A2(n_1607),
.A3(n_1581),
.B1(n_1584),
.B2(n_1594),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1621),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1623),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1633),
.A2(n_1608),
.B1(n_1604),
.B2(n_1596),
.C(n_1554),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1610),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1620),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1627),
.A2(n_1568),
.B(n_1576),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1627),
.B(n_1574),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1623),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1592),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1631),
.B(n_1605),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1611),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1574),
.C(n_1576),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1630),
.A2(n_1631),
.B1(n_1615),
.B2(n_1610),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1630),
.B(n_1595),
.C(n_1499),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.B(n_1562),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1616),
.A2(n_1614),
.B1(n_1617),
.B2(n_1563),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1612),
.C(n_1622),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1641),
.B(n_1629),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1651),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1629),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1652),
.B(n_1632),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1640),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1649),
.B(n_1624),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1638),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1653),
.A2(n_1570),
.B1(n_1573),
.B2(n_1572),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1644),
.B(n_1625),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1660),
.A2(n_1634),
.B(n_1642),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1662),
.A2(n_1636),
.B1(n_1639),
.B2(n_1653),
.C(n_1650),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1654),
.B(n_1642),
.C(n_1645),
.D(n_1647),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1663),
.A2(n_1637),
.B(n_1635),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1655),
.B(n_1646),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1646),
.B(n_1628),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1661),
.Y(n_1670)
);

AOI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1663),
.A2(n_1572),
.B(n_1573),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1658),
.B(n_1597),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1664),
.B(n_1657),
.C(n_1332),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1672),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1665),
.A2(n_1629),
.B1(n_1600),
.B2(n_1570),
.Y(n_1675)
);

AOI211xp5_ASAP7_75t_L g1676 ( 
.A1(n_1666),
.A2(n_1499),
.B(n_1606),
.C(n_1600),
.Y(n_1676)
);

OAI31xp33_ASAP7_75t_L g1677 ( 
.A1(n_1671),
.A2(n_1566),
.A3(n_1527),
.B(n_1528),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1674),
.B(n_1667),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1675),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1669),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1677),
.B(n_1668),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1670),
.Y(n_1683)
);

OAI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1678),
.A2(n_1520),
.B1(n_1528),
.B2(n_1526),
.C1(n_1427),
.C2(n_1423),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1678),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1682),
.Y(n_1686)
);

XNOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1679),
.B(n_1523),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1683),
.Y(n_1688)
);

OR4x2_ASAP7_75t_L g1689 ( 
.A(n_1688),
.B(n_1681),
.C(n_1680),
.D(n_1541),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1685),
.B(n_1541),
.C(n_1427),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_SL g1691 ( 
.A(n_1684),
.B(n_1520),
.C(n_1515),
.Y(n_1691)
);

NAND3x1_ASAP7_75t_L g1692 ( 
.A(n_1689),
.B(n_1686),
.C(n_1687),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1690),
.B1(n_1691),
.B2(n_1385),
.C(n_1494),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1693),
.B(n_1515),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1523),
.B(n_1515),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1694),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1494),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1696),
.A2(n_1433),
.B1(n_1443),
.B2(n_1385),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1697),
.A2(n_1443),
.B1(n_1385),
.B2(n_1404),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1698),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1700),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1701),
.B(n_1699),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1515),
.B1(n_1398),
.B2(n_1410),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1360),
.B(n_1348),
.C(n_1394),
.Y(n_1705)
);


endmodule