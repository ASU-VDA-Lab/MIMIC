module fake_jpeg_1679_n_567 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_567);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_567;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_57),
.Y(n_140)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_64),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_32),
.B(n_0),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_65),
.Y(n_165)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_69),
.B(n_72),
.Y(n_116)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_70),
.Y(n_155)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_92),
.Y(n_157)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_18),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_49),
.Y(n_96)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_105),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_104),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_25),
.B1(n_52),
.B2(n_42),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_108),
.A2(n_142),
.B1(n_144),
.B2(n_24),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_109),
.B(n_118),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_48),
.B1(n_31),
.B2(n_45),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_117),
.A2(n_124),
.B1(n_132),
.B2(n_138),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_25),
.B(n_52),
.C(n_42),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_57),
.A2(n_48),
.B1(n_31),
.B2(n_45),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_47),
.C(n_21),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_126),
.B(n_167),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_48),
.B1(n_31),
.B2(n_54),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_27),
.B1(n_33),
.B2(n_96),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_45),
.B1(n_35),
.B2(n_34),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_55),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_61),
.B1(n_100),
.B2(n_56),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_54),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_38),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_59),
.A2(n_19),
.B1(n_27),
.B2(n_33),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_94),
.B1(n_91),
.B2(n_90),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_67),
.B(n_47),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_111),
.A2(n_27),
.B1(n_33),
.B2(n_22),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_171),
.B(n_182),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_172),
.A2(n_154),
.B1(n_137),
.B2(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_173),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_176),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_177),
.Y(n_279)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_197),
.Y(n_242)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_112),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_188),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_187),
.A2(n_196),
.B1(n_216),
.B2(n_220),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_191),
.B(n_213),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_125),
.B1(n_110),
.B2(n_160),
.Y(n_192)
);

NOR2x1p5_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_114),
.Y(n_256)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_86),
.B1(n_85),
.B2(n_81),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_200),
.B1(n_218),
.B2(n_121),
.Y(n_235)
);

CKINVDCx6p67_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_62),
.B1(n_30),
.B2(n_28),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_209),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_0),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_207),
.B(n_212),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_118),
.A2(n_116),
.B(n_138),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_208),
.A2(n_222),
.B(n_134),
.Y(n_263)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_214),
.Y(n_270)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_113),
.B(n_0),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_110),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_141),
.A2(n_50),
.B1(n_46),
.B2(n_53),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_125),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_53),
.B1(n_50),
.B2(n_46),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_153),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_53),
.B(n_50),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_0),
.Y(n_277)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_114),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_164),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_233),
.B(n_259),
.C(n_265),
.Y(n_310)
);

OA22x2_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_117),
.B1(n_124),
.B2(n_159),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_234),
.A2(n_240),
.B(n_199),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_235),
.A2(n_246),
.B1(n_7),
.B2(n_9),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_203),
.A2(n_161),
.B1(n_121),
.B2(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_147),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_192),
.B1(n_196),
.B2(n_199),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_198),
.B(n_120),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_258),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_134),
.C(n_137),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_220),
.B(n_188),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_181),
.B(n_148),
.C(n_135),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_215),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_156),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_169),
.B(n_135),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_127),
.C(n_156),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_185),
.B(n_156),
.C(n_120),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_177),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_189),
.B(n_175),
.C(n_192),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_286),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_283),
.A2(n_287),
.B1(n_299),
.B2(n_308),
.Y(n_366)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_194),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_248),
.A2(n_192),
.B1(n_196),
.B2(n_175),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_242),
.B(n_233),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_190),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_291),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_193),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_199),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_298),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_301),
.B(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_262),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_248),
.A2(n_196),
.B1(n_175),
.B2(n_219),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_175),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_302),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_201),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_263),
.A2(n_184),
.B(n_211),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_327),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_221),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_312),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_248),
.A2(n_195),
.B1(n_183),
.B2(n_224),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_178),
.B1(n_180),
.B2(n_223),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_316),
.B1(n_317),
.B2(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_229),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_2),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_313),
.B(n_314),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_257),
.A2(n_174),
.B(n_3),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_240),
.B(n_174),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_321),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_256),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_249),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_229),
.Y(n_318)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_5),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_230),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_239),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_241),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_324),
.A2(n_237),
.B1(n_275),
.B2(n_238),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_258),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_325),
.A2(n_231),
.B1(n_254),
.B2(n_252),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_234),
.A2(n_10),
.B(n_11),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_234),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_332),
.Y(n_387)
);

AO22x1_ASAP7_75t_SL g332 ( 
.A1(n_297),
.A2(n_256),
.B1(n_258),
.B2(n_278),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_313),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_341),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_292),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_352),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_345),
.A2(n_354),
.B1(n_370),
.B2(n_316),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_260),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_362),
.C(n_367),
.Y(n_389)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_321),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_299),
.B1(n_287),
.B2(n_283),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_286),
.B(n_276),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_358),
.B(n_371),
.Y(n_392)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_280),
.C(n_272),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_312),
.B(n_265),
.C(n_278),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_291),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_289),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_281),
.B(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_290),
.B(n_270),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_333),
.A2(n_301),
.B(n_304),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_395),
.B(n_396),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_326),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_391),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_354),
.A2(n_327),
.B1(n_328),
.B2(n_306),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_374),
.A2(n_393),
.B1(n_363),
.B2(n_335),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_366),
.A2(n_311),
.B1(n_315),
.B2(n_322),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_379),
.B1(n_383),
.B2(n_384),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_377),
.B(n_332),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_295),
.B1(n_296),
.B2(n_315),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_361),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_380),
.B(n_390),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_281),
.B1(n_305),
.B2(n_293),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_293),
.B1(n_326),
.B2(n_282),
.Y(n_384)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_388),
.B(n_397),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_361),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_371),
.B(n_308),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_282),
.B1(n_309),
.B2(n_303),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_254),
.C(n_261),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_408),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_314),
.B(n_294),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_365),
.A2(n_314),
.B(n_247),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_344),
.A2(n_325),
.B1(n_323),
.B2(n_288),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_398),
.A2(n_344),
.B1(n_338),
.B2(n_364),
.Y(n_418)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_399),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_340),
.B(n_237),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_407),
.Y(n_434)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_359),
.B(n_317),
.Y(n_405)
);

XNOR2x2_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_356),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_358),
.B(n_268),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_335),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_342),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_232),
.C(n_261),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_413),
.Y(n_447)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_400),
.Y(n_415)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_408),
.Y(n_417)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_417),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_418),
.A2(n_433),
.B1(n_398),
.B2(n_386),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_392),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_403),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_420),
.B(n_422),
.Y(n_453)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_403),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_424),
.B(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_356),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_431),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_369),
.Y(n_430)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_432),
.A2(n_435),
.B1(n_442),
.B2(n_345),
.Y(n_460)
);

AOI22x1_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_363),
.B1(n_332),
.B2(n_353),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_388),
.A2(n_353),
.B(n_341),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_387),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_389),
.B(n_392),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_389),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_393),
.A2(n_334),
.B1(n_339),
.B2(n_346),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_383),
.B1(n_374),
.B2(n_376),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_436),
.A2(n_401),
.B1(n_395),
.B2(n_391),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_410),
.A2(n_330),
.B1(n_378),
.B2(n_349),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_469),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_456),
.B(n_471),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_406),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_462),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_416),
.B1(n_413),
.B2(n_409),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_394),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_412),
.B(n_359),
.C(n_401),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_470),
.C(n_417),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_350),
.B1(n_396),
.B2(n_372),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_468),
.B1(n_416),
.B2(n_427),
.Y(n_489)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_467),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_350),
.B1(n_334),
.B2(n_386),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_405),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_425),
.B(n_329),
.C(n_331),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_431),
.B(n_404),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_472),
.B(n_473),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_440),
.C(n_426),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_477),
.B(n_487),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_439),
.Y(n_478)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_428),
.B(n_437),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_479),
.A2(n_490),
.B(n_456),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_443),
.B(n_432),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_443),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_428),
.B(n_426),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_481),
.A2(n_483),
.B(n_484),
.Y(n_503)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_463),
.A2(n_433),
.B(n_435),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_435),
.B(n_434),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_492),
.B1(n_450),
.B2(n_454),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_337),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_488),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_489),
.A2(n_461),
.B1(n_468),
.B2(n_445),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_446),
.A2(n_411),
.B(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_444),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_465),
.B(n_352),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_493),
.B(n_495),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_470),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_494),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_455),
.B(n_329),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_500),
.A2(n_504),
.B(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_484),
.A2(n_452),
.B1(n_471),
.B2(n_441),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_510),
.B1(n_489),
.B2(n_481),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_511),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_459),
.C(n_469),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_507),
.B(n_512),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_479),
.A2(n_441),
.B(n_331),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_508),
.A2(n_476),
.B(n_483),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_475),
.A2(n_360),
.B1(n_357),
.B2(n_355),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_355),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_284),
.C(n_232),
.Y(n_512)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_514),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_497),
.A2(n_490),
.B(n_482),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_516),
.A2(n_518),
.B(n_522),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_530),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_509),
.A2(n_504),
.B(n_503),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_491),
.C(n_474),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_519),
.B(n_520),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_491),
.C(n_480),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_513),
.B(n_498),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_524),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_503),
.A2(n_478),
.B(n_485),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_486),
.C(n_492),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_527),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_501),
.B(n_488),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_266),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_284),
.C(n_236),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_244),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_268),
.B(n_244),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_530),
.A2(n_508),
.B1(n_499),
.B2(n_500),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_540),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_523),
.A2(n_510),
.B1(n_499),
.B2(n_512),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_537),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_517),
.A2(n_247),
.B1(n_238),
.B2(n_266),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_533),
.A2(n_514),
.B1(n_528),
.B2(n_529),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_239),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_16),
.B(n_533),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_13),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_543),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_14),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_525),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_546),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_549),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_535),
.B(n_515),
.C(n_14),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_515),
.C(n_14),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_552),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_16),
.C(n_536),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_542),
.Y(n_557)
);

AO21x1_ASAP7_75t_L g559 ( 
.A1(n_557),
.A2(n_554),
.B(n_548),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_537),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_558),
.A2(n_551),
.B(n_552),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_560),
.Y(n_563)
);

AO21x1_ASAP7_75t_L g561 ( 
.A1(n_555),
.A2(n_538),
.B(n_541),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_561),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_556),
.C(n_544),
.Y(n_564)
);

BUFx24_ASAP7_75t_SL g565 ( 
.A(n_564),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_563),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_545),
.B(n_535),
.Y(n_567)
);


endmodule