module real_jpeg_17786_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_12),
.Y(n_11)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_0),
.A2(n_15),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_2),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_2),
.B(n_5),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_15),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B(n_24),
.C(n_41),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_9),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_9),
.B(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_13),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_22),
.C(n_23),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_28),
.Y(n_27)
);

OR2x4_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B(n_36),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_37),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B(n_50),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);


endmodule