module fake_netlist_6_2272_n_1635 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1635);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1635;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_39),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_68),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_34),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_54),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_14),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_53),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_48),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_94),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_49),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_58),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_9),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_106),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_47),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_4),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_48),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_42),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_30),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_6),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_7),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_5),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_24),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_96),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_101),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_15),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_100),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_17),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_57),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_35),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_75),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_44),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_16),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_66),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_144),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_59),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_46),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_133),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_9),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_38),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_130),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_14),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_142),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_112),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_22),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_34),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_131),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_63),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_126),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_51),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_85),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_18),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_145),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_80),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_22),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_122),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_55),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_32),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_136),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_83),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_115),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_138),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_148),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_113),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_95),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_55),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_20),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_39),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_37),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_109),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_107),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_44),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_78),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_128),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_4),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_120),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_30),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_79),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_36),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_119),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_143),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_12),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_158),
.B(n_0),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_178),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_243),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_205),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_198),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_211),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_R g311 ( 
.A(n_250),
.B(n_212),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_216),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_228),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_231),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_159),
.B(n_2),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_192),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_258),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_241),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_161),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_244),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_192),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_192),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_245),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_192),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_227),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_227),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_253),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_213),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_227),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_254),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_256),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_230),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_166),
.B(n_182),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_152),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_152),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_195),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_197),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_239),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_213),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_239),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_167),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_174),
.B(n_6),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_150),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_199),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_270),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_166),
.B(n_8),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_150),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_198),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_284),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_153),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_200),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_167),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_284),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_298),
.B(n_198),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_353),
.B(n_174),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_309),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_162),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_309),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_320),
.B(n_170),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_182),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_299),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

CKINVDCx8_ASAP7_75t_R g387 ( 
.A(n_359),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_162),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_238),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_208),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_301),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_296),
.B1(n_189),
.B2(n_293),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_303),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_303),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_208),
.Y(n_399)
);

AND3x1_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_238),
.C(n_181),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_359),
.B(n_164),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_334),
.B(n_164),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_184),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_346),
.B(n_173),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_318),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_341),
.Y(n_420)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_184),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_352),
.A2(n_296),
.B1(n_293),
.B2(n_163),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_291),
.B1(n_206),
.B2(n_242),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_373),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_L g437 ( 
.A(n_374),
.B(n_304),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_368),
.B(n_310),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_367),
.B(n_364),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_399),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_391),
.B(n_188),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_368),
.B(n_312),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_391),
.A2(n_316),
.B1(n_236),
.B2(n_255),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_405),
.B(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_398),
.Y(n_458)
);

BUFx8_ASAP7_75t_SL g459 ( 
.A(n_392),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_377),
.B(n_314),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_374),
.B(n_322),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_372),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_388),
.B(n_324),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_378),
.B(n_328),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_402),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_401),
.B(n_357),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_394),
.A2(n_321),
.B1(n_313),
.B2(n_317),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_402),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_413),
.A2(n_302),
.B1(n_300),
.B2(n_305),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_400),
.B(n_188),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_415),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_399),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_421),
.B(n_332),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_388),
.B(n_336),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_421),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_367),
.B(n_345),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_337),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_382),
.B(n_267),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_378),
.B(n_344),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_376),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_382),
.B(n_267),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_422),
.B(n_354),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_365),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_316),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_387),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_363),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_392),
.B(n_362),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_422),
.B(n_361),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_365),
.Y(n_508)
);

NOR2x1p5_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_236),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_382),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_376),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_366),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_392),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_427),
.B(n_362),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_393),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_406),
.A2(n_154),
.B(n_151),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_366),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_369),
.B(n_160),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_398),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_398),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_427),
.A2(n_201),
.B1(n_234),
.B2(n_246),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_398),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_394),
.B(n_305),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_393),
.B(n_311),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_370),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_403),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_403),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_403),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_379),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_370),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_428),
.B(n_305),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_427),
.B(n_306),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_371),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_379),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_398),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_173),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_371),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_379),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_375),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_427),
.B(n_187),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_424),
.B(n_358),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_407),
.B(n_294),
.Y(n_549)
);

NOR2x1p5_ASAP7_75t_L g550 ( 
.A(n_387),
.B(n_161),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_379),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_375),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_425),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_426),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_425),
.B(n_235),
.C(n_240),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_380),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_407),
.B(n_155),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_423),
.B(n_177),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_380),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_407),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_426),
.B(n_177),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_420),
.B(n_156),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_384),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_420),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_407),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_407),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_385),
.B(n_179),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_385),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_410),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_445),
.B(n_410),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_516),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_514),
.B(n_179),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_485),
.B(n_183),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_445),
.B(n_410),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_438),
.A2(n_183),
.B1(n_219),
.B2(n_259),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_464),
.B(n_410),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_440),
.B(n_348),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_467),
.B(n_410),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_514),
.B(n_487),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_448),
.B(n_442),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_435),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_440),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_432),
.B(n_163),
.Y(n_589)
);

BUFx5_ASAP7_75t_L g590 ( 
.A(n_492),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_410),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_565),
.B(n_417),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_456),
.A2(n_259),
.B1(n_263),
.B2(n_266),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_453),
.B(n_229),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_535),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_436),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_490),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_442),
.B(n_219),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_553),
.B(n_263),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_459),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_528),
.B(n_417),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_439),
.B(n_417),
.Y(n_603)
);

NAND3xp33_ASAP7_75t_L g604 ( 
.A(n_553),
.B(n_209),
.C(n_226),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_436),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_441),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_442),
.B(n_266),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_439),
.B(n_506),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_503),
.A2(n_225),
.B1(n_157),
.B2(n_165),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_479),
.B(n_268),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_540),
.Y(n_611)
);

BUFx5_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

OAI221xp5_ASAP7_75t_L g613 ( 
.A1(n_454),
.A2(n_248),
.B1(n_224),
.B2(n_220),
.C(n_249),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_544),
.B(n_417),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_551),
.B(n_417),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_479),
.B(n_268),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_481),
.A2(n_261),
.B1(n_190),
.B2(n_214),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_449),
.B(n_390),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_496),
.B(n_269),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_559),
.B(n_395),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_479),
.B(n_229),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_554),
.B(n_564),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_554),
.B(n_564),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_548),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_532),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_441),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_560),
.B(n_395),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_463),
.B(n_269),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_560),
.B(n_396),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_554),
.B(n_272),
.Y(n_633)
);

INVx6_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_570),
.B(n_396),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_443),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_443),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_446),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_538),
.B(n_272),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_503),
.B(n_229),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_570),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_532),
.B(n_510),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_456),
.B(n_196),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_510),
.B(n_404),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_511),
.B(n_404),
.Y(n_646)
);

OAI221xp5_ASAP7_75t_L g647 ( 
.A1(n_524),
.A2(n_274),
.B1(n_276),
.B2(n_280),
.C(n_289),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_446),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_525),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_503),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_511),
.B(n_408),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_538),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_215),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_495),
.B(n_273),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_517),
.B(n_408),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_447),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_517),
.B(n_409),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_503),
.B(n_262),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_520),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_455),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_429),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_507),
.B(n_481),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_523),
.A2(n_191),
.B(n_218),
.C(n_221),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_523),
.B(n_409),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_481),
.B(n_278),
.Y(n_667)
);

NOR2x1p5_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_501),
.Y(n_668)
);

NOR2xp67_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_412),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_509),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_525),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_518),
.A2(n_172),
.B1(n_215),
.B2(n_251),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_456),
.A2(n_437),
.B1(n_509),
.B2(n_527),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_497),
.B(n_172),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_447),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_414),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_497),
.B(n_172),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_531),
.B(n_414),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_531),
.A2(n_176),
.B(n_203),
.C(n_223),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_429),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_SL g682 ( 
.A1(n_477),
.A2(n_171),
.B1(n_169),
.B2(n_175),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_471),
.B(n_416),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_533),
.B(n_416),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_533),
.A2(n_260),
.B(n_193),
.C(n_194),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_555),
.B(n_281),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_537),
.A2(n_286),
.B1(n_288),
.B2(n_292),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_534),
.B(n_423),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_534),
.B(n_423),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_505),
.B(n_288),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_431),
.B(n_247),
.C(n_233),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_492),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_455),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_486),
.B(n_60),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_518),
.B(n_423),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_518),
.B(n_423),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_450),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_569),
.B(n_423),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_491),
.B(n_423),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_468),
.B(n_202),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_515),
.B(n_542),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_562),
.B(n_204),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_519),
.B(n_210),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_492),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_465),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_460),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_529),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_520),
.B(n_262),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_536),
.B(n_290),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_550),
.B(n_295),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_450),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_547),
.B(n_207),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_539),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_525),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_539),
.B(n_172),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_547),
.B(n_217),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_543),
.B(n_172),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_470),
.B(n_252),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_547),
.B(n_543),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_550),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_546),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_583),
.A2(n_458),
.B(n_461),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_584),
.B(n_546),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_584),
.B(n_552),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_SL g727 ( 
.A1(n_600),
.A2(n_279),
.B1(n_168),
.B2(n_169),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_588),
.B(n_552),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_588),
.B(n_556),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_SL g730 ( 
.A(n_707),
.B(n_262),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_578),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_586),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_598),
.B(n_556),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_580),
.A2(n_458),
.B(n_461),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_700),
.A2(n_458),
.B(n_461),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_602),
.A2(n_561),
.B(n_444),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_571),
.A2(n_561),
.B(n_444),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_SL g738 ( 
.A(n_675),
.B(n_168),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_573),
.A2(n_483),
.B(n_433),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_598),
.B(n_433),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_581),
.B(n_558),
.Y(n_741)
);

NAND2x1_ASAP7_75t_L g742 ( 
.A(n_634),
.B(n_475),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_581),
.B(n_675),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_608),
.B(n_434),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_596),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_642),
.B(n_434),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_577),
.A2(n_444),
.B(n_472),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_703),
.A2(n_549),
.B(n_557),
.C(n_563),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_591),
.A2(n_444),
.B(n_472),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_674),
.B(n_521),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_652),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_594),
.B(n_563),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_696),
.A2(n_482),
.B(n_451),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_592),
.B(n_451),
.Y(n_754)
);

NOR2x1p5_ASAP7_75t_SL g755 ( 
.A(n_590),
.B(n_460),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_603),
.B(n_452),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_521),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_678),
.B(n_664),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_600),
.B(n_563),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_585),
.B(n_521),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_611),
.Y(n_761)
);

BUFx8_ASAP7_75t_L g762 ( 
.A(n_710),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_623),
.B(n_563),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_572),
.B(n_452),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_650),
.B(n_522),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_721),
.A2(n_492),
.B1(n_500),
.B2(n_566),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_697),
.A2(n_483),
.B(n_457),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_574),
.B(n_457),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_582),
.B(n_466),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_669),
.B(n_488),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_627),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_617),
.A2(n_484),
.B1(n_475),
.B2(n_498),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_699),
.A2(n_430),
.B(n_541),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_627),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_631),
.A2(n_498),
.B(n_484),
.C(n_475),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_661),
.A2(n_430),
.B(n_541),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_576),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_644),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_582),
.B(n_466),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_636),
.B(n_484),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_631),
.A2(n_498),
.B(n_512),
.C(n_478),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_661),
.A2(n_430),
.B(n_525),
.Y(n_782)
);

NOR2x2_ASAP7_75t_L g783 ( 
.A(n_712),
.B(n_171),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_541),
.B(n_512),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_617),
.A2(n_500),
.B1(n_492),
.B2(n_480),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_576),
.B(n_348),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_615),
.A2(n_541),
.B(n_512),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_640),
.B(n_473),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_643),
.A2(n_673),
.B(n_721),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_713),
.A2(n_541),
.B(n_488),
.Y(n_790)
);

AOI21xp33_ASAP7_75t_L g791 ( 
.A1(n_701),
.A2(n_189),
.B(n_287),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_673),
.A2(n_494),
.B(n_478),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_590),
.B(n_522),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_650),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_627),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_713),
.A2(n_488),
.B(n_567),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_473),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_619),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_621),
.A2(n_568),
.B(n_567),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_SL g800 ( 
.A1(n_667),
.A2(n_482),
.B(n_499),
.C(n_494),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_658),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_621),
.A2(n_568),
.B(n_567),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_627),
.Y(n_803)
);

OAI21xp33_ASAP7_75t_L g804 ( 
.A1(n_654),
.A2(n_285),
.B(n_282),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_670),
.A2(n_500),
.B1(n_526),
.B2(n_566),
.Y(n_805)
);

BUFx12f_ASAP7_75t_L g806 ( 
.A(n_712),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_626),
.B(n_628),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_701),
.A2(n_480),
.B(n_489),
.C(n_499),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_663),
.B(n_489),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_522),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_619),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_662),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_683),
.B(n_526),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_709),
.B(n_545),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_649),
.A2(n_568),
.B(n_567),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_715),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_689),
.A2(n_476),
.B(n_462),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_649),
.A2(n_568),
.B(n_567),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_590),
.B(n_500),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_723),
.B(n_545),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_690),
.A2(n_476),
.B(n_462),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_645),
.A2(n_651),
.B(n_646),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_587),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_671),
.A2(n_568),
.B(n_567),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_604),
.B(n_469),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_590),
.B(n_566),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_722),
.B(n_474),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_662),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_622),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_671),
.A2(n_716),
.B(n_595),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_595),
.B(n_545),
.Y(n_831)
);

NOR2x1p5_ASAP7_75t_SL g832 ( 
.A(n_590),
.B(n_493),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_630),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_655),
.A2(n_500),
.B(n_568),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_SL g835 ( 
.A(n_601),
.B(n_275),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_716),
.A2(n_500),
.B(n_358),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_654),
.A2(n_275),
.B(n_180),
.C(n_185),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_684),
.A2(n_500),
.B1(n_215),
.B2(n_265),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_702),
.A2(n_351),
.B(n_350),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_613),
.A2(n_351),
.B(n_350),
.C(n_215),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_632),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_657),
.A2(n_222),
.B(n_279),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_579),
.A2(n_282),
.B(n_277),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_666),
.A2(n_215),
.B(n_65),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_624),
.B(n_215),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_635),
.B(n_215),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_662),
.A2(n_277),
.B(n_265),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_681),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_692),
.A2(n_215),
.B1(n_222),
.B2(n_257),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_681),
.A2(n_257),
.B(n_186),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_712),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_644),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_625),
.B(n_186),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_641),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_597),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_618),
.B(n_185),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_722),
.B(n_705),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_634),
.Y(n_858)
);

BUFx8_ASAP7_75t_L g859 ( 
.A(n_659),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_714),
.A2(n_180),
.B(n_175),
.C(n_17),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_668),
.B(n_146),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_681),
.A2(n_129),
.B(n_125),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_714),
.A2(n_10),
.B(n_12),
.C(n_18),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_590),
.B(n_123),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_691),
.B(n_19),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_677),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_589),
.B(n_575),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_681),
.A2(n_118),
.B(n_116),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_644),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_698),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_SL g871 ( 
.A1(n_665),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_698),
.B(n_21),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_698),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_698),
.A2(n_110),
.B(n_104),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_679),
.A2(n_103),
.B(n_98),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_685),
.A2(n_91),
.B(n_90),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_694),
.A2(n_87),
.B(n_81),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_620),
.B(n_72),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_718),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_708),
.B(n_25),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_634),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_605),
.B(n_26),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_653),
.A2(n_62),
.B(n_27),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_606),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_629),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_637),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_638),
.A2(n_26),
.B(n_27),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_639),
.A2(n_28),
.B(n_31),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_648),
.A2(n_31),
.B(n_32),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_620),
.Y(n_890)
);

BUFx4f_ASAP7_75t_L g891 ( 
.A(n_656),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_599),
.B(n_607),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_676),
.B(n_33),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_704),
.A2(n_40),
.B(n_43),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_612),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_870),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_829),
.B(n_833),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_777),
.B(n_693),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_732),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_841),
.B(n_718),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_731),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_738),
.B(n_660),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_745),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_887),
.A2(n_889),
.B1(n_692),
.B2(n_758),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_777),
.B(n_693),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_866),
.B(n_633),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_819),
.A2(n_695),
.B(n_706),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_751),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_761),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_759),
.B(n_798),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_780),
.B(n_660),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_858),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_763),
.A2(n_720),
.B1(n_687),
.B2(n_610),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_806),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_741),
.A2(n_593),
.B(n_688),
.C(n_616),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_816),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_751),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_758),
.A2(n_711),
.B1(n_647),
.B2(n_682),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_786),
.B(n_706),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_807),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_798),
.A2(n_719),
.B1(n_717),
.B2(n_686),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_811),
.B(n_612),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_811),
.B(n_612),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_789),
.A2(n_680),
.B(n_612),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_823),
.Y(n_925)
);

INVxp67_ASAP7_75t_SL g926 ( 
.A(n_870),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_870),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_895),
.A2(n_612),
.B(n_693),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_864),
.A2(n_612),
.B(n_693),
.C(n_706),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_807),
.B(n_45),
.Y(n_930)
);

O2A1O1Ixp5_ASAP7_75t_SL g931 ( 
.A1(n_791),
.A2(n_50),
.B(n_52),
.C(n_693),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_743),
.B(n_693),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_794),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_853),
.A2(n_706),
.B(n_50),
.C(n_52),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_870),
.Y(n_935)
);

OAI22x1_ASAP7_75t_L g936 ( 
.A1(n_743),
.A2(n_706),
.B1(n_853),
.B2(n_857),
.Y(n_936)
);

O2A1O1Ixp5_ASAP7_75t_L g937 ( 
.A1(n_845),
.A2(n_706),
.B(n_750),
.C(n_788),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_725),
.A2(n_726),
.B1(n_757),
.B2(n_733),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_873),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_752),
.A2(n_857),
.B1(n_892),
.B2(n_878),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_895),
.A2(n_767),
.B(n_753),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_SL g942 ( 
.A(n_804),
.B(n_730),
.C(n_842),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_728),
.B(n_729),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_769),
.Y(n_944)
);

CKINVDCx11_ASAP7_75t_R g945 ( 
.A(n_851),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_SL g946 ( 
.A1(n_760),
.A2(n_757),
.B(n_875),
.C(n_876),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_797),
.B(n_740),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_890),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_739),
.A2(n_724),
.B(n_734),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_852),
.B(n_849),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_744),
.B(n_754),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_779),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_827),
.B(n_801),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_867),
.B(n_794),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_762),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_764),
.B(n_768),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_756),
.B(n_865),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_873),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_785),
.A2(n_750),
.B1(n_891),
.B2(n_881),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_835),
.B(n_762),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_765),
.B(n_760),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_890),
.B(n_856),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_825),
.A2(n_780),
.B1(n_778),
.B2(n_852),
.Y(n_963)
);

INVx6_ASAP7_75t_L g964 ( 
.A(n_881),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_SL g965 ( 
.A1(n_864),
.A2(n_775),
.B(n_781),
.C(n_879),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_854),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_747),
.A2(n_735),
.B(n_790),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_746),
.B(n_771),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_737),
.A2(n_749),
.B(n_773),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_771),
.B(n_837),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_885),
.B(n_886),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_873),
.B(n_774),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_855),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_872),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_884),
.B(n_812),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_812),
.B(n_828),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_SL g977 ( 
.A(n_873),
.B(n_774),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_843),
.B(n_727),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_774),
.B(n_803),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_809),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_860),
.A2(n_792),
.B(n_808),
.C(n_748),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_880),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_785),
.A2(n_891),
.B1(n_766),
.B2(n_805),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_854),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_774),
.A2(n_803),
.B1(n_795),
.B2(n_828),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_882),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_847),
.B(n_850),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_736),
.A2(n_776),
.B(n_782),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_803),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_748),
.A2(n_877),
.B(n_838),
.C(n_863),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_803),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_795),
.B(n_848),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_861),
.B(n_849),
.Y(n_994)
);

O2A1O1Ixp5_ASAP7_75t_L g995 ( 
.A1(n_834),
.A2(n_846),
.B(n_822),
.C(n_826),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_893),
.A2(n_871),
.B(n_800),
.C(n_840),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_810),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_793),
.A2(n_826),
.B(n_831),
.C(n_814),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_839),
.B(n_770),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_859),
.B(n_813),
.Y(n_1001)
);

CKINVDCx6p67_ASAP7_75t_R g1002 ( 
.A(n_820),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_772),
.B(n_830),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_793),
.A2(n_787),
.B(n_784),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_817),
.B(n_821),
.Y(n_1005)
);

OAI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_894),
.A2(n_888),
.B(n_840),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_742),
.B(n_836),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_796),
.A2(n_883),
.B1(n_874),
.B2(n_868),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_783),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_844),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_755),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_832),
.B(n_862),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_799),
.B(n_802),
.C(n_815),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_818),
.B(n_824),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_741),
.A2(n_584),
.B(n_438),
.C(n_448),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_777),
.B(n_584),
.Y(n_1016)
);

AO21x1_ASAP7_75t_L g1017 ( 
.A1(n_758),
.A2(n_750),
.B(n_664),
.Y(n_1017)
);

BUFx4f_ASAP7_75t_L g1018 ( 
.A(n_806),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_870),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_819),
.A2(n_895),
.B(n_583),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_819),
.A2(n_895),
.B(n_583),
.Y(n_1021)
);

INVx3_ASAP7_75t_SL g1022 ( 
.A(n_783),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_SL g1023 ( 
.A1(n_970),
.A2(n_996),
.B(n_959),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_901),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_945),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_924),
.A2(n_937),
.B(n_995),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_947),
.B(n_897),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_903),
.Y(n_1029)
);

AOI221x1_ASAP7_75t_L g1030 ( 
.A1(n_934),
.A2(n_936),
.B1(n_1006),
.B2(n_938),
.C(n_969),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_994),
.A2(n_1003),
.B(n_1008),
.C(n_1014),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_907),
.A2(n_1005),
.B(n_1021),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_SL g1033 ( 
.A1(n_983),
.A2(n_922),
.B(n_923),
.Y(n_1033)
);

NAND3x1_ASAP7_75t_L g1034 ( 
.A(n_1001),
.B(n_963),
.C(n_954),
.Y(n_1034)
);

AO32x2_ASAP7_75t_L g1035 ( 
.A1(n_918),
.A2(n_921),
.A3(n_985),
.B1(n_931),
.B2(n_965),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_957),
.B(n_956),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_909),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_1003),
.A2(n_1004),
.B(n_967),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_961),
.A2(n_932),
.B(n_1020),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_986),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_943),
.A2(n_919),
.B(n_989),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_1016),
.B(n_906),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_1014),
.A2(n_932),
.A3(n_1012),
.B(n_988),
.Y(n_1043)
);

CKINVDCx11_ASAP7_75t_R g1044 ( 
.A(n_955),
.Y(n_1044)
);

AO32x2_ASAP7_75t_L g1045 ( 
.A1(n_920),
.A2(n_950),
.A3(n_917),
.B1(n_912),
.B2(n_910),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_929),
.A2(n_999),
.B(n_928),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_950),
.A2(n_940),
.B1(n_962),
.B2(n_974),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_1013),
.A2(n_905),
.B(n_898),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_972),
.A2(n_1007),
.B(n_968),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_984),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1007),
.A2(n_898),
.B(n_905),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_980),
.A2(n_982),
.B(n_987),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_988),
.A2(n_1000),
.B(n_926),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_926),
.A2(n_935),
.B(n_939),
.Y(n_1054)
);

AO21x1_ASAP7_75t_L g1055 ( 
.A1(n_979),
.A2(n_913),
.B(n_998),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_944),
.B(n_952),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_962),
.B(n_974),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_966),
.Y(n_1058)
);

AO31x2_ASAP7_75t_L g1059 ( 
.A1(n_953),
.A2(n_975),
.A3(n_971),
.B(n_976),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1011),
.A2(n_954),
.B(n_916),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_SL g1061 ( 
.A(n_902),
.B(n_977),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_930),
.B(n_911),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_902),
.B(n_908),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_SL g1064 ( 
.A1(n_911),
.A2(n_992),
.B(n_908),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_964),
.A2(n_933),
.B1(n_925),
.B2(n_973),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_993),
.A2(n_1011),
.B(n_912),
.Y(n_1066)
);

AOI221x1_ASAP7_75t_L g1067 ( 
.A1(n_1001),
.A2(n_896),
.B1(n_1019),
.B2(n_990),
.C(n_927),
.Y(n_1067)
);

AOI221x1_ASAP7_75t_L g1068 ( 
.A1(n_896),
.A2(n_1019),
.B1(n_958),
.B2(n_927),
.C(n_990),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_899),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_933),
.A2(n_1022),
.B(n_948),
.C(n_1009),
.Y(n_1070)
);

AOI221x1_ASAP7_75t_L g1071 ( 
.A1(n_958),
.A2(n_990),
.B1(n_1002),
.B2(n_1022),
.C(n_960),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_964),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_964),
.A2(n_1018),
.B(n_997),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_1018),
.B(n_960),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_914),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_901),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1077)
);

AO32x2_ASAP7_75t_L g1078 ( 
.A1(n_938),
.A2(n_918),
.A3(n_959),
.B1(n_609),
.B2(n_983),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_901),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_964),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_908),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1015),
.A2(n_978),
.B1(n_738),
.B2(n_942),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_947),
.B(n_588),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_964),
.Y(n_1088)
);

CKINVDCx8_ASAP7_75t_R g1089 ( 
.A(n_984),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_948),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_901),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1093)
);

AO21x2_ASAP7_75t_L g1094 ( 
.A1(n_949),
.A2(n_946),
.B(n_941),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1015),
.A2(n_915),
.B(n_584),
.C(n_448),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_900),
.B(n_777),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_900),
.B(n_777),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_900),
.B(n_777),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_978),
.A2(n_942),
.B1(n_950),
.B2(n_791),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_908),
.Y(n_1101)
);

INVx3_ASAP7_75t_SL g1102 ( 
.A(n_984),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_994),
.A2(n_938),
.B(n_961),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1015),
.B(n_448),
.C(n_438),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1017),
.A2(n_970),
.B(n_889),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_947),
.B(n_588),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1015),
.A2(n_445),
.B1(n_904),
.B2(n_897),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_964),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_901),
.Y(n_1110)
);

AO21x1_ASAP7_75t_L g1111 ( 
.A1(n_994),
.A2(n_938),
.B(n_961),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1015),
.A2(n_915),
.B(n_791),
.C(n_942),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_1001),
.Y(n_1117)
);

OAI22x1_ASAP7_75t_L g1118 ( 
.A1(n_978),
.A2(n_940),
.B1(n_963),
.B2(n_743),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_977),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_908),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1122)
);

AOI221x1_ASAP7_75t_L g1123 ( 
.A1(n_1015),
.A2(n_934),
.B1(n_991),
.B2(n_936),
.C(n_1006),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_941),
.A2(n_991),
.B(n_981),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1015),
.A2(n_915),
.B(n_584),
.C(n_448),
.Y(n_1125)
);

BUFx8_ASAP7_75t_L g1126 ( 
.A(n_955),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_908),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_947),
.B(n_588),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1015),
.A2(n_915),
.B(n_584),
.C(n_448),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_945),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1015),
.B(n_448),
.C(n_438),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1015),
.A2(n_445),
.B1(n_904),
.B2(n_897),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_947),
.B(n_588),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_SL g1140 ( 
.A(n_959),
.B(n_858),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_941),
.A2(n_991),
.B(n_981),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1015),
.A2(n_981),
.B(n_991),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_948),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_967),
.A2(n_1004),
.B(n_989),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1015),
.A2(n_981),
.B(n_991),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1015),
.A2(n_981),
.B(n_991),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1017),
.A2(n_991),
.A3(n_981),
.B(n_1010),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_941),
.A2(n_949),
.B(n_951),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1099),
.A2(n_1133),
.B1(n_1104),
.B2(n_1142),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_1044),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_SL g1151 ( 
.A1(n_1104),
.A2(n_1133),
.B1(n_1137),
.B2(n_1107),
.Y(n_1151)
);

OAI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_1095),
.A2(n_1129),
.B(n_1125),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1028),
.B(n_1036),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1028),
.A2(n_1084),
.B1(n_1036),
.B2(n_1047),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1142),
.A2(n_1145),
.B1(n_1146),
.B2(n_1137),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1026),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1110),
.Y(n_1157)
);

INVx6_ASAP7_75t_L g1158 ( 
.A(n_1082),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1083),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1084),
.A2(n_1047),
.B1(n_1097),
.B2(n_1057),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_SL g1161 ( 
.A1(n_1107),
.A2(n_1145),
.B1(n_1146),
.B2(n_1124),
.Y(n_1161)
);

OAI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1087),
.A2(n_1106),
.B1(n_1128),
.B2(n_1139),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1090),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1034),
.A2(n_1118),
.B1(n_1042),
.B2(n_1063),
.Y(n_1164)
);

OAI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1087),
.A2(n_1106),
.B1(n_1128),
.B2(n_1139),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1024),
.Y(n_1166)
);

OAI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1056),
.A2(n_1123),
.B1(n_1071),
.B2(n_1052),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1089),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1082),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1124),
.A2(n_1141),
.B1(n_1023),
.B2(n_1096),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1103),
.A2(n_1111),
.B1(n_1141),
.B2(n_1098),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1037),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1076),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

BUFx8_ASAP7_75t_L g1175 ( 
.A(n_1130),
.Y(n_1175)
);

CKINVDCx11_ASAP7_75t_R g1176 ( 
.A(n_1058),
.Y(n_1176)
);

OAI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1065),
.A2(n_1143),
.B1(n_1060),
.B2(n_1101),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1088),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1081),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1113),
.A2(n_1119),
.B1(n_1127),
.B2(n_1121),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1092),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1105),
.A2(n_1033),
.B1(n_1039),
.B2(n_1094),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1069),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1102),
.Y(n_1184)
);

CKINVDCx11_ASAP7_75t_R g1185 ( 
.A(n_1050),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1117),
.Y(n_1186)
);

CKINVDCx11_ASAP7_75t_R g1187 ( 
.A(n_1075),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1059),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1060),
.B(n_1043),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1072),
.B(n_1061),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1059),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1059),
.Y(n_1192)
);

BUFx8_ASAP7_75t_SL g1193 ( 
.A(n_1074),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1075),
.A2(n_1109),
.B1(n_1117),
.B2(n_1070),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1039),
.A2(n_1094),
.B1(n_1055),
.B2(n_1148),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1045),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1073),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1140),
.A2(n_1078),
.B1(n_1027),
.B2(n_1126),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1048),
.B(n_1054),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1075),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_1126),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1043),
.B(n_1025),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1064),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1080),
.Y(n_1205)
);

CKINVDCx11_ASAP7_75t_R g1206 ( 
.A(n_1078),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1080),
.B(n_1086),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_1045),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1077),
.A2(n_1115),
.B1(n_1138),
.B2(n_1134),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1078),
.A2(n_1027),
.B1(n_1120),
.B2(n_1116),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1045),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1049),
.A2(n_1053),
.B1(n_1132),
.B2(n_1085),
.Y(n_1212)
);

CKINVDCx11_ASAP7_75t_R g1213 ( 
.A(n_1035),
.Y(n_1213)
);

BUFx4_ASAP7_75t_SL g1214 ( 
.A(n_1030),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1035),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1051),
.A2(n_1041),
.B1(n_1066),
.B2(n_1035),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1032),
.A2(n_1046),
.B1(n_1144),
.B2(n_1093),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1038),
.A2(n_1031),
.B1(n_1147),
.B2(n_1091),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1079),
.A2(n_1122),
.B1(n_1100),
.B2(n_1136),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1147),
.B(n_1091),
.Y(n_1220)
);

CKINVDCx6p67_ASAP7_75t_R g1221 ( 
.A(n_1108),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1112),
.A2(n_1135),
.B1(n_1114),
.B2(n_1131),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1112),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1135),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_1133),
.B2(n_942),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1040),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_1133),
.B2(n_942),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1044),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1036),
.B(n_1028),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1088),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1095),
.A2(n_1015),
.B(n_1125),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1062),
.B(n_911),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1029),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_SL g1234 ( 
.A(n_1026),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1040),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_1133),
.B2(n_942),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1083),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1082),
.B(n_977),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1087),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1029),
.Y(n_1240)
);

BUFx2_ASAP7_75t_SL g1241 ( 
.A(n_1040),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1099),
.A2(n_1104),
.B1(n_1133),
.B2(n_942),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1104),
.A2(n_738),
.B1(n_950),
.B2(n_1133),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1082),
.B(n_977),
.Y(n_1244)
);

CKINVDCx6p67_ASAP7_75t_R g1245 ( 
.A(n_1058),
.Y(n_1245)
);

AOI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_1133),
.B(n_1113),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1089),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1104),
.A2(n_738),
.B1(n_950),
.B2(n_1133),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1104),
.A2(n_738),
.B1(n_950),
.B2(n_1133),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1104),
.A2(n_738),
.B1(n_950),
.B2(n_1133),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1040),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1082),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1189),
.B(n_1211),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1199),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1217),
.A2(n_1219),
.B(n_1200),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1188),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1159),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1166),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1158),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1237),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1206),
.B(n_1151),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1246),
.A2(n_1216),
.B(n_1218),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1191),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1192),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1223),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1208),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1195),
.A2(n_1209),
.B(n_1203),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1163),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1229),
.B(n_1153),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1217),
.A2(n_1219),
.B(n_1200),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1202),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1205),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1207),
.B(n_1196),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1160),
.B(n_1154),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1220),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1180),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1208),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1216),
.A2(n_1218),
.B(n_1212),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1158),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1225),
.A2(n_1242),
.B(n_1236),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1222),
.A2(n_1209),
.B(n_1195),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1204),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1224),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1168),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1224),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1239),
.B(n_1155),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1221),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1155),
.B(n_1149),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1204),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1172),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1241),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1173),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1179),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1181),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_1186),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1164),
.B(n_1157),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1214),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1158),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1214),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1151),
.B(n_1149),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1190),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1183),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1161),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1161),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1233),
.B(n_1227),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1182),
.A2(n_1231),
.B(n_1152),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1225),
.A2(n_1227),
.B(n_1242),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1210),
.A2(n_1213),
.A3(n_1215),
.B(n_1182),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1240),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1183),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1162),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1162),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1198),
.B(n_1250),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1198),
.B(n_1250),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1194),
.B(n_1238),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1165),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1236),
.B(n_1171),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1177),
.A2(n_1197),
.B1(n_1243),
.B2(n_1249),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1171),
.B(n_1210),
.Y(n_1320)
);

AO21x1_ASAP7_75t_SL g1321 ( 
.A1(n_1167),
.A2(n_1243),
.B(n_1249),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1248),
.B(n_1170),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1183),
.Y(n_1323)
);

AOI222xp33_ASAP7_75t_L g1324 ( 
.A1(n_1234),
.A2(n_1175),
.B1(n_1167),
.B2(n_1228),
.C1(n_1150),
.C2(n_1176),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1248),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1232),
.A2(n_1245),
.B1(n_1234),
.B2(n_1178),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1247),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1230),
.B(n_1232),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1280),
.A2(n_1307),
.B(n_1274),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1254),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1322),
.B(n_1201),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1322),
.B(n_1244),
.Y(n_1332)
);

NAND4xp25_ASAP7_75t_SL g1333 ( 
.A(n_1324),
.B(n_1202),
.C(n_1187),
.D(n_1193),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1303),
.B(n_1251),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1290),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1273),
.B(n_1253),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1304),
.B(n_1235),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1281),
.A2(n_1156),
.B(n_1169),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1306),
.A2(n_1169),
.B(n_1252),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1281),
.A2(n_1174),
.B(n_1226),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1304),
.B(n_1174),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1319),
.B(n_1226),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1300),
.A2(n_1184),
.B(n_1175),
.C(n_1226),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1300),
.B(n_1185),
.C(n_1288),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1293),
.B(n_1308),
.Y(n_1345)
);

AO32x2_ASAP7_75t_L g1346 ( 
.A1(n_1273),
.A2(n_1253),
.A3(n_1308),
.B1(n_1262),
.B2(n_1298),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1261),
.A2(n_1313),
.B(n_1315),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1255),
.A2(n_1270),
.B(n_1265),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1308),
.B(n_1294),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1289),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1308),
.B(n_1294),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1256),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1288),
.A2(n_1261),
.B(n_1318),
.C(n_1315),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1263),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1318),
.A2(n_1296),
.B(n_1305),
.C(n_1325),
.Y(n_1355)
);

OAI211xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1291),
.A2(n_1269),
.B(n_1325),
.C(n_1326),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1263),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1268),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1297),
.A2(n_1299),
.B1(n_1316),
.B2(n_1295),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1308),
.B(n_1258),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1257),
.B(n_1260),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1264),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1270),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1297),
.A2(n_1299),
.B1(n_1316),
.B2(n_1295),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1276),
.A2(n_1311),
.B(n_1317),
.Y(n_1366)
);

NAND2x1_ASAP7_75t_L g1367 ( 
.A(n_1287),
.B(n_1283),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1292),
.B(n_1278),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1311),
.A2(n_1314),
.B1(n_1312),
.B2(n_1317),
.C(n_1313),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1271),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1278),
.A2(n_1267),
.B(n_1262),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1267),
.A2(n_1262),
.B(n_1320),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1320),
.B(n_1301),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1312),
.A2(n_1314),
.B(n_1286),
.C(n_1282),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1275),
.B(n_1267),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1352),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1345),
.B(n_1267),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1375),
.B(n_1275),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1342),
.A2(n_1321),
.B1(n_1286),
.B2(n_1266),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1340),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1364),
.B(n_1285),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1368),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1375),
.B(n_1264),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1345),
.B(n_1360),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1330),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1330),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1372),
.B(n_1354),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1354),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1357),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1340),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1329),
.B(n_1316),
.C(n_1309),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1340),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1363),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1336),
.B(n_1265),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1348),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1346),
.B(n_1272),
.Y(n_1397)
);

AND2x4_ASAP7_75t_SL g1398 ( 
.A(n_1385),
.B(n_1350),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1384),
.B(n_1346),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1388),
.B(n_1371),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1389),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1389),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1384),
.B(n_1346),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_1388),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1335),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1379),
.A2(n_1329),
.B1(n_1353),
.B2(n_1344),
.C(n_1355),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1391),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1396),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1379),
.A2(n_1347),
.B1(n_1369),
.B2(n_1356),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1396),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1381),
.B(n_1364),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1390),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1384),
.B(n_1387),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1390),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1394),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1392),
.A2(n_1347),
.B1(n_1333),
.B2(n_1366),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1387),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1394),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1376),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1392),
.A2(n_1343),
.B1(n_1374),
.B2(n_1359),
.C(n_1365),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1392),
.A2(n_1277),
.B1(n_1266),
.B2(n_1337),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1391),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1377),
.B(n_1373),
.Y(n_1423)
);

NOR2x1_ASAP7_75t_L g1424 ( 
.A(n_1391),
.B(n_1367),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1391),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1377),
.B(n_1373),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_1364),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_L g1428 ( 
.A(n_1388),
.B(n_1339),
.C(n_1289),
.Y(n_1428)
);

OAI31xp33_ASAP7_75t_L g1429 ( 
.A1(n_1385),
.A2(n_1277),
.A3(n_1332),
.B(n_1331),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1419),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1398),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1404),
.B(n_1383),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1399),
.B(n_1377),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1404),
.B(n_1383),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1419),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1400),
.B(n_1395),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1401),
.B(n_1395),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1408),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1401),
.B(n_1395),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.B(n_1386),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1399),
.B(n_1397),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1414),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1414),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1408),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1399),
.B(n_1397),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1408),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1424),
.B(n_1391),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1412),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1424),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1408),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1402),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_L g1453 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1411),
.B(n_1380),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1403),
.B(n_1393),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1412),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1402),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1415),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1407),
.B(n_1338),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1406),
.B(n_1370),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1418),
.B(n_1382),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1438),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1430),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1436),
.B(n_1416),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1436),
.B(n_1416),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1450),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1463),
.B(n_1370),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1431),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1440),
.B(n_1432),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1432),
.B(n_1423),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1430),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1435),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_1405),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1431),
.A2(n_1406),
.B1(n_1409),
.B2(n_1420),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1479)
);

NOR2x1_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1420),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1434),
.B(n_1423),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1448),
.A2(n_1409),
.B1(n_1428),
.B2(n_1421),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1452),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1435),
.Y(n_1484)
);

NAND2x1_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1407),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1449),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1448),
.A2(n_1428),
.B(n_1429),
.C(n_1421),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1459),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1433),
.B(n_1413),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1444),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1444),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1448),
.B(n_1417),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1434),
.B(n_1405),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1437),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1449),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1448),
.A2(n_1332),
.B1(n_1411),
.B2(n_1341),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1441),
.B(n_1417),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1437),
.A2(n_1411),
.B1(n_1341),
.B2(n_1334),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1456),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1441),
.B(n_1417),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1439),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1439),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1441),
.B(n_1427),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1471),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1476),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1426),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1473),
.B(n_1457),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1486),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1499),
.B(n_1445),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1482),
.B(n_1429),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1483),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1489),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1486),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1445),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1502),
.B(n_1445),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1497),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1457),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1502),
.B(n_1454),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1470),
.B(n_1284),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1506),
.B(n_1447),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1479),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1497),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1501),
.Y(n_1529)
);

BUFx2_ASAP7_75t_SL g1530 ( 
.A(n_1469),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1426),
.Y(n_1531)
);

INVx3_ASAP7_75t_SL g1532 ( 
.A(n_1504),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_SL g1533 ( 
.A(n_1487),
.B(n_1350),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1479),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1501),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1506),
.B(n_1447),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1504),
.B(n_1462),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1485),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1447),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1466),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1475),
.Y(n_1541)
);

NAND2x1_ASAP7_75t_SL g1542 ( 
.A(n_1532),
.B(n_1443),
.Y(n_1542)
);

OAI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1533),
.A2(n_1485),
.B1(n_1503),
.B2(n_1498),
.C(n_1469),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1508),
.B(n_1516),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1532),
.B(n_1495),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1515),
.A2(n_1524),
.B(n_1517),
.Y(n_1546)
);

OAI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1511),
.A2(n_1453),
.B(n_1500),
.C(n_1422),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1530),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1507),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1507),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

NOR3xp33_ASAP7_75t_L g1552 ( 
.A(n_1538),
.B(n_1505),
.C(n_1358),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1474),
.Y(n_1553)
);

CKINVDCx14_ASAP7_75t_R g1554 ( 
.A(n_1525),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

AOI211xp5_ASAP7_75t_L g1556 ( 
.A1(n_1532),
.A2(n_1453),
.B(n_1454),
.C(n_1494),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1530),
.Y(n_1558)
);

AND2x4_ASAP7_75t_SL g1559 ( 
.A(n_1523),
.B(n_1443),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1488),
.Y(n_1560)
);

OAI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1527),
.A2(n_1495),
.B1(n_1477),
.B2(n_1461),
.C(n_1481),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1477),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1513),
.Y(n_1563)
);

AOI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1512),
.A2(n_1522),
.B(n_1537),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1518),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1518),
.Y(n_1566)
);

AOI322xp5_ASAP7_75t_L g1567 ( 
.A1(n_1544),
.A2(n_1455),
.A3(n_1526),
.B1(n_1536),
.B2(n_1539),
.C1(n_1514),
.C2(n_1520),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1554),
.B(n_1526),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1565),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1565),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1543),
.A2(n_1534),
.B1(n_1527),
.B2(n_1536),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1549),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1542),
.A2(n_1546),
.B(n_1548),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1558),
.B(n_1534),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1559),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1540),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1554),
.A2(n_1541),
.B(n_1522),
.Y(n_1577)
);

OAI322xp33_ASAP7_75t_L g1578 ( 
.A1(n_1545),
.A2(n_1541),
.A3(n_1512),
.B1(n_1535),
.B2(n_1521),
.C1(n_1529),
.C2(n_1528),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1550),
.Y(n_1579)
);

OAI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1547),
.A2(n_1537),
.B1(n_1531),
.B2(n_1535),
.C(n_1529),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1521),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_1514),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1519),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1564),
.B(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1559),
.Y(n_1585)
);

AOI31xp33_ASAP7_75t_L g1586 ( 
.A1(n_1573),
.A2(n_1556),
.A3(n_1563),
.B(n_1557),
.Y(n_1586)
);

OAI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1584),
.A2(n_1561),
.B1(n_1553),
.B2(n_1562),
.C(n_1555),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1568),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1584),
.A2(n_1566),
.B(n_1551),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1577),
.B(n_1472),
.C(n_1465),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1569),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1575),
.Y(n_1592)
);

AOI32xp33_ASAP7_75t_L g1593 ( 
.A1(n_1585),
.A2(n_1520),
.A3(n_1519),
.B1(n_1523),
.B2(n_1407),
.Y(n_1593)
);

AOI211xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1578),
.A2(n_1523),
.B(n_1460),
.C(n_1484),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1575),
.B(n_1488),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1588),
.B(n_1581),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1595),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1574),
.Y(n_1598)
);

AOI221x1_ASAP7_75t_L g1599 ( 
.A1(n_1591),
.A2(n_1570),
.B1(n_1572),
.B2(n_1579),
.C(n_1571),
.Y(n_1599)
);

AOI21xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1586),
.A2(n_1581),
.B(n_1576),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1594),
.B(n_1593),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1586),
.B(n_1567),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_L g1603 ( 
.A(n_1590),
.B(n_1580),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1589),
.B(n_1583),
.C(n_1582),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1600),
.B(n_1587),
.Y(n_1605)
);

AOI31xp33_ASAP7_75t_L g1606 ( 
.A1(n_1596),
.A2(n_1302),
.A3(n_1323),
.B(n_1310),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1597),
.B(n_1490),
.Y(n_1607)
);

AOI211xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1603),
.A2(n_1460),
.B(n_1442),
.C(n_1491),
.Y(n_1608)
);

OAI211xp5_ASAP7_75t_L g1609 ( 
.A1(n_1602),
.A2(n_1425),
.B(n_1422),
.C(n_1323),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1605),
.A2(n_1601),
.B(n_1598),
.C(n_1604),
.Y(n_1610)
);

AOI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_1599),
.B(n_1362),
.C(n_1310),
.Y(n_1611)
);

NAND4xp75_ASAP7_75t_L g1612 ( 
.A(n_1607),
.B(n_1442),
.C(n_1492),
.D(n_1491),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1608),
.B(n_1490),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1606),
.A2(n_1425),
.B(n_1422),
.C(n_1361),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1608),
.A2(n_1425),
.B1(n_1461),
.B2(n_1472),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1613),
.Y(n_1616)
);

XNOR2xp5_ASAP7_75t_L g1617 ( 
.A(n_1611),
.B(n_1334),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1612),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1615),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1610),
.B(n_1614),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1616),
.Y(n_1621)
);

AOI221x1_ASAP7_75t_L g1622 ( 
.A1(n_1618),
.A2(n_1493),
.B1(n_1492),
.B2(n_1465),
.C(n_1462),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_SL g1623 ( 
.A(n_1616),
.B(n_1461),
.C(n_1493),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1621),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1620),
.B1(n_1619),
.B2(n_1623),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_1617),
.B1(n_1622),
.B2(n_1455),
.Y(n_1626)
);

XNOR2x1_ASAP7_75t_L g1627 ( 
.A(n_1626),
.B(n_1337),
.Y(n_1627)
);

XNOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1627),
.B(n_1331),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1628),
.A2(n_1446),
.B(n_1444),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1629),
.A2(n_1446),
.B(n_1451),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1629),
.A2(n_1446),
.B(n_1451),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1630),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1631),
.Y(n_1633)
);

OAI221xp5_ASAP7_75t_R g1634 ( 
.A1(n_1633),
.A2(n_1461),
.B1(n_1451),
.B2(n_1458),
.C(n_1455),
.Y(n_1634)
);

AOI211xp5_ASAP7_75t_L g1635 ( 
.A1(n_1634),
.A2(n_1632),
.B(n_1279),
.C(n_1259),
.Y(n_1635)
);


endmodule