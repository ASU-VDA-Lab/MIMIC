module fake_ariane_2274_n_974 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_974);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_974;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_307;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_269;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_485;
wire n_401;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_840;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_689;
wire n_694;
wire n_400;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_260;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_262;
wire n_490;
wire n_743;
wire n_907;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_527;
wire n_290;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_609;
wire n_444;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_437;
wire n_697;
wire n_622;
wire n_274;
wire n_337;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_548;
wire n_542;
wire n_289;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_114),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_58),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_10),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_158),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_90),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_132),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_111),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_83),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_49),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_118),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_112),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_215),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_124),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_13),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_59),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_110),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_161),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_174),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_98),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_187),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_146),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_44),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_122),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_96),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_84),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_2),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_186),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_137),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_24),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_200),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_103),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_82),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_144),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_80),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_169),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_176),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_172),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_177),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_97),
.B(n_232),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_117),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_104),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_15),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_30),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_107),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_120),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_35),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_123),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_69),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_224),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_142),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_23),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_133),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_147),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_99),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_31),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_57),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_67),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_206),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_113),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_210),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_18),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_164),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_101),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_63),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_139),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_213),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_196),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_173),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_106),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_226),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_8),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_8),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_79),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_85),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_119),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_30),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_17),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_195),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_189),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_135),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_153),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_18),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_38),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_205),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_170),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_68),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_13),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_72),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_163),
.B(n_179),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_55),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_33),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_102),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_28),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_130),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_86),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_56),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_236),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_115),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_191),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_9),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_175),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_109),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_227),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_218),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_0),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_121),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_100),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_145),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_127),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_81),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_220),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_43),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_39),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_216),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_125),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_162),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_152),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_52),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_211),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_105),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_75),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_204),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_9),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_47),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_292),
.B(n_0),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_315),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

OAI22x1_ASAP7_75t_R g412 ( 
.A1(n_240),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_238),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_292),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_309),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_315),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_296),
.B(n_1),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_298),
.B(n_3),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_296),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_330),
.B(n_4),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_242),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_4),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_387),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_243),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_245),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_273),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_256),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_288),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_241),
.B(n_14),
.Y(n_431)
);

CKINVDCx11_ASAP7_75t_R g432 ( 
.A(n_379),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_280),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g434 ( 
.A(n_299),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_324),
.B(n_20),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_318),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_262),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_284),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_328),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_300),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_340),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

BUFx12f_ASAP7_75t_L g446 ( 
.A(n_272),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_287),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_21),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_364),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_355),
.B(n_22),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_346),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_346),
.B(n_45),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_376),
.B(n_22),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_244),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_247),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_283),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_251),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_254),
.B(n_24),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_257),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_258),
.Y(n_466)
);

BUFx12f_ASAP7_75t_L g467 ( 
.A(n_281),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_259),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_314),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_285),
.B(n_25),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_294),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_263),
.A2(n_26),
.B(n_29),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_266),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_305),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_335),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_329),
.Y(n_476)
);

OA21x2_ASAP7_75t_L g477 ( 
.A1(n_268),
.A2(n_31),
.B(n_32),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_332),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_347),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_271),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_275),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_286),
.B(n_34),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_291),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_352),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_353),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_338),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_293),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_297),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_360),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_365),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_302),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_303),
.B(n_36),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_306),
.B(n_36),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_357),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_317),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_320),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_277),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_323),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_310),
.B(n_37),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_370),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_325),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_326),
.B(n_37),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_336),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_343),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_319),
.B(n_40),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_237),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_350),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_356),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_358),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_351),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_363),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_362),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_367),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_374),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_380),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_333),
.B(n_41),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_316),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_377),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_349),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_381),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_383),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_361),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_386),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_378),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_392),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_373),
.A2(n_48),
.B(n_46),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_395),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_403),
.B(n_51),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_239),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_316),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_385),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_246),
.Y(n_534)
);

BUFx8_ASAP7_75t_SL g535 ( 
.A(n_389),
.Y(n_535)
);

XNOR2x2_ASAP7_75t_L g536 ( 
.A(n_253),
.B(n_42),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_535),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_413),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_439),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_438),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_447),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_393),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_R g546 ( 
.A(n_421),
.B(n_248),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_421),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_406),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_510),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_476),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_486),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_512),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_506),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_432),
.Y(n_557)
);

BUFx6f_ASAP7_75t_SL g558 ( 
.A(n_420),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_524),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_533),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_427),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_518),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_469),
.B(n_391),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_446),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_467),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_489),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_442),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_518),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_R g571 ( 
.A(n_475),
.B(n_249),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_534),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_R g577 ( 
.A(n_485),
.B(n_250),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_534),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_530),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_R g580 ( 
.A(n_500),
.B(n_252),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_R g581 ( 
.A(n_409),
.B(n_255),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_440),
.Y(n_582)
);

AND3x2_ASAP7_75t_L g583 ( 
.A(n_453),
.B(n_393),
.C(n_368),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_484),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_415),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_415),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g589 ( 
.A(n_416),
.B(n_402),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

AND3x2_ASAP7_75t_L g591 ( 
.A(n_459),
.B(n_368),
.C(n_311),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_437),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_490),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_R g594 ( 
.A(n_532),
.B(n_508),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_462),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_441),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_419),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_462),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_496),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_498),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_523),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_521),
.B(n_260),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_474),
.Y(n_603)
);

AND3x2_ASAP7_75t_L g604 ( 
.A(n_408),
.B(n_304),
.C(n_279),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_452),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_414),
.B(n_313),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_494),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_448),
.Y(n_608)
);

NOR2xp67_ASAP7_75t_L g609 ( 
.A(n_494),
.B(n_261),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_461),
.B(n_264),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_449),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_543),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_544),
.B(n_408),
.C(n_420),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_610),
.B(n_422),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_593),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_610),
.B(n_422),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_547),
.B(n_433),
.C(n_423),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_546),
.B(n_414),
.C(n_418),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_470),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_600),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_470),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_601),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_558),
.B(n_461),
.Y(n_625)
);

AO221x1_ASAP7_75t_L g626 ( 
.A1(n_597),
.A2(n_412),
.B1(n_425),
.B2(n_536),
.C(n_471),
.Y(n_626)
);

AO221x1_ASAP7_75t_L g627 ( 
.A1(n_574),
.A2(n_455),
.B1(n_451),
.B2(n_466),
.C(n_465),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_575),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_558),
.B(n_463),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_590),
.B(n_417),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_561),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_539),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_540),
.A2(n_499),
.B1(n_505),
.B2(n_516),
.Y(n_633)
);

AND2x4_ASAP7_75t_SL g634 ( 
.A(n_595),
.B(n_499),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_602),
.B(n_572),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_594),
.B(n_582),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_SL g637 ( 
.A(n_585),
.B(n_478),
.C(n_428),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_596),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_578),
.B(n_505),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_608),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_592),
.B(n_463),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_546),
.B(n_464),
.C(n_431),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_571),
.B(n_435),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_604),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_577),
.B(n_482),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_573),
.Y(n_648)
);

BUFx8_ASAP7_75t_L g649 ( 
.A(n_557),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_549),
.Y(n_650)
);

BUFx5_ASAP7_75t_L g651 ( 
.A(n_609),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_586),
.B(n_480),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_580),
.B(n_497),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_583),
.B(n_497),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_581),
.B(n_492),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_591),
.B(n_519),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_588),
.B(n_519),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_581),
.B(n_493),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_589),
.B(n_502),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_559),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_605),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_603),
.B(n_522),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_560),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_569),
.B(n_426),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_564),
.B(n_487),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_607),
.B(n_522),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_598),
.B(n_488),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_556),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_556),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_537),
.B(n_434),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_551),
.B(n_495),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_538),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_650),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_673),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_674),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_615),
.B(n_541),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_631),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_643),
.A2(n_611),
.B1(n_531),
.B2(n_483),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_662),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_612),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_620),
.A2(n_503),
.B1(n_504),
.B2(n_460),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_665),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_675),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_666),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_630),
.B(n_542),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_639),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_624),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_634),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_637),
.A2(n_511),
.B1(n_513),
.B2(n_509),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_616),
.Y(n_695)
);

BUFx8_ASAP7_75t_L g696 ( 
.A(n_645),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_642),
.B(n_495),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_649),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_619),
.A2(n_527),
.B1(n_515),
.B2(n_468),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_673),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_622),
.B(n_570),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_623),
.B(n_621),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_652),
.B(n_555),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_614),
.B(n_550),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_636),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_618),
.B(n_553),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_638),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_625),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_613),
.B(n_507),
.Y(n_710)
);

AO22x1_ASAP7_75t_L g711 ( 
.A1(n_629),
.A2(n_565),
.B1(n_567),
.B2(n_566),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_639),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_646),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_628),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_654),
.B(n_514),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_635),
.B(n_554),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_646),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_644),
.B(n_563),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_632),
.B(n_633),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_667),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_SL g721 ( 
.A1(n_626),
.A2(n_472),
.B1(n_477),
.B2(n_454),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_656),
.B(n_514),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_641),
.B(n_520),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_647),
.A2(n_658),
.B1(n_655),
.B2(n_661),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_669),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_646),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_640),
.B(n_468),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_SL g728 ( 
.A(n_670),
.B(n_267),
.C(n_265),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_617),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_627),
.A2(n_481),
.B1(n_491),
.B2(n_473),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_671),
.A2(n_411),
.B(n_410),
.C(n_472),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_672),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_653),
.B(n_481),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_648),
.B(n_552),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_651),
.B(n_491),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_660),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_663),
.Y(n_738)
);

AND2x6_ASAP7_75t_L g739 ( 
.A(n_657),
.B(n_382),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_680),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_676),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_SL g742 ( 
.A1(n_685),
.A2(n_397),
.B(n_668),
.C(n_664),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_702),
.A2(n_411),
.B(n_410),
.C(n_477),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_724),
.A2(n_526),
.B(n_525),
.C(n_501),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_679),
.B(n_525),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_697),
.A2(n_270),
.B(n_269),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_701),
.A2(n_528),
.B(n_274),
.C(n_276),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_706),
.B(n_528),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_714),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_695),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_710),
.A2(n_707),
.B(n_704),
.C(n_719),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_687),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_718),
.B(n_278),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_692),
.A2(n_684),
.B(n_703),
.C(n_723),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_690),
.A2(n_529),
.B(n_289),
.C(n_290),
.Y(n_755)
);

CKINVDCx11_ASAP7_75t_R g756 ( 
.A(n_688),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_282),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_736),
.A2(n_301),
.B(n_295),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_689),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_709),
.B(n_307),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_677),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_722),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_725),
.A2(n_458),
.B(n_401),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_693),
.B(n_308),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_720),
.B(n_312),
.Y(n_765)
);

CKINVDCx8_ASAP7_75t_R g766 ( 
.A(n_698),
.Y(n_766)
);

BUFx12f_ASAP7_75t_L g767 ( 
.A(n_696),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_734),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_708),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_694),
.B(n_321),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_716),
.B(n_715),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_699),
.B(n_327),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_731),
.A2(n_337),
.B(n_334),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_730),
.B(n_341),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_681),
.A2(n_344),
.B(n_342),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_683),
.B(n_345),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_680),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_700),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_729),
.A2(n_401),
.B(n_322),
.C(n_54),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_732),
.B(n_354),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_SL g782 ( 
.A(n_721),
.B(n_369),
.C(n_366),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_728),
.A2(n_400),
.B(n_371),
.C(n_375),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_682),
.A2(n_396),
.B(n_390),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_686),
.B(n_399),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_749),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_740),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_750),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_772),
.B(n_711),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_744),
.A2(n_733),
.B(n_738),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_763),
.A2(n_713),
.B(n_682),
.Y(n_791)
);

AO21x2_ASAP7_75t_L g792 ( 
.A1(n_743),
.A2(n_737),
.B(n_717),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_740),
.Y(n_793)
);

OAI21x1_ASAP7_75t_L g794 ( 
.A1(n_774),
.A2(n_717),
.B(n_713),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_781),
.A2(n_735),
.B(n_691),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_751),
.A2(n_712),
.B(n_726),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_757),
.A2(n_691),
.B(n_680),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_780),
.A2(n_705),
.B(n_691),
.Y(n_798)
);

BUFx8_ASAP7_75t_L g799 ( 
.A(n_767),
.Y(n_799)
);

AO21x1_ASAP7_75t_L g800 ( 
.A1(n_753),
.A2(n_739),
.B(n_401),
.Y(n_800)
);

BUFx12f_ASAP7_75t_L g801 ( 
.A(n_756),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_761),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_759),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_745),
.B(n_739),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_740),
.B(n_778),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_769),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_782),
.A2(n_705),
.B(n_739),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_778),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_779),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_771),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_785),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_752),
.B(n_705),
.Y(n_813)
);

AO21x2_ASAP7_75t_L g814 ( 
.A1(n_747),
.A2(n_401),
.B(n_322),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_748),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_741),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_777),
.B(n_322),
.Y(n_817)
);

INVx6_ASAP7_75t_L g818 ( 
.A(n_762),
.Y(n_818)
);

AO21x2_ASAP7_75t_L g819 ( 
.A1(n_742),
.A2(n_401),
.B(n_322),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_754),
.Y(n_820)
);

OA21x2_ASAP7_75t_L g821 ( 
.A1(n_783),
.A2(n_456),
.B(n_444),
.Y(n_821)
);

AO21x2_ASAP7_75t_L g822 ( 
.A1(n_746),
.A2(n_457),
.B(n_456),
.Y(n_822)
);

OA21x2_ASAP7_75t_L g823 ( 
.A1(n_770),
.A2(n_457),
.B(n_444),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_766),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_773),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_760),
.B(n_430),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_764),
.B(n_64),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_776),
.A2(n_784),
.B(n_755),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_775),
.B(n_430),
.Y(n_829)
);

INVx11_ASAP7_75t_L g830 ( 
.A(n_799),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_789),
.A2(n_817),
.B1(n_765),
.B2(n_813),
.Y(n_831)
);

BUFx8_ASAP7_75t_L g832 ( 
.A(n_801),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_793),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_807),
.Y(n_835)
);

OR2x6_ASAP7_75t_L g836 ( 
.A(n_818),
.B(n_758),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_804),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_786),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_800),
.A2(n_797),
.B(n_821),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_803),
.B(n_65),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_811),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_802),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_816),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_812),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_815),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_793),
.B(n_78),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_825),
.A2(n_820),
.B1(n_827),
.B2(n_805),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_796),
.B(n_87),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_787),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_827),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_792),
.A2(n_93),
.B(n_94),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_787),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_791),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_802),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_793),
.B(n_228),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_795),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_790),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_806),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_801),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_809),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_824),
.B(n_116),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_837),
.Y(n_863)
);

CKINVDCx12_ASAP7_75t_R g864 ( 
.A(n_830),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_847),
.B(n_808),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_R g866 ( 
.A(n_848),
.B(n_821),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_855),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_833),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_849),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_841),
.B(n_810),
.Y(n_870)
);

AO31x2_ASAP7_75t_L g871 ( 
.A1(n_858),
.A2(n_797),
.A3(n_826),
.B(n_823),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_860),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_853),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_SL g874 ( 
.A1(n_831),
.A2(n_829),
.B(n_828),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_834),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_854),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_847),
.B(n_823),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_840),
.B(n_829),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_832),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_856),
.B(n_794),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_856),
.B(n_819),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_842),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_838),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_853),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_857),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_862),
.B(n_814),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_845),
.B(n_814),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_859),
.B(n_798),
.Y(n_888)
);

AOI21xp33_ASAP7_75t_L g889 ( 
.A1(n_848),
.A2(n_823),
.B(n_822),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_835),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_890),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_863),
.B(n_852),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_875),
.B(n_861),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_836),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_873),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_883),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_887),
.B(n_851),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_885),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_869),
.B(n_851),
.Y(n_899)
);

INVx3_ASAP7_75t_SL g900 ( 
.A(n_879),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_873),
.B(n_839),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_884),
.B(n_850),
.Y(n_902)
);

AND2x6_ASAP7_75t_SL g903 ( 
.A(n_864),
.B(n_836),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_886),
.B(n_844),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_865),
.B(n_844),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_877),
.B(n_846),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_876),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_876),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_882),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_870),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_871),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_868),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_881),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_871),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_881),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_878),
.B(n_843),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_891),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_911),
.A2(n_889),
.B(n_874),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_909),
.B(n_867),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_894),
.B(n_880),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_900),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_896),
.Y(n_922)
);

AOI21xp33_ASAP7_75t_L g923 ( 
.A1(n_905),
.A2(n_866),
.B(n_889),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_910),
.B(n_868),
.Y(n_924)
);

INVx5_ASAP7_75t_L g925 ( 
.A(n_903),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_893),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_892),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_913),
.B(n_872),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_916),
.B(n_126),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_915),
.B(n_866),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_SL g931 ( 
.A1(n_904),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_895),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_930),
.B(n_920),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_922),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_926),
.B(n_901),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_917),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_917),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_927),
.B(n_901),
.Y(n_938)
);

AND2x4_ASAP7_75t_SL g939 ( 
.A(n_920),
.B(n_908),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_928),
.B(n_907),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_925),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_912),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_932),
.B(n_897),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_936),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_934),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_933),
.B(n_919),
.Y(n_946)
);

AOI32xp33_ASAP7_75t_L g947 ( 
.A1(n_943),
.A2(n_931),
.A3(n_929),
.B1(n_902),
.B2(n_924),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_937),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_SL g949 ( 
.A1(n_942),
.A2(n_921),
.B(n_923),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_937),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_949),
.B(n_941),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_L g952 ( 
.A1(n_947),
.A2(n_938),
.B(n_935),
.Y(n_952)
);

AOI21xp33_ASAP7_75t_L g953 ( 
.A1(n_945),
.A2(n_918),
.B(n_908),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_946),
.B(n_940),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_952),
.B(n_939),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_954),
.Y(n_956)
);

OAI222xp33_ASAP7_75t_L g957 ( 
.A1(n_951),
.A2(n_899),
.B1(n_906),
.B2(n_948),
.C1(n_944),
.C2(n_950),
.Y(n_957)
);

NAND2x1_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_953),
.Y(n_958)
);

AO21x1_ASAP7_75t_L g959 ( 
.A1(n_958),
.A2(n_955),
.B(n_957),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_959),
.A2(n_898),
.B(n_914),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_138),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_962),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_963),
.A2(n_141),
.B1(n_149),
.B2(n_150),
.Y(n_964)
);

OA22x2_ASAP7_75t_L g965 ( 
.A1(n_963),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_965),
.Y(n_966)
);

AOI31xp33_ASAP7_75t_L g967 ( 
.A1(n_964),
.A2(n_157),
.A3(n_159),
.B(n_160),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_SL g968 ( 
.A1(n_966),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_SL g969 ( 
.A1(n_967),
.A2(n_178),
.B1(n_180),
.B2(n_182),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_968),
.A2(n_183),
.B1(n_185),
.B2(n_188),
.Y(n_970)
);

XNOR2xp5_ASAP7_75t_L g971 ( 
.A(n_970),
.B(n_969),
.Y(n_971)
);

AOI222xp33_ASAP7_75t_L g972 ( 
.A1(n_971),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.C1(n_202),
.C2(n_203),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_972),
.B(n_207),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_973),
.A2(n_208),
.B1(n_214),
.B2(n_217),
.Y(n_974)
);


endmodule