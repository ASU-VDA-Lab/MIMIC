module fake_jpeg_1038_n_54 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_30),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_33)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_23),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_26),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.C(n_28),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_31),
.B(n_27),
.C(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

AOI322xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_33),
.A3(n_31),
.B1(n_27),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_29),
.C(n_6),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_7),
.Y(n_48)
);

AOI322xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.A3(n_49),
.B1(n_46),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_45),
.A3(n_42),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_5),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_8),
.B(n_11),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_13),
.C(n_14),
.Y(n_54)
);


endmodule