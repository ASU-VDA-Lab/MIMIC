module fake_jpeg_14951_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_27),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_80),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_76),
.B(n_82),
.Y(n_91)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_0),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_84),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_41),
.B1(n_48),
.B2(n_36),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_0),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_101),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_11),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_50),
.B(n_67),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_103),
.B(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_16),
.B1(n_18),
.B2(n_64),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_68),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_27),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_87),
.C(n_27),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_16),
.B1(n_18),
.B2(n_59),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_11),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_108),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_55),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_114),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_63),
.B(n_83),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_117),
.B(n_125),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_13),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_83),
.B(n_62),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_80),
.B1(n_59),
.B2(n_69),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_76),
.B1(n_82),
.B2(n_42),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_124),
.B1(n_100),
.B2(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_42),
.B1(n_61),
.B2(n_36),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_0),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_1),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_91),
.B(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_92),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_156),
.B(n_126),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_139),
.B(n_153),
.Y(n_167)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_104),
.B1(n_91),
.B2(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_128),
.B1(n_130),
.B2(n_124),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_145),
.B1(n_130),
.B2(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_96),
.B1(n_95),
.B2(n_57),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_21),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_144),
.Y(n_162)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_164),
.B1(n_25),
.B2(n_35),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_136),
.B(n_116),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_175),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_125),
.B(n_126),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_174),
.A2(n_78),
.B(n_13),
.C(n_14),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_121),
.B1(n_57),
.B2(n_114),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_177),
.B1(n_137),
.B2(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_66),
.B1(n_25),
.B2(n_85),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_85),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_21),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_132),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_153),
.B1(n_154),
.B2(n_135),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_134),
.C(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_189),
.C(n_174),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_145),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_134),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_138),
.C(n_150),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_142),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_135),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_196),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_181),
.B1(n_173),
.B2(n_178),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_44),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_78),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_167),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_178),
.B1(n_172),
.B2(n_158),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_198),
.B1(n_202),
.B2(n_196),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_213),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_157),
.B1(n_169),
.B2(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_172),
.B1(n_177),
.B2(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_179),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_211),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_165),
.B1(n_159),
.B2(n_166),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_158),
.B1(n_162),
.B2(n_180),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_164),
.B1(n_175),
.B2(n_26),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_13),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_14),
.C(n_19),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_191),
.A2(n_22),
.B1(n_26),
.B2(n_20),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_198),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_194),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_229),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_22),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_13),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_235),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_9),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_236),
.C(n_17),
.Y(n_239)
);

AOI321xp33_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_217),
.A3(n_220),
.B1(n_216),
.B2(n_219),
.C(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_203),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_240),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_249),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_35),
.C(n_30),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_30),
.C(n_28),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_244),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_14),
.C(n_21),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_21),
.C(n_23),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_24),
.C(n_23),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_24),
.C(n_2),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_254),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_222),
.B(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_236),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_1),
.C(n_3),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_260),
.B1(n_256),
.B2(n_6),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_1),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_3),
.C(n_4),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_269),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_1),
.B(n_3),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_266),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_4),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_4),
.C(n_5),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_4),
.B(n_5),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_265),
.B(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_5),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_261),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_273),
.B(n_270),
.C(n_271),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_274),
.B(n_7),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_280),
.B(n_7),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_6),
.C(n_7),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_8),
.Y(n_285)
);


endmodule