module real_jpeg_20006_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_96)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_60),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_27),
.B1(n_81),
.B2(n_90),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_10),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_27),
.B1(n_42),
.B2(n_43),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_12),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_25),
.A3(n_34),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_14),
.B(n_43),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_13),
.B(n_38),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_25),
.B(n_150),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_14),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_58)
);

BUFx3_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_100),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_98),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_71),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_19),
.B(n_71),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_54),
.C(n_63),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_20),
.A2(n_21),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_49),
.C(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_35),
.B2(n_38),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_25),
.B(n_51),
.Y(n_82)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_26),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_26),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_29),
.A2(n_32),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_34),
.A2(n_57),
.B(n_68),
.C(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_42),
.B(n_127),
.Y(n_126)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_47),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_45),
.A2(n_46),
.B1(n_108),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_45),
.A2(n_70),
.B1(n_111),
.B2(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_80),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_51),
.B(n_81),
.C(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_81),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_54),
.A2(n_63),
.B1(n_64),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_54),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_55),
.A2(n_58),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_55),
.A2(n_58),
.B1(n_119),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_55),
.A2(n_58),
.B1(n_59),
.B2(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_68),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_69),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_67),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_81),
.CON(n_80),
.SN(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_78),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_86),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_84),
.B2(n_85),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_157),
.B(n_163),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_143),
.B(n_156),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_131),
.B(n_142),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_120),
.B(n_130),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_112),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_133),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.C(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_159),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);


endmodule