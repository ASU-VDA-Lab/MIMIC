module fake_jpeg_25589_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_8),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_3),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_18),
.B1(n_28),
.B2(n_27),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_34),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_55),
.Y(n_64)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_17),
.B(n_29),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_19),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_4),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_5),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_21),
.B1(n_25),
.B2(n_10),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_7),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_58),
.B1(n_47),
.B2(n_12),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_77),
.B1(n_69),
.B2(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_58),
.B1(n_47),
.B2(n_13),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_67),
.B(n_71),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

AOI321xp33_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_74),
.A3(n_77),
.B1(n_7),
.B2(n_70),
.C(n_22),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_11),
.B(n_14),
.Y(n_88)
);


endmodule