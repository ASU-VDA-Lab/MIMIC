module fake_jpeg_7611_n_59 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_33),
.B(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_2),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_45),
.B(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_3),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_27),
.B1(n_13),
.B2(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_15),
.B1(n_20),
.B2(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_43),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_3),
.C(n_4),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_47),
.B(n_41),
.C(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_48),
.Y(n_55)
);

OAI322xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_55),
.A3(n_39),
.B1(n_40),
.B2(n_11),
.C1(n_16),
.C2(n_19),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_8),
.B(n_9),
.Y(n_59)
);


endmodule