module real_aes_9708_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_1802;
wire n_397;
wire n_1855;
wire n_1056;
wire n_727;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_1226;
wire n_525;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1564 ( .A1(n_0), .A2(n_144), .B1(n_1534), .B2(n_1555), .C(n_1565), .Y(n_1564) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_1), .A2(n_93), .B1(n_872), .B2(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1360 ( .A(n_2), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_2), .A2(n_8), .B1(n_749), .B2(n_1377), .Y(n_1376) );
AOI22xp5_ASAP7_75t_L g1533 ( .A1(n_3), .A2(n_128), .B1(n_1534), .B2(n_1538), .Y(n_1533) );
AOI22xp33_ASAP7_75t_SL g1070 ( .A1(n_4), .A2(n_16), .B1(n_822), .B2(n_1071), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_4), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_5), .A2(n_246), .B1(n_513), .B2(n_976), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_5), .A2(n_246), .B1(n_824), .B2(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1353 ( .A(n_6), .Y(n_1353) );
INVx1_ASAP7_75t_L g1019 ( .A(n_7), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_7), .A2(n_270), .B1(n_749), .B2(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1359 ( .A(n_8), .Y(n_1359) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_9), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_9), .A2(n_67), .B1(n_712), .B2(n_714), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_10), .A2(n_303), .B1(n_698), .B2(n_805), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_10), .A2(n_303), .B1(n_815), .B2(n_816), .Y(n_814) );
INVxp33_ASAP7_75t_SL g1065 ( .A(n_11), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_11), .A2(n_332), .B1(n_805), .B2(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g594 ( .A(n_12), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_12), .A2(n_223), .B1(n_614), .B2(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g965 ( .A(n_13), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_13), .A2(n_72), .B1(n_982), .B2(n_983), .Y(n_981) );
AOI221xp5_ASAP7_75t_L g1831 ( .A1(n_14), .A2(n_209), .B1(n_633), .B2(n_693), .C(n_1832), .Y(n_1831) );
OAI22xp33_ASAP7_75t_L g1843 ( .A1(n_14), .A2(n_326), .B1(n_1844), .B2(n_1847), .Y(n_1843) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_15), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_15), .A2(n_232), .B1(n_675), .B2(n_730), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1092 ( .A(n_16), .Y(n_1092) );
INVx1_ASAP7_75t_L g801 ( .A(n_17), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_17), .A2(n_57), .B1(n_633), .B2(n_693), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g1856 ( .A1(n_18), .A2(n_1857), .B1(n_1858), .B2(n_1859), .Y(n_1856) );
CKINVDCx5p33_ASAP7_75t_R g1857 ( .A(n_18), .Y(n_1857) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_19), .A2(n_259), .B1(n_756), .B2(n_1192), .Y(n_1261) );
AOI221xp5_ASAP7_75t_SL g1274 ( .A1(n_19), .A2(n_551), .B1(n_1275), .B2(n_1276), .C(n_1284), .Y(n_1274) );
INVx1_ASAP7_75t_L g1352 ( .A(n_20), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_20), .A2(n_65), .B1(n_753), .B2(n_983), .Y(n_1379) );
INVx1_ASAP7_75t_L g1566 ( .A(n_21), .Y(n_1566) );
INVxp33_ASAP7_75t_SL g792 ( .A(n_22), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_22), .A2(n_109), .B1(n_558), .B2(n_609), .Y(n_820) );
INVxp33_ASAP7_75t_L g733 ( .A(n_23), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_23), .A2(n_35), .B1(n_542), .B2(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g1442 ( .A(n_24), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1454 ( .A1(n_24), .A2(n_337), .B1(n_845), .B2(n_884), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_25), .A2(n_365), .B1(n_767), .B2(n_1034), .Y(n_1037) );
INVx1_ASAP7_75t_L g1043 ( .A(n_25), .Y(n_1043) );
XOR2x2_ASAP7_75t_L g1052 ( .A(n_26), .B(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1479 ( .A(n_27), .Y(n_1479) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_28), .A2(n_268), .B1(n_513), .B2(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g988 ( .A1(n_28), .A2(n_268), .B1(n_872), .B2(n_989), .Y(n_988) );
OAI211xp5_ASAP7_75t_L g886 ( .A1(n_29), .A2(n_654), .B(n_887), .C(n_890), .Y(n_886) );
INVx1_ASAP7_75t_L g918 ( .A(n_29), .Y(n_918) );
OAI222xp33_ASAP7_75t_L g573 ( .A1(n_30), .A2(n_84), .B1(n_238), .B2(n_574), .C1(n_577), .C2(n_583), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_30), .A2(n_197), .B1(n_633), .B2(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g1410 ( .A(n_31), .Y(n_1410) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_31), .A2(n_210), .B1(n_940), .B2(n_994), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g1784 ( .A1(n_32), .A2(n_370), .B1(n_1785), .B2(n_1786), .Y(n_1784) );
INVxp67_ASAP7_75t_SL g1819 ( .A(n_32), .Y(n_1819) );
AOI22xp33_ASAP7_75t_SL g1884 ( .A1(n_33), .A2(n_97), .B1(n_510), .B2(n_688), .Y(n_1884) );
AOI22xp33_ASAP7_75t_L g1893 ( .A1(n_33), .A2(n_97), .B1(n_614), .B2(n_714), .Y(n_1893) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_34), .Y(n_929) );
INVx1_ASAP7_75t_L g727 ( .A(n_35), .Y(n_727) );
INVx1_ASAP7_75t_L g1473 ( .A(n_36), .Y(n_1473) );
INVx1_ASAP7_75t_L g590 ( .A(n_37), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_37), .A2(n_190), .B1(n_510), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g1330 ( .A(n_38), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g1335 ( .A1(n_38), .A2(n_231), .B1(n_845), .B2(n_848), .Y(n_1335) );
INVx1_ASAP7_75t_L g954 ( .A(n_39), .Y(n_954) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_39), .A2(n_168), .B1(n_940), .B2(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g789 ( .A(n_40), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_41), .A2(n_143), .B1(n_712), .B2(n_1071), .Y(n_1304) );
INVxp67_ASAP7_75t_SL g1316 ( .A(n_41), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_42), .A2(n_87), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_42), .A2(n_87), .B1(n_547), .B2(n_702), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g1236 ( .A1(n_43), .A2(n_501), .B(n_1000), .C(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1270 ( .A(n_43), .Y(n_1270) );
INVx1_ASAP7_75t_L g381 ( .A(n_44), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g1293 ( .A1(n_45), .A2(n_501), .B(n_1294), .C(n_1295), .Y(n_1293) );
INVx1_ASAP7_75t_L g1309 ( .A(n_45), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_46), .A2(n_63), .B1(n_390), .B2(n_500), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1222 ( .A1(n_46), .A2(n_355), .B1(n_845), .B2(n_884), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_47), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_47), .A2(n_203), .B1(n_749), .B2(n_750), .Y(n_1174) );
AOI22xp5_ASAP7_75t_L g1589 ( .A1(n_48), .A2(n_152), .B1(n_1534), .B2(n_1538), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_49), .A2(n_239), .B1(n_638), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_49), .A2(n_239), .B1(n_614), .B2(n_702), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_50), .A2(n_124), .B1(n_845), .B2(n_848), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_50), .A2(n_124), .B1(n_515), .B2(n_805), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_51), .A2(n_357), .B1(n_638), .B2(n_640), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_51), .A2(n_251), .B1(n_816), .B2(n_875), .Y(n_874) );
INVxp33_ASAP7_75t_L g1881 ( .A(n_52), .Y(n_1881) );
AOI22xp33_ASAP7_75t_L g1895 ( .A1(n_52), .A2(n_300), .B1(n_621), .B2(n_986), .Y(n_1895) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_53), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_53), .A2(n_299), .B1(n_805), .B2(n_809), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_54), .A2(n_324), .B1(n_976), .B2(n_1190), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_54), .A2(n_324), .B1(n_547), .B2(n_989), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_55), .A2(n_206), .B1(n_983), .B2(n_1192), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_55), .A2(n_206), .B1(n_767), .B2(n_1034), .Y(n_1419) );
AO221x2_ASAP7_75t_L g1552 ( .A1(n_56), .A2(n_282), .B1(n_1553), .B2(n_1555), .C(n_1557), .Y(n_1552) );
INVxp33_ASAP7_75t_SL g796 ( .A(n_57), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_58), .A2(n_89), .B1(n_902), .B2(n_906), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_58), .A2(n_89), .B1(n_547), .B2(n_1181), .Y(n_1184) );
INVx1_ASAP7_75t_L g1782 ( .A(n_59), .Y(n_1782) );
INVxp33_ASAP7_75t_SL g859 ( .A(n_60), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_60), .A2(n_174), .B1(n_815), .B2(n_816), .Y(n_877) );
INVxp67_ASAP7_75t_SL g1102 ( .A(n_61), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_61), .A2(n_226), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_62), .A2(n_367), .B1(n_902), .B2(n_906), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_62), .A2(n_367), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_63), .A2(n_191), .B1(n_438), .B2(n_1203), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1238 ( .A1(n_64), .A2(n_146), .B1(n_390), .B2(n_500), .Y(n_1238) );
INVx1_ASAP7_75t_L g1267 ( .A(n_64), .Y(n_1267) );
INVx1_ASAP7_75t_L g1356 ( .A(n_65), .Y(n_1356) );
INVx1_ASAP7_75t_L g1363 ( .A(n_66), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_66), .A2(n_264), .B1(n_986), .B2(n_987), .Y(n_1386) );
INVxp33_ASAP7_75t_SL g678 ( .A(n_67), .Y(n_678) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_68), .A2(n_652), .B1(n_717), .B2(n_718), .Y(n_651) );
CKINVDCx14_ASAP7_75t_R g717 ( .A(n_68), .Y(n_717) );
INVx1_ASAP7_75t_L g957 ( .A(n_69), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_69), .A2(n_182), .B1(n_657), .B2(n_766), .Y(n_992) );
OAI211xp5_ASAP7_75t_L g999 ( .A1(n_69), .A2(n_501), .B(n_1000), .C(n_1002), .Y(n_999) );
XNOR2xp5_ASAP7_75t_L g1011 ( .A(n_70), .B(n_1012), .Y(n_1011) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_71), .Y(n_589) );
INVx1_ASAP7_75t_L g969 ( .A(n_72), .Y(n_969) );
OAI211xp5_ASAP7_75t_L g1006 ( .A1(n_72), .A2(n_654), .B(n_1007), .C(n_1008), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_73), .A2(n_1226), .B1(n_1286), .B2(n_1287), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_73), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_74), .A2(n_313), .B1(n_1534), .B2(n_1538), .Y(n_1572) );
AOI22xp5_ASAP7_75t_L g1521 ( .A1(n_75), .A2(n_350), .B1(n_1522), .B2(n_1530), .Y(n_1521) );
INVx1_ASAP7_75t_L g662 ( .A(n_76), .Y(n_662) );
INVx1_ASAP7_75t_L g448 ( .A(n_77), .Y(n_448) );
INVx1_ASAP7_75t_L g1471 ( .A(n_78), .Y(n_1471) );
INVx1_ASAP7_75t_L g966 ( .A(n_79), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_79), .A2(n_341), .B1(n_749), .B2(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g1211 ( .A(n_80), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g1458 ( .A(n_81), .Y(n_1458) );
AO22x1_ASAP7_75t_L g1575 ( .A1(n_82), .A2(n_262), .B1(n_1538), .B2(n_1576), .Y(n_1575) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_83), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_83), .A2(n_310), .B1(n_696), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g600 ( .A(n_84), .Y(n_600) );
XOR2xp5_ASAP7_75t_L g829 ( .A(n_85), .B(n_830), .Y(n_829) );
AO22x1_ASAP7_75t_L g1577 ( .A1(n_85), .A2(n_260), .B1(n_1522), .B2(n_1530), .Y(n_1577) );
INVx1_ASAP7_75t_L g839 ( .A(n_86), .Y(n_839) );
OAI222xp33_ASAP7_75t_L g852 ( .A1(n_86), .A2(n_187), .B1(n_284), .B2(n_480), .C1(n_853), .C2(n_856), .Y(n_852) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_88), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_88), .A2(n_104), .B1(n_1279), .B2(n_1282), .Y(n_1278) );
INVx1_ASAP7_75t_L g1302 ( .A(n_90), .Y(n_1302) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_91), .A2(n_271), .B1(n_696), .B2(n_924), .C(n_926), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_91), .A2(n_271), .B1(n_939), .B2(n_940), .Y(n_938) );
OAI21xp33_ASAP7_75t_SL g834 ( .A1(n_92), .A2(n_835), .B(n_838), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_92), .A2(n_318), .B1(n_750), .B2(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g1047 ( .A(n_93), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1758 ( .A(n_94), .Y(n_1758) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_95), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_96), .A2(n_256), .B1(n_902), .B2(n_906), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_96), .A2(n_256), .B1(n_824), .B2(n_939), .Y(n_945) );
BUFx2_ASAP7_75t_L g460 ( .A(n_98), .Y(n_460) );
BUFx2_ASAP7_75t_L g506 ( .A(n_98), .Y(n_506) );
INVx1_ASAP7_75t_L g535 ( .A(n_98), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_99), .A2(n_258), .B1(n_706), .B2(n_737), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g1086 ( .A(n_99), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_100), .A2(n_361), .B1(n_614), .B2(n_1075), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_100), .A2(n_361), .B1(n_805), .B2(n_809), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_101), .A2(n_336), .B1(n_756), .B2(n_1192), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_101), .A2(n_336), .B1(n_767), .B2(n_771), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_102), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_102), .A2(n_317), .B1(n_480), .B2(n_675), .Y(n_674) );
AO22x2_ASAP7_75t_L g568 ( .A1(n_103), .A2(n_569), .B1(n_570), .B2(n_648), .Y(n_568) );
INVx1_ASAP7_75t_L g648 ( .A(n_103), .Y(n_648) );
INVxp67_ASAP7_75t_SL g1260 ( .A(n_104), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_105), .A2(n_294), .B1(n_556), .B2(n_737), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_105), .A2(n_294), .B1(n_529), .B2(n_693), .Y(n_1083) );
INVx1_ASAP7_75t_L g1396 ( .A(n_106), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_106), .A2(n_363), .B1(n_513), .B2(n_911), .Y(n_1416) );
XNOR2xp5_ASAP7_75t_L g1146 ( .A(n_107), .B(n_1147), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_108), .Y(n_899) );
INVx1_ASAP7_75t_L g788 ( .A(n_109), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_110), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_111), .A2(n_251), .B1(n_529), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_111), .A2(n_357), .B1(n_870), .B2(n_873), .Y(n_869) );
INVx1_ASAP7_75t_L g1506 ( .A(n_112), .Y(n_1506) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_113), .A2(n_114), .B1(n_902), .B2(n_906), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_113), .A2(n_114), .B1(n_547), .B2(n_1311), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_115), .A2(n_122), .B1(n_583), .B2(n_1401), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_115), .A2(n_122), .B1(n_675), .B2(n_730), .Y(n_1405) );
AO221x1_ASAP7_75t_L g1540 ( .A1(n_116), .A2(n_129), .B1(n_1534), .B2(n_1538), .C(n_1541), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_117), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_117), .A2(n_249), .B1(n_510), .B2(n_526), .Y(n_525) );
AO221x1_ASAP7_75t_L g1547 ( .A1(n_118), .A2(n_330), .B1(n_1534), .B2(n_1538), .C(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1223 ( .A(n_119), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_120), .A2(n_275), .B1(n_609), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_120), .A2(n_275), .B1(n_644), .B2(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g1500 ( .A(n_121), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_123), .A2(n_162), .B1(n_672), .B2(n_761), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_123), .A2(n_162), .B1(n_986), .B2(n_987), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_125), .Y(n_927) );
INVx1_ASAP7_75t_L g1482 ( .A(n_126), .Y(n_1482) );
OAI22xp33_ASAP7_75t_SL g1512 ( .A1(n_126), .A2(n_229), .B1(n_390), .B2(n_902), .Y(n_1512) );
INVx1_ASAP7_75t_L g1545 ( .A(n_127), .Y(n_1545) );
AOI22xp5_ASAP7_75t_L g1588 ( .A1(n_130), .A2(n_161), .B1(n_1522), .B2(n_1530), .Y(n_1588) );
INVx1_ASAP7_75t_L g1828 ( .A(n_131), .Y(n_1828) );
OAI22xp33_ASAP7_75t_L g1848 ( .A1(n_131), .A2(n_209), .B1(n_1849), .B2(n_1851), .Y(n_1848) );
INVxp33_ASAP7_75t_SL g1878 ( .A(n_132), .Y(n_1878) );
AOI22xp33_ASAP7_75t_L g1896 ( .A1(n_132), .A2(n_230), .B1(n_616), .B2(n_1897), .Y(n_1896) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_133), .A2(n_266), .B1(n_737), .B2(n_1123), .Y(n_1122) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_133), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_134), .A2(n_220), .B1(n_560), .B2(n_616), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_134), .A2(n_220), .B1(n_638), .B2(n_640), .Y(n_637) );
XOR2xp5_ASAP7_75t_L g1425 ( .A(n_135), .B(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1788 ( .A(n_136), .Y(n_1788) );
OAI221xp5_ASAP7_75t_L g1809 ( .A1(n_136), .A2(n_1810), .B1(n_1812), .B2(n_1817), .C(n_1820), .Y(n_1809) );
INVx1_ASAP7_75t_L g1558 ( .A(n_137), .Y(n_1558) );
INVx1_ASAP7_75t_L g734 ( .A(n_138), .Y(n_734) );
INVx1_ASAP7_75t_L g1018 ( .A(n_139), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_139), .A2(n_272), .B1(n_756), .B2(n_982), .Y(n_1031) );
INVx1_ASAP7_75t_L g1106 ( .A(n_140), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_140), .A2(n_314), .B1(n_856), .B2(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g1885 ( .A1(n_141), .A2(n_308), .B1(n_633), .B2(n_635), .Y(n_1885) );
AOI22xp33_ASAP7_75t_L g1892 ( .A1(n_141), .A2(n_308), .B1(n_621), .B2(n_706), .Y(n_1892) );
INVxp33_ASAP7_75t_SL g1865 ( .A(n_142), .Y(n_1865) );
AOI22xp33_ASAP7_75t_L g1887 ( .A1(n_142), .A2(n_353), .B1(n_638), .B2(n_1888), .Y(n_1887) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_143), .Y(n_1320) );
INVx1_ASAP7_75t_L g1496 ( .A(n_145), .Y(n_1496) );
OAI22xp33_ASAP7_75t_L g1502 ( .A1(n_145), .A2(n_151), .B1(n_845), .B2(n_848), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1228 ( .A1(n_146), .A2(n_356), .B1(n_884), .B2(n_885), .Y(n_1228) );
INVxp33_ASAP7_75t_L g745 ( .A(n_147), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_147), .A2(n_334), .B1(n_756), .B2(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g1439 ( .A(n_148), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_148), .A2(n_301), .B1(n_848), .B2(n_885), .Y(n_1460) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_149), .A2(n_782), .B1(n_825), .B2(n_826), .Y(n_781) );
INVxp67_ASAP7_75t_L g825 ( .A(n_149), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_150), .A2(n_192), .B1(n_390), .B2(n_500), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_150), .A2(n_284), .B1(n_540), .B2(n_873), .Y(n_876) );
INVx1_ASAP7_75t_L g1499 ( .A(n_151), .Y(n_1499) );
INVx1_ASAP7_75t_L g1526 ( .A(n_153), .Y(n_1526) );
OAI211xp5_ASAP7_75t_L g1162 ( .A1(n_154), .A2(n_501), .B(n_1163), .C(n_1165), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_154), .A2(n_269), .B1(n_1034), .B2(n_1179), .Y(n_1183) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_155), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_155), .A2(n_305), .B1(n_518), .B2(n_529), .Y(n_528) );
INVxp33_ASAP7_75t_SL g1098 ( .A(n_156), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_156), .A2(n_200), .B1(n_491), .B2(n_1111), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1394 ( .A(n_157), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_158), .A2(n_372), .B1(n_390), .B2(n_500), .Y(n_1292) );
INVx1_ASAP7_75t_L g1307 ( .A(n_158), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_159), .A2(n_244), .B1(n_759), .B2(n_1170), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_159), .A2(n_244), .B1(n_547), .B2(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_160), .A2(n_255), .B1(n_672), .B2(n_753), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_160), .A2(n_255), .B1(n_657), .B2(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1549 ( .A(n_163), .Y(n_1549) );
INVx1_ASAP7_75t_L g1871 ( .A(n_164), .Y(n_1871) );
OAI22xp5_ASAP7_75t_L g1876 ( .A1(n_164), .A2(n_298), .B1(n_480), .B2(n_856), .Y(n_1876) );
AO22x2_ASAP7_75t_SL g1093 ( .A1(n_165), .A2(n_1094), .B1(n_1095), .B2(n_1138), .Y(n_1093) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_165), .Y(n_1094) );
INVx1_ASAP7_75t_L g1450 ( .A(n_166), .Y(n_1450) );
OAI22xp33_ASAP7_75t_SL g1465 ( .A1(n_166), .A2(n_179), .B1(n_390), .B2(n_902), .Y(n_1465) );
INVxp33_ASAP7_75t_SL g1056 ( .A(n_167), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_167), .A2(n_176), .B1(n_515), .B2(n_693), .Y(n_1080) );
INVx1_ASAP7_75t_L g955 ( .A(n_168), .Y(n_955) );
INVx1_ASAP7_75t_L g1527 ( .A(n_169), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_169), .B(n_1525), .Y(n_1532) );
INVxp33_ASAP7_75t_SL g669 ( .A(n_170), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_170), .A2(n_342), .B1(n_706), .B2(n_709), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_171), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_172), .A2(n_237), .B1(n_694), .B2(n_761), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_172), .A2(n_237), .B1(n_767), .B2(n_1034), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_173), .A2(n_185), .B1(n_845), .B2(n_848), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_173), .A2(n_319), .B1(n_909), .B2(n_912), .C(n_914), .Y(n_908) );
INVxp33_ASAP7_75t_L g858 ( .A(n_174), .Y(n_858) );
INVx2_ASAP7_75t_L g393 ( .A(n_175), .Y(n_393) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_176), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1793 ( .A1(n_177), .A2(n_215), .B1(n_1794), .B2(n_1798), .Y(n_1793) );
INVx1_ASAP7_75t_L g1836 ( .A(n_177), .Y(n_1836) );
INVxp33_ASAP7_75t_L g1864 ( .A(n_178), .Y(n_1864) );
AOI22xp33_ASAP7_75t_L g1890 ( .A1(n_178), .A2(n_345), .B1(n_644), .B2(n_694), .Y(n_1890) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_179), .A2(n_297), .B1(n_547), .B2(n_824), .Y(n_1452) );
INVx1_ASAP7_75t_L g1325 ( .A(n_180), .Y(n_1325) );
OAI22xp33_ASAP7_75t_L g1338 ( .A1(n_180), .A2(n_372), .B1(n_884), .B2(n_885), .Y(n_1338) );
BUFx3_ASAP7_75t_L g415 ( .A(n_181), .Y(n_415) );
INVx1_ASAP7_75t_L g433 ( .A(n_181), .Y(n_433) );
INVx1_ASAP7_75t_L g961 ( .A(n_182), .Y(n_961) );
INVx1_ASAP7_75t_L g490 ( .A(n_183), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_183), .A2(n_263), .B1(n_556), .B2(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g442 ( .A(n_184), .Y(n_442) );
INVx1_ASAP7_75t_L g915 ( .A(n_185), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g1413 ( .A1(n_186), .A2(n_252), .B1(n_513), .B2(n_976), .Y(n_1413) );
AOI22xp33_ASAP7_75t_SL g1420 ( .A1(n_186), .A2(n_252), .B1(n_824), .B2(n_994), .Y(n_1420) );
INVx1_ASAP7_75t_L g840 ( .A(n_187), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_188), .A2(n_368), .B1(n_515), .B2(n_518), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_188), .A2(n_368), .B1(n_540), .B2(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g1393 ( .A(n_189), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g1417 ( .A1(n_189), .A2(n_321), .B1(n_983), .B2(n_1192), .Y(n_1417) );
INVx1_ASAP7_75t_L g587 ( .A(n_190), .Y(n_587) );
OAI211xp5_ASAP7_75t_SL g1206 ( .A1(n_191), .A2(n_501), .B(n_1207), .C(n_1210), .Y(n_1206) );
INVx1_ASAP7_75t_L g842 ( .A(n_192), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_193), .A2(n_248), .B1(n_909), .B2(n_912), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_193), .A2(n_248), .B1(n_560), .B2(n_816), .Y(n_1120) );
INVx1_ASAP7_75t_L g1790 ( .A(n_194), .Y(n_1790) );
OAI211xp5_ASAP7_75t_SL g1821 ( .A1(n_194), .A2(n_1822), .B(n_1824), .C(n_1833), .Y(n_1821) );
INVx1_ASAP7_75t_L g425 ( .A(n_195), .Y(n_425) );
INVx1_ASAP7_75t_L g1332 ( .A(n_196), .Y(n_1332) );
OAI211xp5_ASAP7_75t_L g1336 ( .A1(n_196), .A2(n_654), .B(n_835), .C(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g585 ( .A(n_197), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g1110 ( .A1(n_198), .A2(n_364), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
AOI22xp33_ASAP7_75t_SL g1121 ( .A1(n_198), .A2(n_364), .B1(n_540), .B2(n_542), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_199), .A2(n_355), .B1(n_756), .B2(n_761), .Y(n_1196) );
INVx1_ASAP7_75t_L g1217 ( .A(n_199), .Y(n_1217) );
INVx1_ASAP7_75t_L g1104 ( .A(n_200), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_201), .A2(n_1290), .B1(n_1339), .B2(n_1340), .Y(n_1289) );
INVx1_ASAP7_75t_L g1340 ( .A(n_201), .Y(n_1340) );
INVx1_ASAP7_75t_L g1155 ( .A(n_202), .Y(n_1155) );
INVx1_ASAP7_75t_L g1158 ( .A(n_203), .Y(n_1158) );
INVx1_ASAP7_75t_L g728 ( .A(n_204), .Y(n_728) );
XNOR2xp5_ASAP7_75t_L g879 ( .A(n_205), .B(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g1483 ( .A(n_207), .Y(n_1483) );
OAI211xp5_ASAP7_75t_SL g1510 ( .A1(n_207), .A2(n_501), .B(n_1163), .C(n_1511), .Y(n_1510) );
AO22x2_ASAP7_75t_L g720 ( .A1(n_208), .A2(n_721), .B1(n_775), .B2(n_776), .Y(n_720) );
INVx1_ASAP7_75t_L g775 ( .A(n_208), .Y(n_775) );
INVx1_ASAP7_75t_L g1408 ( .A(n_210), .Y(n_1408) );
INVx1_ASAP7_75t_L g458 ( .A(n_211), .Y(n_458) );
INVx1_ASAP7_75t_L g1764 ( .A(n_211), .Y(n_1764) );
INVxp33_ASAP7_75t_SL g463 ( .A(n_212), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_212), .A2(n_247), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g1212 ( .A(n_213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1303 ( .A(n_214), .Y(n_1303) );
INVx1_ASAP7_75t_L g1840 ( .A(n_215), .Y(n_1840) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_216), .A2(n_219), .B1(n_515), .B2(n_693), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_216), .A2(n_219), .B1(n_706), .B2(n_737), .Y(n_813) );
INVxp67_ASAP7_75t_L g1370 ( .A(n_217), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_217), .A2(n_302), .B1(n_940), .B2(n_994), .Y(n_1387) );
INVx1_ASAP7_75t_L g1023 ( .A(n_218), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_218), .A2(n_338), .B1(n_480), .B2(n_856), .Y(n_1044) );
INVxp67_ASAP7_75t_SL g1435 ( .A(n_221), .Y(n_1435) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_221), .A2(n_344), .B1(n_824), .B2(n_872), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_222), .A2(n_362), .B1(n_513), .B2(n_976), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_222), .A2(n_362), .B1(n_712), .B2(n_774), .Y(n_1035) );
INVx1_ASAP7_75t_L g593 ( .A(n_223), .Y(n_593) );
INVx1_ASAP7_75t_L g1542 ( .A(n_224), .Y(n_1542) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_225), .A2(n_374), .B1(n_1522), .B2(n_1530), .Y(n_1573) );
INVxp33_ASAP7_75t_SL g1099 ( .A(n_226), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_227), .A2(n_311), .B1(n_774), .B2(n_872), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_227), .A2(n_311), .B1(n_902), .B2(n_906), .Y(n_1205) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_228), .A2(n_319), .B1(n_884), .B2(n_885), .Y(n_883) );
INVx1_ASAP7_75t_L g900 ( .A(n_228), .Y(n_900) );
INVx1_ASAP7_75t_L g1486 ( .A(n_229), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1879 ( .A(n_230), .Y(n_1879) );
INVx1_ASAP7_75t_L g1323 ( .A(n_231), .Y(n_1323) );
INVxp67_ASAP7_75t_SL g1062 ( .A(n_232), .Y(n_1062) );
INVxp33_ASAP7_75t_L g724 ( .A(n_233), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_233), .A2(n_327), .B1(n_547), .B2(n_774), .Y(n_773) );
INVxp33_ASAP7_75t_L g744 ( .A(n_234), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_234), .A2(n_290), .B1(n_630), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_235), .A2(n_359), .B1(n_753), .B2(n_756), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_235), .A2(n_359), .B1(n_766), .B2(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g1101 ( .A(n_236), .Y(n_1101) );
INVx1_ASAP7_75t_L g599 ( .A(n_238), .Y(n_599) );
INVx1_ASAP7_75t_L g1064 ( .A(n_240), .Y(n_1064) );
INVx1_ASAP7_75t_L g1431 ( .A(n_241), .Y(n_1431) );
INVxp33_ASAP7_75t_SL g665 ( .A(n_242), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_242), .A2(n_257), .B1(n_644), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g1154 ( .A(n_243), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_245), .A2(n_315), .B1(n_845), .B2(n_848), .Y(n_1233) );
INVx1_ASAP7_75t_L g1249 ( .A(n_245), .Y(n_1249) );
INVxp33_ASAP7_75t_SL g472 ( .A(n_247), .Y(n_472) );
INVxp33_ASAP7_75t_SL g418 ( .A(n_249), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_250), .A2(n_276), .B1(n_756), .B2(n_761), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_250), .A2(n_276), .B1(n_986), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1232 ( .A(n_253), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_254), .A2(n_287), .B1(n_976), .B2(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1221 ( .A(n_254), .Y(n_1221) );
INVx1_ASAP7_75t_L g656 ( .A(n_257), .Y(n_656) );
INVxp67_ASAP7_75t_SL g1089 ( .A(n_258), .Y(n_1089) );
INVxp67_ASAP7_75t_SL g1277 ( .A(n_259), .Y(n_1277) );
INVx1_ASAP7_75t_L g1487 ( .A(n_261), .Y(n_1487) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_261), .A2(n_273), .B1(n_500), .B2(n_906), .Y(n_1509) );
INVxp33_ASAP7_75t_SL g497 ( .A(n_263), .Y(n_497) );
INVxp33_ASAP7_75t_L g1367 ( .A(n_264), .Y(n_1367) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_265), .Y(n_897) );
INVxp33_ASAP7_75t_L g1137 ( .A(n_266), .Y(n_1137) );
BUFx3_ASAP7_75t_L g417 ( .A(n_267), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_267), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_269), .A2(n_340), .B1(n_390), .B2(n_500), .Y(n_1166) );
INVx1_ASAP7_75t_L g1016 ( .A(n_270), .Y(n_1016) );
INVx1_ASAP7_75t_L g1021 ( .A(n_272), .Y(n_1021) );
OAI22xp5_ASAP7_75t_L g1503 ( .A1(n_273), .A2(n_280), .B1(n_884), .B2(n_885), .Y(n_1503) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_274), .Y(n_389) );
INVx1_ASAP7_75t_L g537 ( .A(n_274), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_274), .B(n_349), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_274), .B(n_467), .Y(n_1804) );
AO22x2_ASAP7_75t_L g402 ( .A1(n_277), .A2(n_403), .B1(n_566), .B2(n_567), .Y(n_402) );
INVx1_ASAP7_75t_L g566 ( .A(n_277), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_278), .A2(n_322), .B1(n_644), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_278), .A2(n_322), .B1(n_609), .B2(n_621), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g1459 ( .A(n_279), .Y(n_1459) );
INVx1_ASAP7_75t_L g1497 ( .A(n_280), .Y(n_1497) );
INVx1_ASAP7_75t_L g1231 ( .A(n_281), .Y(n_1231) );
XNOR2xp5_ASAP7_75t_L g1466 ( .A(n_283), .B(n_1467), .Y(n_1466) );
INVx2_ASAP7_75t_L g410 ( .A(n_285), .Y(n_410) );
OR2x2_ASAP7_75t_L g1846 ( .A(n_285), .B(n_1764), .Y(n_1846) );
INVx1_ASAP7_75t_L g1348 ( .A(n_286), .Y(n_1348) );
INVxp67_ASAP7_75t_SL g1220 ( .A(n_287), .Y(n_1220) );
INVx1_ASAP7_75t_L g603 ( .A(n_288), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_288), .A2(n_293), .B1(n_609), .B2(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g1867 ( .A(n_289), .Y(n_1867) );
INVxp33_ASAP7_75t_L g742 ( .A(n_290), .Y(n_742) );
INVxp33_ASAP7_75t_SL g785 ( .A(n_291), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_291), .A2(n_295), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g1507 ( .A(n_292), .Y(n_1507) );
INVx1_ASAP7_75t_L g597 ( .A(n_293), .Y(n_597) );
INVxp33_ASAP7_75t_SL g786 ( .A(n_295), .Y(n_786) );
OAI211xp5_ASAP7_75t_L g1229 ( .A1(n_296), .A2(n_654), .B(n_1007), .C(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1250 ( .A(n_296), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1462 ( .A1(n_297), .A2(n_337), .B1(n_500), .B2(n_906), .Y(n_1462) );
INVx1_ASAP7_75t_L g1872 ( .A(n_298), .Y(n_1872) );
INVxp33_ASAP7_75t_SL g797 ( .A(n_299), .Y(n_797) );
INVxp67_ASAP7_75t_SL g1875 ( .A(n_300), .Y(n_1875) );
INVx1_ASAP7_75t_L g1437 ( .A(n_301), .Y(n_1437) );
INVx1_ASAP7_75t_L g1368 ( .A(n_302), .Y(n_1368) );
AO22x2_ASAP7_75t_L g950 ( .A1(n_304), .A2(n_951), .B1(n_995), .B2(n_996), .Y(n_950) );
INVxp67_ASAP7_75t_L g995 ( .A(n_304), .Y(n_995) );
INVx1_ASAP7_75t_L g435 ( .A(n_305), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_306), .A2(n_348), .B1(n_510), .B2(n_511), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_306), .A2(n_348), .B1(n_545), .B2(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g1451 ( .A(n_307), .Y(n_1451) );
OAI211xp5_ASAP7_75t_SL g1463 ( .A1(n_307), .A2(n_501), .B(n_1163), .C(n_1464), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_309), .A2(n_346), .B1(n_574), .B2(n_583), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_309), .A2(n_346), .B1(n_675), .B2(n_1132), .Y(n_1365) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_310), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g1791 ( .A1(n_312), .A2(n_351), .B1(n_548), .B2(n_1792), .Y(n_1791) );
OAI22xp5_ASAP7_75t_L g1801 ( .A1(n_312), .A2(n_351), .B1(n_1802), .B2(n_1805), .Y(n_1801) );
AOI222xp33_ASAP7_75t_L g1751 ( .A1(n_313), .A2(n_1752), .B1(n_1853), .B2(n_1855), .C1(n_1898), .C2(n_1902), .Y(n_1751) );
INVx1_ASAP7_75t_L g1755 ( .A(n_313), .Y(n_1755) );
INVx1_ASAP7_75t_L g1107 ( .A(n_314), .Y(n_1107) );
INVx1_ASAP7_75t_L g1242 ( .A(n_315), .Y(n_1242) );
INVx1_ASAP7_75t_L g1407 ( .A(n_316), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_316), .A2(n_352), .B1(n_987), .B2(n_1034), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_317), .Y(n_660) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_318), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_320), .Y(n_962) );
INVx1_ASAP7_75t_L g1399 ( .A(n_321), .Y(n_1399) );
INVx1_ASAP7_75t_L g790 ( .A(n_323), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_325), .A2(n_340), .B1(n_845), .B2(n_884), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_325), .A2(n_354), .B1(n_982), .B2(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1830 ( .A(n_326), .Y(n_1830) );
INVxp33_ASAP7_75t_L g725 ( .A(n_327), .Y(n_725) );
INVx1_ASAP7_75t_L g1476 ( .A(n_328), .Y(n_1476) );
INVx1_ASAP7_75t_L g731 ( .A(n_329), .Y(n_731) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_331), .B(n_381), .Y(n_1529) );
AND3x2_ASAP7_75t_L g1537 ( .A(n_331), .B(n_381), .C(n_1526), .Y(n_1537) );
INVxp33_ASAP7_75t_SL g1057 ( .A(n_332), .Y(n_1057) );
INVx2_ASAP7_75t_L g394 ( .A(n_333), .Y(n_394) );
INVx1_ASAP7_75t_L g739 ( .A(n_334), .Y(n_739) );
INVx1_ASAP7_75t_L g1297 ( .A(n_335), .Y(n_1297) );
INVx1_ASAP7_75t_L g1022 ( .A(n_338), .Y(n_1022) );
INVx1_ASAP7_75t_L g793 ( .A(n_339), .Y(n_793) );
INVx1_ASAP7_75t_L g971 ( .A(n_341), .Y(n_971) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_342), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_343), .Y(n_891) );
INVxp67_ASAP7_75t_SL g1433 ( .A(n_344), .Y(n_1433) );
INVxp67_ASAP7_75t_SL g1870 ( .A(n_345), .Y(n_1870) );
INVx1_ASAP7_75t_L g1430 ( .A(n_347), .Y(n_1430) );
INVx1_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
INVx2_ASAP7_75t_L g467 ( .A(n_349), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g1389 ( .A(n_350), .B(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1404 ( .A(n_352), .Y(n_1404) );
INVxp33_ASAP7_75t_L g1868 ( .A(n_353), .Y(n_1868) );
INVx1_ASAP7_75t_L g1151 ( .A(n_354), .Y(n_1151) );
INVx1_ASAP7_75t_L g1246 ( .A(n_356), .Y(n_1246) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_358), .Y(n_892) );
INVx1_ASAP7_75t_L g1296 ( .A(n_360), .Y(n_1296) );
INVx1_ASAP7_75t_L g1397 ( .A(n_363), .Y(n_1397) );
INVx1_ASAP7_75t_L g1049 ( .A(n_365), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_366), .A2(n_373), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
INVxp33_ASAP7_75t_L g1134 ( .A(n_366), .Y(n_1134) );
INVx1_ASAP7_75t_L g1781 ( .A(n_369), .Y(n_1781) );
INVxp33_ASAP7_75t_SL g1818 ( .A(n_370), .Y(n_1818) );
INVx1_ASAP7_75t_L g1443 ( .A(n_371), .Y(n_1443) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_373), .Y(n_1135) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_397), .B(n_1515), .Y(n_375) );
HB1xp67_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1854 ( .A(n_379), .B(n_385), .Y(n_1854) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1901 ( .A(n_380), .Y(n_1901) );
NAND2xp5_ASAP7_75t_L g1906 ( .A(n_380), .B(n_382), .Y(n_1906) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1900 ( .A(n_382), .B(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x6_ASAP7_75t_L g505 ( .A(n_387), .B(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g679 ( .A(n_387), .B(n_506), .Y(n_679) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g523 ( .A(n_388), .B(n_396), .Y(n_523) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_389), .B(n_466), .Y(n_1263) );
INVx8_ASAP7_75t_L g498 ( .A(n_390), .Y(n_498) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
OR2x6_ASAP7_75t_L g500 ( .A(n_391), .B(n_465), .Y(n_500) );
INVx2_ASAP7_75t_SL g917 ( .A(n_391), .Y(n_917) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_391), .Y(n_928) );
INVx1_ASAP7_75t_L g1329 ( .A(n_391), .Y(n_1329) );
HB1xp67_ASAP7_75t_L g1441 ( .A(n_391), .Y(n_1441) );
INVx2_ASAP7_75t_SL g1492 ( .A(n_391), .Y(n_1492) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_L g469 ( .A(n_393), .Y(n_469) );
AND2x4_ASAP7_75t_L g476 ( .A(n_393), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g486 ( .A(n_393), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_393), .Y(n_495) );
AND2x2_ASAP7_75t_L g517 ( .A(n_393), .B(n_394), .Y(n_517) );
INVx1_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
INVx2_ASAP7_75t_L g477 ( .A(n_394), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_394), .Y(n_482) );
INVx1_ASAP7_75t_L g855 ( .A(n_394), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_394), .B(n_469), .Y(n_905) );
AND2x4_ASAP7_75t_L g481 ( .A(n_395), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g675 ( .A(n_396), .B(n_485), .Y(n_675) );
OR2x2_ASAP7_75t_L g856 ( .A(n_396), .B(n_485), .Y(n_856) );
XNOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_1140), .Y(n_397) );
XNOR2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_946), .Y(n_398) );
XOR2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_779), .Y(n_399) );
AO22x2_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_649), .B1(n_650), .B2(n_778), .Y(n_400) );
INVx1_ASAP7_75t_L g778 ( .A(n_401), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_568), .Y(n_401) );
INVx1_ASAP7_75t_L g567 ( .A(n_403), .Y(n_567) );
AOI221x1_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_455), .B1(n_461), .B2(n_504), .C(n_507), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_424), .C(n_434), .D(n_451), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_418), .B2(n_419), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_407), .A2(n_419), .B1(n_665), .B2(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_407), .A2(n_419), .B1(n_796), .B2(n_797), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_407), .A2(n_419), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_407), .A2(n_419), .B1(n_453), .B2(n_1056), .C(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_407), .A2(n_419), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AOI22xp5_ASAP7_75t_SL g1351 ( .A1(n_407), .A2(n_426), .B1(n_1352), .B2(n_1353), .Y(n_1351) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
AND2x6_ASAP7_75t_L g430 ( .A(n_408), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g586 ( .A(n_408), .B(n_411), .Y(n_586) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g575 ( .A(n_409), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g421 ( .A(n_410), .Y(n_421) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_410), .Y(n_428) );
AND2x2_ASAP7_75t_L g553 ( .A(n_410), .B(n_458), .Y(n_553) );
INVx2_ASAP7_75t_L g565 ( .A(n_410), .Y(n_565) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_412), .Y(n_541) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_412), .Y(n_557) );
INVx2_ASAP7_75t_L g610 ( .A(n_412), .Y(n_610) );
INVx2_ASAP7_75t_SL g708 ( .A(n_412), .Y(n_708) );
INVx2_ASAP7_75t_L g1124 ( .A(n_412), .Y(n_1124) );
INVx1_ASAP7_75t_L g1203 ( .A(n_412), .Y(n_1203) );
INVx1_ASAP7_75t_L g1382 ( .A(n_412), .Y(n_1382) );
INVx6_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g426 ( .A(n_413), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g772 ( .A(n_413), .Y(n_772) );
BUFx2_ASAP7_75t_L g986 ( .A(n_413), .Y(n_986) );
AND2x2_ASAP7_75t_L g1761 ( .A(n_413), .B(n_1762), .Y(n_1761) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g450 ( .A(n_414), .Y(n_450) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g422 ( .A(n_415), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g441 ( .A(n_415), .B(n_417), .Y(n_441) );
INVx1_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g432 ( .A(n_417), .B(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_419), .A2(n_585), .B1(n_586), .B2(n_587), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_419), .A2(n_586), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx6p67_ASAP7_75t_R g848 ( .A(n_419), .Y(n_848) );
AOI22xp5_ASAP7_75t_SL g964 ( .A1(n_419), .A2(n_586), .B1(n_965), .B2(n_966), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_419), .A2(n_430), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_419), .A2(n_430), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_419), .A2(n_430), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AOI22xp5_ASAP7_75t_L g1395 ( .A1(n_419), .A2(n_430), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1863 ( .A1(n_419), .A2(n_586), .B1(n_1864), .B2(n_1865), .Y(n_1863) );
AND2x6_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
INVx1_ASAP7_75t_L g846 ( .A(n_420), .Y(n_846) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_420), .B(n_767), .Y(n_1355) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x6_ASAP7_75t_L g449 ( .A(n_421), .B(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_422), .Y(n_547) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_422), .Y(n_560) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_422), .Y(n_615) );
INVx2_ASAP7_75t_SL g713 ( .A(n_422), .Y(n_713) );
BUFx2_ASAP7_75t_L g815 ( .A(n_422), .Y(n_815) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_422), .Y(n_872) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_422), .Y(n_939) );
BUFx3_ASAP7_75t_L g994 ( .A(n_422), .Y(n_994) );
BUFx2_ASAP7_75t_L g1272 ( .A(n_422), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1897 ( .A(n_422), .Y(n_1897) );
INVx1_ASAP7_75t_L g582 ( .A(n_423), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_429), .B2(n_430), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_425), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_426), .A2(n_430), .B1(n_589), .B2(n_590), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_426), .A2(n_430), .B1(n_662), .B2(n_663), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_426), .A2(n_430), .B1(n_453), .B2(n_734), .C(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_426), .A2(n_430), .B1(n_793), .B2(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_426), .A2(n_430), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx4_ASAP7_75t_L g884 ( .A(n_426), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_426), .A2(n_430), .B1(n_962), .B2(n_971), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_426), .A2(n_430), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_426), .A2(n_430), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_426), .A2(n_430), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
AOI22xp5_ASAP7_75t_SL g1392 ( .A1(n_426), .A2(n_586), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1866 ( .A1(n_426), .A2(n_430), .B1(n_1867), .B2(n_1868), .Y(n_1866) );
AND2x4_ASAP7_75t_L g444 ( .A(n_427), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_SL g740 ( .A(n_427), .B(n_445), .Y(n_740) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx4_ASAP7_75t_L g885 ( .A(n_430), .Y(n_885) );
INVx2_ASAP7_75t_L g549 ( .A(n_431), .Y(n_549) );
INVx1_ASAP7_75t_L g703 ( .A(n_431), .Y(n_703) );
INVx1_ASAP7_75t_L g715 ( .A(n_431), .Y(n_715) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_431), .Y(n_774) );
BUFx6f_ASAP7_75t_L g940 ( .A(n_431), .Y(n_940) );
INVx1_ASAP7_75t_L g1040 ( .A(n_431), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g619 ( .A(n_432), .Y(n_619) );
INVx1_ASAP7_75t_L g817 ( .A(n_432), .Y(n_817) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_432), .Y(n_824) );
INVx1_ASAP7_75t_L g990 ( .A(n_432), .Y(n_990) );
INVx1_ASAP7_75t_L g581 ( .A(n_433), .Y(n_581) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_442), .B2(n_443), .C1(n_448), .C2(n_449), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g800 ( .A1(n_438), .A2(n_449), .B1(n_740), .B2(n_789), .C1(n_790), .C2(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g621 ( .A(n_439), .Y(n_621) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g453 ( .A(n_440), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g658 ( .A(n_440), .Y(n_658) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_440), .Y(n_738) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_440), .Y(n_767) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_441), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g478 ( .A1(n_442), .A2(n_448), .B1(n_479), .B2(n_483), .C1(n_490), .C2(n_491), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g967 ( .A1(n_443), .A2(n_449), .B1(n_958), .B2(n_959), .C1(n_968), .C2(n_969), .Y(n_967) );
AOI222xp33_ASAP7_75t_L g1103 ( .A1(n_443), .A2(n_449), .B1(n_1104), .B2(n_1105), .C1(n_1106), .C2(n_1107), .Y(n_1103) );
BUFx4f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_444), .A2(n_449), .B1(n_656), .B2(n_657), .C1(n_659), .C2(n_660), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_444), .A2(n_449), .B1(n_891), .B2(n_892), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_444), .A2(n_449), .B1(n_958), .B2(n_959), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_444), .A2(n_449), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_444), .A2(n_449), .B1(n_1296), .B2(n_1297), .Y(n_1337) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g576 ( .A(n_446), .Y(n_576) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g1281 ( .A(n_447), .Y(n_1281) );
INVx3_ASAP7_75t_L g583 ( .A(n_449), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g736 ( .A1(n_449), .A2(n_728), .B1(n_731), .B2(n_737), .C1(n_739), .C2(n_740), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_449), .A2(n_575), .B1(n_839), .B2(n_840), .Y(n_838) );
AOI222xp33_ASAP7_75t_L g1020 ( .A1(n_449), .A2(n_558), .B1(n_740), .B2(n_1021), .C1(n_1022), .C2(n_1023), .Y(n_1020) );
AOI222xp33_ASAP7_75t_L g1058 ( .A1(n_449), .A2(n_740), .B1(n_1059), .B2(n_1060), .C1(n_1061), .C2(n_1062), .Y(n_1058) );
AOI222xp33_ASAP7_75t_L g1150 ( .A1(n_449), .A2(n_740), .B1(n_1151), .B2(n_1152), .C1(n_1154), .C2(n_1155), .Y(n_1150) );
AOI222xp33_ASAP7_75t_L g1216 ( .A1(n_449), .A2(n_575), .B1(n_1211), .B2(n_1212), .C1(n_1217), .C2(n_1218), .Y(n_1216) );
AOI222xp33_ASAP7_75t_L g1456 ( .A1(n_449), .A2(n_575), .B1(n_1443), .B2(n_1457), .C1(n_1458), .C2(n_1459), .Y(n_1456) );
AOI222xp33_ASAP7_75t_L g1505 ( .A1(n_449), .A2(n_575), .B1(n_621), .B2(n_1500), .C1(n_1506), .C2(n_1507), .Y(n_1505) );
AOI222xp33_ASAP7_75t_L g1869 ( .A1(n_449), .A2(n_740), .B1(n_987), .B2(n_1870), .C1(n_1871), .C2(n_1872), .Y(n_1869) );
BUFx3_ASAP7_75t_L g1283 ( .A(n_450), .Y(n_1283) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND4xp25_ASAP7_75t_L g963 ( .A(n_452), .B(n_964), .C(n_967), .D(n_970), .Y(n_963) );
NAND4xp25_ASAP7_75t_L g1013 ( .A(n_452), .B(n_1014), .C(n_1017), .D(n_1020), .Y(n_1013) );
NAND4xp25_ASAP7_75t_SL g1096 ( .A(n_452), .B(n_1097), .C(n_1100), .D(n_1103), .Y(n_1096) );
NAND4xp25_ASAP7_75t_L g1350 ( .A(n_452), .B(n_1351), .C(n_1354), .D(n_1358), .Y(n_1350) );
NAND4xp25_ASAP7_75t_L g1391 ( .A(n_452), .B(n_1392), .C(n_1395), .D(n_1398), .Y(n_1391) );
NAND4xp25_ASAP7_75t_SL g1862 ( .A(n_452), .B(n_1863), .C(n_1866), .D(n_1869), .Y(n_1862) );
INVx5_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_453), .B(n_573), .Y(n_572) );
CKINVDCx8_ASAP7_75t_R g654 ( .A(n_453), .Y(n_654) );
NOR2xp33_ASAP7_75t_SL g833 ( .A(n_453), .B(n_834), .Y(n_833) );
AOI221x1_ASAP7_75t_L g570 ( .A1(n_455), .A2(n_504), .B1(n_571), .B2(n_591), .C(n_605), .Y(n_570) );
AOI221x1_ASAP7_75t_L g951 ( .A1(n_455), .A2(n_504), .B1(n_952), .B2(n_963), .C(n_972), .Y(n_951) );
OAI31xp33_ASAP7_75t_L g1004 ( .A1(n_455), .A2(n_1005), .A3(n_1006), .B(n_1009), .Y(n_1004) );
AOI211x1_ASAP7_75t_SL g1095 ( .A1(n_455), .A2(n_1096), .B(n_1108), .C(n_1128), .Y(n_1095) );
OAI31xp33_ASAP7_75t_L g1227 ( .A1(n_455), .A2(n_1228), .A3(n_1229), .B(n_1233), .Y(n_1227) );
AOI211xp5_ASAP7_75t_L g1861 ( .A1(n_455), .A2(n_1862), .B(n_1873), .C(n_1882), .Y(n_1861) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI211x1_ASAP7_75t_SL g652 ( .A1(n_456), .A2(n_653), .B(n_667), .C(n_680), .Y(n_652) );
AOI221x1_ASAP7_75t_L g721 ( .A1(n_456), .A2(n_504), .B1(n_722), .B2(n_735), .C(n_746), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_456), .A2(n_504), .B1(n_783), .B2(n_794), .C(n_802), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g831 ( .A1(n_456), .A2(n_832), .B(n_844), .Y(n_831) );
INVx1_ASAP7_75t_L g1066 ( .A(n_456), .Y(n_1066) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
AND2x4_ASAP7_75t_L g893 ( .A(n_457), .B(n_459), .Y(n_893) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g564 ( .A(n_458), .B(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
OR2x6_ASAP7_75t_L g1262 ( .A(n_460), .B(n_1263), .Y(n_1262) );
NAND4xp25_ASAP7_75t_SL g461 ( .A(n_462), .B(n_478), .C(n_496), .D(n_501), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B1(n_472), .B2(n_473), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_464), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_464), .A2(n_595), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_464), .A2(n_473), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_464), .A2(n_595), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_464), .A2(n_473), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_464), .A2(n_595), .B1(n_954), .B2(n_955), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_464), .A2(n_473), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI22xp5_ASAP7_75t_SL g1090 ( .A1(n_464), .A2(n_473), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_464), .A2(n_595), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g1366 ( .A1(n_464), .A2(n_498), .B1(n_1367), .B2(n_1368), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_464), .A2(n_498), .B1(n_1407), .B2(n_1408), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g1877 ( .A1(n_464), .A2(n_473), .B1(n_1878), .B2(n_1879), .Y(n_1877) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_468), .Y(n_464) );
AND2x4_ASAP7_75t_L g473 ( .A(n_465), .B(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g595 ( .A(n_465), .B(n_474), .Y(n_595) );
INVx1_ASAP7_75t_L g903 ( .A(n_465), .Y(n_903) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g489 ( .A(n_467), .Y(n_489) );
BUFx2_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
INVx1_ASAP7_75t_L g639 ( .A(n_468), .Y(n_639) );
INVx1_ASAP7_75t_L g697 ( .A(n_468), .Y(n_697) );
BUFx6f_ASAP7_75t_L g749 ( .A(n_468), .Y(n_749) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_468), .Y(n_911) );
BUFx6f_ASAP7_75t_L g976 ( .A(n_468), .Y(n_976) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_468), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_468), .B(n_1804), .Y(n_1803) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g1839 ( .A(n_469), .Y(n_1839) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_475), .Y(n_1378) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_476), .Y(n_513) );
INVx1_ASAP7_75t_L g631 ( .A(n_476), .Y(n_631) );
INVx3_ASAP7_75t_L g691 ( .A(n_476), .Y(n_691) );
AND2x4_ASAP7_75t_L g494 ( .A(n_477), .B(n_495), .Y(n_494) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_479), .A2(n_597), .B1(n_598), .B2(n_599), .C1(n_600), .C2(n_601), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g956 ( .A1(n_479), .A2(n_601), .B1(n_756), .B2(n_957), .C1(n_958), .C2(n_959), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_479), .A2(n_483), .B1(n_1231), .B2(n_1232), .Y(n_1237) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g730 ( .A(n_481), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_481), .A2(n_601), .B1(n_636), .B2(n_788), .C1(n_789), .C2(n_790), .Y(n_787) );
AOI222xp33_ASAP7_75t_SL g896 ( .A1(n_481), .A2(n_518), .B1(n_601), .B2(n_891), .C1(n_892), .C2(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g1132 ( .A(n_481), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_481), .A2(n_483), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1464 ( .A1(n_481), .A2(n_483), .B1(n_1458), .B2(n_1459), .Y(n_1464) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_481), .A2(n_483), .B1(n_1506), .B2(n_1507), .Y(n_1511) );
HB1xp67_ASAP7_75t_L g1835 ( .A(n_482), .Y(n_1835) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_483), .A2(n_729), .B1(n_958), .B2(n_959), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_483), .A2(n_729), .B1(n_1154), .B2(n_1155), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_483), .A2(n_729), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
AND2x4_ASAP7_75t_L g601 ( .A(n_484), .B(n_487), .Y(n_601) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g854 ( .A(n_486), .B(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_486), .B(n_855), .Y(n_922) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g503 ( .A(n_488), .Y(n_503) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_489), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g518 ( .A(n_492), .Y(n_518) );
INVx1_ASAP7_75t_L g598 ( .A(n_492), .Y(n_598) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g726 ( .A1(n_493), .A2(n_601), .B1(n_727), .B2(n_728), .C1(n_729), .C2(n_731), .Y(n_726) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g502 ( .A(n_494), .B(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_494), .Y(n_636) );
BUFx3_ASAP7_75t_L g647 ( .A(n_494), .Y(n_647) );
INVx1_ASAP7_75t_L g673 ( .A(n_494), .Y(n_673) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_494), .Y(n_694) );
BUFx3_ASAP7_75t_L g983 ( .A(n_494), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_498), .A2(n_589), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_498), .A2(n_499), .B1(n_662), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_498), .A2(n_499), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_498), .A2(n_604), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_498), .A2(n_604), .B1(n_899), .B2(n_900), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_498), .A2(n_604), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_498), .A2(n_604), .B1(n_1015), .B2(n_1049), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_498), .A2(n_604), .B1(n_1064), .B2(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_498), .A2(n_499), .B1(n_1101), .B2(n_1137), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g1880 ( .A1(n_498), .A2(n_499), .B1(n_1867), .B2(n_1881), .Y(n_1880) );
AOI22xp33_ASAP7_75t_SL g1369 ( .A1(n_499), .A2(n_595), .B1(n_1353), .B2(n_1370), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_499), .A2(n_595), .B1(n_1394), .B2(n_1410), .Y(n_1409) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g604 ( .A(n_500), .Y(n_604) );
NAND4xp25_ASAP7_75t_SL g591 ( .A(n_501), .B(n_592), .C(n_596), .D(n_602), .Y(n_591) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_501), .B(n_723), .C(n_726), .D(n_732), .Y(n_722) );
NAND4xp25_ASAP7_75t_L g783 ( .A(n_501), .B(n_784), .C(n_787), .D(n_791), .Y(n_783) );
NAND3xp33_ASAP7_75t_SL g895 ( .A(n_501), .B(n_896), .C(n_898), .Y(n_895) );
NAND4xp25_ASAP7_75t_L g952 ( .A(n_501), .B(n_953), .C(n_956), .D(n_960), .Y(n_952) );
CKINVDCx11_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_502), .A2(n_671), .B(n_672), .C(n_674), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g850 ( .A(n_502), .B(n_851), .C(n_852), .Y(n_850) );
AOI211xp5_ASAP7_75t_L g1042 ( .A1(n_502), .A2(n_693), .B(n_1043), .C(n_1044), .Y(n_1042) );
AOI211xp5_ASAP7_75t_L g1085 ( .A1(n_502), .A2(n_756), .B(n_1086), .C(n_1087), .Y(n_1085) );
AOI211xp5_ASAP7_75t_L g1129 ( .A1(n_502), .A2(n_756), .B(n_1130), .C(n_1131), .Y(n_1129) );
AOI211xp5_ASAP7_75t_L g1362 ( .A1(n_502), .A2(n_1363), .B(n_1364), .C(n_1365), .Y(n_1362) );
AOI211xp5_ASAP7_75t_L g1403 ( .A1(n_502), .A2(n_685), .B(n_1404), .C(n_1405), .Y(n_1403) );
AOI211xp5_ASAP7_75t_L g1874 ( .A1(n_502), .A2(n_693), .B(n_1875), .C(n_1876), .Y(n_1874) );
OAI21xp5_ASAP7_75t_L g894 ( .A1(n_504), .A2(n_895), .B(n_901), .Y(n_894) );
OAI31xp33_ASAP7_75t_L g997 ( .A1(n_504), .A2(n_998), .A3(n_999), .B(n_1003), .Y(n_997) );
OAI31xp33_ASAP7_75t_L g1160 ( .A1(n_504), .A2(n_1161), .A3(n_1162), .B(n_1166), .Y(n_1160) );
OAI31xp33_ASAP7_75t_SL g1204 ( .A1(n_504), .A2(n_1205), .A3(n_1206), .B(n_1213), .Y(n_1204) );
OAI31xp33_ASAP7_75t_L g1234 ( .A1(n_504), .A2(n_1235), .A3(n_1236), .B(n_1238), .Y(n_1234) );
OAI31xp33_ASAP7_75t_L g1291 ( .A1(n_504), .A2(n_1292), .A3(n_1293), .B(n_1298), .Y(n_1291) );
OAI31xp33_ASAP7_75t_SL g1461 ( .A1(n_504), .A2(n_1462), .A3(n_1463), .B(n_1465), .Y(n_1461) );
OAI31xp33_ASAP7_75t_SL g1508 ( .A1(n_504), .A2(n_1509), .A3(n_1510), .B(n_1512), .Y(n_1508) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
AOI31xp33_ASAP7_75t_L g1041 ( .A1(n_505), .A2(n_1042), .A3(n_1045), .B(n_1048), .Y(n_1041) );
AOI31xp33_ASAP7_75t_SL g1084 ( .A1(n_505), .A2(n_1085), .A3(n_1088), .B(n_1090), .Y(n_1084) );
AOI31xp33_ASAP7_75t_L g1128 ( .A1(n_505), .A2(n_1129), .A3(n_1133), .B(n_1136), .Y(n_1128) );
AOI31xp33_ASAP7_75t_L g1873 ( .A1(n_505), .A2(n_1874), .A3(n_1877), .B(n_1880), .Y(n_1873) );
AND2x4_ASAP7_75t_L g563 ( .A(n_506), .B(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_L g716 ( .A(n_506), .B(n_564), .Y(n_716) );
AND2x4_ASAP7_75t_L g1760 ( .A(n_506), .B(n_1761), .Y(n_1760) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_508), .B(n_524), .C(n_538), .D(n_554), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .C(n_519), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g527 ( .A(n_513), .Y(n_527) );
INVx2_ASAP7_75t_SL g913 ( .A(n_513), .Y(n_913) );
BUFx3_ASAP7_75t_L g1117 ( .A(n_513), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1111 ( .A(n_515), .Y(n_1111) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_SL g531 ( .A(n_516), .Y(n_531) );
INVx2_ASAP7_75t_SL g634 ( .A(n_516), .Y(n_634) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_517), .Y(n_755) );
AOI33xp33_ASAP7_75t_L g1109 ( .A1(n_519), .A2(n_867), .A3(n_1110), .B1(n_1114), .B2(n_1115), .B3(n_1118), .Y(n_1109) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI33xp33_ASAP7_75t_L g626 ( .A1(n_521), .A2(n_532), .A3(n_627), .B1(n_632), .B2(n_637), .B3(n_643), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_521), .B(n_748), .C(n_752), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_521), .B(n_804), .C(n_806), .Y(n_803) );
BUFx3_ASAP7_75t_L g930 ( .A(n_521), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g974 ( .A(n_521), .B(n_975), .C(n_977), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_521), .B(n_1026), .C(n_1027), .Y(n_1025) );
NAND3xp33_ASAP7_75t_L g1168 ( .A(n_521), .B(n_1169), .C(n_1172), .Y(n_1168) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_521), .B(n_1189), .C(n_1191), .Y(n_1188) );
NAND3xp33_ASAP7_75t_L g1372 ( .A(n_521), .B(n_1373), .C(n_1374), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1412 ( .A(n_521), .B(n_1413), .C(n_1414), .Y(n_1412) );
NAND3xp33_ASAP7_75t_L g1883 ( .A(n_521), .B(n_1884), .C(n_1885), .Y(n_1883) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
OR2x6_ASAP7_75t_L g551 ( .A(n_522), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g624 ( .A(n_522), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g683 ( .A(n_522), .B(n_523), .Y(n_683) );
AND2x2_ASAP7_75t_L g762 ( .A(n_522), .B(n_763), .Y(n_762) );
OR2x2_ASAP7_75t_L g932 ( .A(n_522), .B(n_552), .Y(n_932) );
INVx2_ASAP7_75t_L g1766 ( .A(n_522), .Y(n_1766) );
INVx1_ASAP7_75t_L g1816 ( .A(n_523), .Y(n_1816) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .C(n_532), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g1817 ( .A1(n_527), .A2(n_1434), .B1(n_1818), .B2(n_1819), .Y(n_1817) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g644 ( .A(n_531), .Y(n_644) );
AOI33xp33_ASAP7_75t_L g681 ( .A1(n_532), .A2(n_682), .A3(n_684), .B1(n_687), .B2(n_692), .B3(n_695), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_532), .B(n_808), .C(n_811), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g1076 ( .A(n_532), .B(n_1077), .C(n_1080), .Y(n_1076) );
NAND3xp33_ASAP7_75t_L g1173 ( .A(n_532), .B(n_1174), .C(n_1175), .Y(n_1173) );
NAND3xp33_ASAP7_75t_L g1886 ( .A(n_532), .B(n_1887), .C(n_1890), .Y(n_1886) );
INVx5_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx6_ASAP7_75t_L g867 ( .A(n_533), .Y(n_867) );
OR2x6_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g1777 ( .A(n_534), .B(n_1762), .Y(n_1777) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g1845 ( .A(n_535), .B(n_1846), .Y(n_1845) );
INVx2_ASAP7_75t_L g763 ( .A(n_536), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .C(n_550), .Y(n_538) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g766 ( .A(n_541), .Y(n_766) );
INVx1_ASAP7_75t_L g875 ( .A(n_541), .Y(n_875) );
BUFx4f_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g558 ( .A(n_543), .Y(n_558) );
INVx2_ASAP7_75t_SL g612 ( .A(n_543), .Y(n_612) );
INVx1_ASAP7_75t_L g710 ( .A(n_543), .Y(n_710) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_543), .Y(n_987) );
INVx1_ASAP7_75t_L g1153 ( .A(n_543), .Y(n_1153) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g822 ( .A(n_547), .Y(n_822) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g561 ( .A(n_549), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g1484 ( .A1(n_549), .A2(n_1485), .B1(n_1486), .B2(n_1487), .Y(n_1484) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g700 ( .A(n_551), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_551), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_551), .A2(n_1264), .B1(n_1301), .B2(n_1305), .Y(n_1300) );
OAI22xp5_ASAP7_75t_SL g1778 ( .A1(n_551), .A2(n_1264), .B1(n_1779), .B2(n_1787), .Y(n_1778) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g625 ( .A(n_553), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .C(n_562), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_562), .B(n_820), .C(n_821), .Y(n_819) );
AOI33xp33_ASAP7_75t_L g1119 ( .A1(n_562), .A2(n_818), .A3(n_1120), .B1(n_1121), .B2(n_1122), .B3(n_1125), .Y(n_1119) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx4f_ASAP7_75t_L g607 ( .A(n_563), .Y(n_607) );
INVx4_ASAP7_75t_L g941 ( .A(n_563), .Y(n_941) );
AND2x4_ASAP7_75t_L g1762 ( .A(n_565), .B(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_584), .C(n_588), .Y(n_571) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g1401 ( .A(n_575), .Y(n_1401) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_579), .Y(n_1007) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g837 ( .A(n_580), .Y(n_837) );
BUFx2_ASAP7_75t_L g889 ( .A(n_580), .Y(n_889) );
INVx2_ASAP7_75t_L g937 ( .A(n_580), .Y(n_937) );
BUFx4f_ASAP7_75t_L g944 ( .A(n_580), .Y(n_944) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
OR2x2_ASAP7_75t_L g847 ( .A(n_581), .B(n_582), .Y(n_847) );
INVx5_ASAP7_75t_SL g906 ( .A(n_595), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_626), .Y(n_605) );
AOI33xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .A3(n_613), .B1(n_620), .B2(n_622), .B3(n_623), .Y(n_606) );
AOI33xp33_ASAP7_75t_L g868 ( .A1(n_607), .A2(n_700), .A3(n_869), .B1(n_874), .B2(n_876), .B3(n_877), .Y(n_868) );
NAND3xp33_ASAP7_75t_L g1068 ( .A(n_607), .B(n_1069), .C(n_1070), .Y(n_1068) );
CKINVDCx5p33_ASAP7_75t_R g1264 ( .A(n_607), .Y(n_1264) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g873 ( .A(n_612), .Y(n_873) );
INVx1_ASAP7_75t_L g1179 ( .A(n_612), .Y(n_1179) );
INVx1_ASAP7_75t_L g1457 ( .A(n_612), .Y(n_1457) );
BUFx4f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1472 ( .A(n_615), .Y(n_1472) );
BUFx2_ASAP7_75t_L g1785 ( .A(n_615), .Y(n_1785) );
INVx1_ASAP7_75t_L g1852 ( .A(n_615), .Y(n_1852) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g1071 ( .A(n_617), .Y(n_1071) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_618), .Y(n_1311) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1127 ( .A(n_619), .Y(n_1127) );
NAND3xp33_ASAP7_75t_L g764 ( .A(n_623), .B(n_765), .C(n_768), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_623), .B(n_985), .C(n_988), .Y(n_984) );
NAND3xp33_ASAP7_75t_L g1032 ( .A(n_623), .B(n_1033), .C(n_1035), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g1177 ( .A(n_623), .B(n_1178), .C(n_1180), .Y(n_1177) );
NAND3xp33_ASAP7_75t_L g1197 ( .A(n_623), .B(n_1198), .C(n_1199), .Y(n_1197) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_623), .B(n_1381), .C(n_1383), .Y(n_1380) );
NAND3xp33_ASAP7_75t_L g1418 ( .A(n_623), .B(n_1419), .C(n_1420), .Y(n_1418) );
NAND3xp33_ASAP7_75t_L g1891 ( .A(n_623), .B(n_1892), .C(n_1893), .Y(n_1891) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_SL g1445 ( .A1(n_624), .A2(n_941), .B1(n_1446), .B2(n_1449), .Y(n_1445) );
INVx1_ASAP7_75t_L g1829 ( .A(n_628), .Y(n_1829) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g1806 ( .A(n_630), .B(n_1807), .Y(n_1806) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g642 ( .A(n_631), .Y(n_642) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_634), .B(n_1768), .Y(n_1767) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g686 ( .A(n_636), .Y(n_686) );
BUFx2_ASAP7_75t_L g866 ( .A(n_636), .Y(n_866) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g810 ( .A(n_642), .Y(n_810) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g862 ( .A(n_646), .Y(n_862) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_647), .Y(n_756) );
AND2x4_ASAP7_75t_L g1823 ( .A(n_647), .B(n_1807), .Y(n_1823) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_719), .B1(n_720), .B2(n_777), .Y(n_650) );
INVx1_ASAP7_75t_L g777 ( .A(n_651), .Y(n_777) );
INVx1_ASAP7_75t_L g718 ( .A(n_652), .Y(n_718) );
NAND4xp25_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .C(n_661), .D(n_664), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g794 ( .A(n_654), .B(n_795), .C(n_798), .D(n_800), .Y(n_794) );
NAND3xp33_ASAP7_75t_SL g1149 ( .A(n_654), .B(n_1150), .C(n_1156), .Y(n_1149) );
NAND3xp33_ASAP7_75t_SL g1215 ( .A(n_654), .B(n_1216), .C(n_1219), .Y(n_1215) );
NAND2xp5_ASAP7_75t_SL g1455 ( .A(n_654), .B(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_SL g1504 ( .A(n_654), .B(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g1775 ( .A(n_658), .Y(n_1775) );
AOI31xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .A3(n_676), .B(n_679), .Y(n_667) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AO21x1_ASAP7_75t_SL g849 ( .A1(n_679), .A2(n_850), .B(n_857), .Y(n_849) );
AOI31xp33_ASAP7_75t_L g1361 ( .A1(n_679), .A2(n_1362), .A3(n_1366), .B(n_1369), .Y(n_1361) );
AOI31xp33_ASAP7_75t_L g1402 ( .A1(n_679), .A2(n_1403), .A3(n_1406), .B(n_1409), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_699), .Y(n_680) );
BUFx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI33xp33_ASAP7_75t_L g860 ( .A1(n_683), .A2(n_861), .A3(n_863), .B1(n_864), .B2(n_865), .B3(n_867), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g1081 ( .A(n_683), .B(n_1082), .C(n_1083), .Y(n_1081) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g1176 ( .A(n_686), .Y(n_1176) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g698 ( .A(n_689), .Y(n_698) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g925 ( .A(n_690), .Y(n_925) );
INVx2_ASAP7_75t_L g1171 ( .A(n_690), .Y(n_1171) );
INVx2_ASAP7_75t_L g1889 ( .A(n_690), .Y(n_1889) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_691), .Y(n_751) );
INVx3_ASAP7_75t_L g1079 ( .A(n_691), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g1113 ( .A(n_694), .Y(n_1113) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g759 ( .A(n_697), .Y(n_759) );
INVx1_ASAP7_75t_L g805 ( .A(n_697), .Y(n_805) );
AOI33xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .A3(n_704), .B1(n_705), .B2(n_711), .B3(n_716), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g1075 ( .A(n_703), .Y(n_1075) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g1384 ( .A(n_713), .Y(n_1384) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g1273 ( .A(n_715), .Y(n_1273) );
NAND3xp33_ASAP7_75t_L g769 ( .A(n_716), .B(n_770), .C(n_773), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g991 ( .A(n_716), .B(n_992), .C(n_993), .Y(n_991) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_716), .B(n_1037), .C(n_1038), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g1182 ( .A(n_716), .B(n_1183), .C(n_1184), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1200 ( .A(n_716), .B(n_1201), .C(n_1202), .Y(n_1200) );
NAND3xp33_ASAP7_75t_L g1385 ( .A(n_716), .B(n_1386), .C(n_1387), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g1421 ( .A(n_716), .B(n_1422), .C(n_1423), .Y(n_1421) );
INVx1_ASAP7_75t_L g1488 ( .A(n_716), .Y(n_1488) );
NAND3xp33_ASAP7_75t_L g1894 ( .A(n_716), .B(n_1895), .C(n_1896), .Y(n_1894) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g776 ( .A(n_721), .Y(n_776) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_741), .C(n_743), .Y(n_735) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_757), .C(n_764), .D(n_769), .Y(n_746) );
INVx1_ASAP7_75t_L g1326 ( .A(n_750), .Y(n_1326) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_L g980 ( .A(n_751), .Y(n_980) );
INVx2_ASAP7_75t_SL g1030 ( .A(n_751), .Y(n_1030) );
INVx2_ASAP7_75t_L g1190 ( .A(n_751), .Y(n_1190) );
INVx2_ASAP7_75t_L g1195 ( .A(n_751), .Y(n_1195) );
INVx2_ASAP7_75t_L g1259 ( .A(n_751), .Y(n_1259) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_SL g761 ( .A(n_754), .Y(n_761) );
INVx2_ASAP7_75t_L g1192 ( .A(n_754), .Y(n_1192) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
BUFx2_ASAP7_75t_L g982 ( .A(n_755), .Y(n_982) );
AND2x4_ASAP7_75t_L g1811 ( .A(n_755), .B(n_1804), .Y(n_1811) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .C(n_762), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_762), .B(n_979), .C(n_981), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g1028 ( .A(n_762), .B(n_1029), .C(n_1031), .Y(n_1028) );
NAND3xp33_ASAP7_75t_L g1375 ( .A(n_762), .B(n_1376), .C(n_1379), .Y(n_1375) );
NAND3xp33_ASAP7_75t_L g1415 ( .A(n_762), .B(n_1416), .C(n_1417), .Y(n_1415) );
INVx1_ASAP7_75t_L g1444 ( .A(n_762), .Y(n_1444) );
INVx2_ASAP7_75t_SL g1832 ( .A(n_763), .Y(n_1832) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_767), .Y(n_968) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_767), .Y(n_1105) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g1034 ( .A(n_772), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1557 ( .A1(n_775), .A2(n_1558), .B1(n_1559), .B2(n_1560), .Y(n_1557) );
XNOR2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_827), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g826 ( .A(n_782), .Y(n_826) );
NAND4xp25_ASAP7_75t_SL g802 ( .A(n_803), .B(n_807), .C(n_812), .D(n_819), .Y(n_802) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .C(n_818), .Y(n_812) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g1786 ( .A(n_817), .Y(n_1786) );
NAND3xp33_ASAP7_75t_L g1072 ( .A(n_818), .B(n_1073), .C(n_1074), .Y(n_1072) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx6f_ASAP7_75t_L g1181 ( .A(n_824), .Y(n_1181) );
INVx1_ASAP7_75t_L g1474 ( .A(n_824), .Y(n_1474) );
XOR2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_878), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND4xp25_ASAP7_75t_L g830 ( .A(n_831), .B(n_849), .C(n_860), .D(n_868), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_841), .Y(n_832) );
OAI221xp5_ASAP7_75t_L g1446 ( .A1(n_835), .A2(n_1430), .B1(n_1431), .B2(n_1447), .C(n_1448), .Y(n_1446) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_837), .Y(n_1308) );
OR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx2_ASAP7_75t_L g935 ( .A(n_847), .Y(n_935) );
INVx1_ASAP7_75t_L g1285 ( .A(n_847), .Y(n_1285) );
BUFx2_ASAP7_75t_L g1306 ( .A(n_847), .Y(n_1306) );
INVx1_ASAP7_75t_L g1478 ( .A(n_847), .Y(n_1478) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_853), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_926) );
INVx1_ASAP7_75t_L g1001 ( .A(n_853), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1294 ( .A(n_853), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_853), .A2(n_1491), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
INVx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_854), .Y(n_1164) );
INVx2_ASAP7_75t_L g1209 ( .A(n_854), .Y(n_1209) );
INVx2_ASAP7_75t_L g1331 ( .A(n_854), .Y(n_1331) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_867), .A2(n_908), .B1(n_923), .B2(n_930), .C(n_931), .Y(n_907) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_867), .B(n_1194), .C(n_1196), .Y(n_1193) );
INVx2_ASAP7_75t_L g1252 ( .A(n_867), .Y(n_1252) );
INVx1_ASAP7_75t_L g1333 ( .A(n_867), .Y(n_1333) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
BUFx3_ASAP7_75t_L g1126 ( .A(n_872), .Y(n_1126) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND3x1_ASAP7_75t_L g880 ( .A(n_881), .B(n_894), .C(n_907), .Y(n_880) );
OAI31xp33_ASAP7_75t_SL g881 ( .A1(n_882), .A2(n_883), .A3(n_886), .B(n_893), .Y(n_881) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g1449 ( .A1(n_888), .A2(n_934), .B1(n_1450), .B2(n_1451), .C(n_1452), .Y(n_1449) );
INVx2_ASAP7_75t_SL g888 ( .A(n_889), .Y(n_888) );
AOI211xp5_ASAP7_75t_L g1012 ( .A1(n_893), .A2(n_1013), .B(n_1024), .C(n_1041), .Y(n_1012) );
OAI21xp5_ASAP7_75t_L g1148 ( .A1(n_893), .A2(n_1149), .B(n_1159), .Y(n_1148) );
OAI21xp5_ASAP7_75t_SL g1214 ( .A1(n_893), .A2(n_1215), .B(n_1222), .Y(n_1214) );
OAI31xp33_ASAP7_75t_SL g1334 ( .A1(n_893), .A2(n_1335), .A3(n_1336), .B(n_1338), .Y(n_1334) );
AOI211xp5_ASAP7_75t_L g1349 ( .A1(n_893), .A2(n_1350), .B(n_1361), .C(n_1371), .Y(n_1349) );
AOI211xp5_ASAP7_75t_L g1390 ( .A1(n_893), .A2(n_1391), .B(n_1402), .C(n_1411), .Y(n_1390) );
OAI31xp33_ASAP7_75t_SL g1453 ( .A1(n_893), .A2(n_1454), .A3(n_1455), .B(n_1460), .Y(n_1453) );
OAI31xp33_ASAP7_75t_L g1501 ( .A1(n_893), .A2(n_1502), .A3(n_1503), .B(n_1504), .Y(n_1501) );
OAI221xp5_ASAP7_75t_L g942 ( .A1(n_897), .A2(n_899), .B1(n_934), .B2(n_943), .C(n_945), .Y(n_942) );
OR2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
INVx2_ASAP7_75t_L g1256 ( .A(n_904), .Y(n_1256) );
BUFx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1245 ( .A(n_905), .Y(n_1245) );
INVx1_ASAP7_75t_L g1319 ( .A(n_905), .Y(n_1319) );
INVx3_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_SL g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B1(n_918), .B2(n_919), .Y(n_914) );
INVx3_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g1429 ( .A1(n_921), .A2(n_928), .B1(n_1430), .B2(n_1431), .Y(n_1429) );
OAI22xp33_ASAP7_75t_L g1490 ( .A1(n_921), .A2(n_1476), .B1(n_1479), .B2(n_1491), .Y(n_1490) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OAI22xp33_ASAP7_75t_SL g1432 ( .A1(n_925), .A2(n_1433), .B1(n_1434), .B2(n_1435), .Y(n_1432) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_927), .A2(n_929), .B1(n_934), .B2(n_936), .C(n_938), .Y(n_933) );
OAI22xp33_ASAP7_75t_SL g1248 ( .A1(n_928), .A2(n_1249), .B1(n_1250), .B2(n_1251), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1313 ( .A1(n_928), .A2(n_1302), .B1(n_1303), .B2(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1814 ( .A(n_928), .Y(n_1814) );
OAI22xp5_ASAP7_75t_SL g931 ( .A1(n_932), .A2(n_933), .B1(n_941), .B2(n_942), .Y(n_931) );
OAI33xp33_ASAP7_75t_L g1469 ( .A1(n_932), .A2(n_1470), .A3(n_1475), .B1(n_1481), .B2(n_1484), .B3(n_1488), .Y(n_1469) );
OAI221xp5_ASAP7_75t_L g1787 ( .A1(n_934), .A2(n_1788), .B1(n_1789), .B2(n_1790), .C(n_1791), .Y(n_1787) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g1266 ( .A(n_935), .Y(n_1266) );
INVx2_ASAP7_75t_L g1447 ( .A(n_935), .Y(n_1447) );
INVx1_ASAP7_75t_L g1850 ( .A(n_935), .Y(n_1850) );
BUFx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1269 ( .A(n_937), .Y(n_1269) );
OR2x6_ASAP7_75t_L g1847 ( .A(n_937), .B(n_1845), .Y(n_1847) );
INVx1_ASAP7_75t_L g1485 ( .A(n_939), .Y(n_1485) );
BUFx2_ASAP7_75t_L g1783 ( .A(n_943), .Y(n_1783) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_L g1480 ( .A(n_944), .Y(n_1480) );
INVx1_ASAP7_75t_L g1789 ( .A(n_944), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
XNOR2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_1050), .Y(n_947) );
AO22x2_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_950), .B1(n_1010), .B2(n_1011), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g1003 ( .A(n_953), .Y(n_1003) );
INVx1_ASAP7_75t_L g998 ( .A(n_960), .Y(n_998) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_964), .Y(n_1005) );
INVxp67_ASAP7_75t_L g1009 ( .A(n_970), .Y(n_1009) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_973), .B(n_997), .C(n_1004), .Y(n_996) );
AND4x1_ASAP7_75t_L g973 ( .A(n_974), .B(n_978), .C(n_984), .D(n_991), .Y(n_973) );
INVx1_ASAP7_75t_L g1321 ( .A(n_980), .Y(n_1321) );
BUFx2_ASAP7_75t_L g1364 ( .A(n_983), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_986), .Y(n_1275) );
BUFx2_ASAP7_75t_SL g1060 ( .A(n_987), .Y(n_1060) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_990), .B(n_1845), .Y(n_1844) );
BUFx3_ASAP7_75t_L g1792 ( .A(n_994), .Y(n_1792) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1028), .C(n_1032), .D(n_1036), .Y(n_1024) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1052), .B1(n_1093), .B2(n_1139), .Y(n_1050) );
INVx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NOR3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1067), .C(n_1084), .Y(n_1053) );
AOI31xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1058), .A3(n_1063), .B(n_1066), .Y(n_1054) );
NAND4xp25_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1072), .C(n_1076), .D(n_1081), .Y(n_1067) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1079), .Y(n_1438) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1093), .Y(n_1139) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1095), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1119), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
BUFx3_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
XNOR2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1344), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1224), .B1(n_1342), .B2(n_1343), .Y(n_1144) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1145), .Y(n_1342) );
XOR2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1185), .Y(n_1145) );
NAND3x1_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1160), .C(n_1167), .Y(n_1147) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1153), .Y(n_1218) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1164), .Y(n_1251) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1164), .Y(n_1314) );
AND4x1_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1173), .C(n_1177), .D(n_1182), .Y(n_1167) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
XOR2xp5_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1223), .Y(n_1185) );
NAND3xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1204), .C(n_1214), .Y(n_1186) );
AND4x1_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1193), .C(n_1197), .D(n_1200), .Y(n_1187) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1190), .Y(n_1247) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_1209), .B(n_1769), .Y(n_1820) );
OAI22xp33_ASAP7_75t_L g1548 ( .A1(n_1223), .A2(n_1543), .B1(n_1546), .B2(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1224), .Y(n_1343) );
AOI22xp5_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1288), .B1(n_1289), .B2(n_1341), .Y(n_1224) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1225), .Y(n_1341) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1226), .Y(n_1286) );
NAND3xp33_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1234), .C(n_1239), .Y(n_1226) );
NOR3xp33_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1253), .C(n_1274), .Y(n_1239) );
NOR3xp33_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1248), .C(n_1252), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1243), .B1(n_1246), .B2(n_1247), .Y(n_1241) );
BUFx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1245), .Y(n_1434) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1245), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1262), .B1(n_1264), .B2(n_1265), .Y(n_1253) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_1255), .A2(n_1257), .B1(n_1258), .B2(n_1260), .C(n_1261), .Y(n_1254) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
OAI33xp33_ASAP7_75t_L g1312 ( .A1(n_1262), .A2(n_1313), .A3(n_1315), .B1(n_1322), .B2(n_1327), .B3(n_1333), .Y(n_1312) );
OAI33xp33_ASAP7_75t_L g1428 ( .A1(n_1262), .A2(n_1429), .A3(n_1432), .B1(n_1436), .B2(n_1440), .B3(n_1444), .Y(n_1428) );
OAI33xp33_ASAP7_75t_L g1489 ( .A1(n_1262), .A2(n_1444), .A3(n_1490), .B1(n_1493), .B2(n_1494), .B3(n_1498), .Y(n_1489) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1267), .B1(n_1268), .B2(n_1270), .C(n_1271), .Y(n_1265) );
OAI221xp5_ASAP7_75t_L g1301 ( .A1(n_1266), .A2(n_1268), .B1(n_1302), .B2(n_1303), .C(n_1304), .Y(n_1301) );
OAI21xp33_ASAP7_75t_SL g1276 ( .A1(n_1268), .A2(n_1277), .B(n_1278), .Y(n_1276) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
NAND2x1p5_ASAP7_75t_L g1796 ( .A(n_1280), .B(n_1797), .Y(n_1796) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx2_ASAP7_75t_L g1799 ( .A(n_1283), .Y(n_1799) );
BUFx2_ASAP7_75t_L g1780 ( .A(n_1284), .Y(n_1780) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1290), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1299), .C(n_1334), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1312), .Y(n_1299) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1307), .B1(n_1308), .B2(n_1309), .C(n_1310), .Y(n_1305) );
OAI221xp5_ASAP7_75t_L g1812 ( .A1(n_1314), .A2(n_1781), .B1(n_1782), .B2(n_1813), .C(n_1815), .Y(n_1812) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_1316), .A2(n_1317), .B1(n_1320), .B2(n_1321), .Y(n_1315) );
INVx2_ASAP7_75t_SL g1317 ( .A(n_1318), .Y(n_1317) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1318), .Y(n_1324) );
BUFx3_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1319), .Y(n_1827) );
OAI22xp5_ASAP7_75t_SL g1322 ( .A1(n_1323), .A2(n_1324), .B1(n_1325), .B2(n_1326), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1330), .B1(n_1331), .B2(n_1332), .Y(n_1327) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
OAI22xp33_ASAP7_75t_L g1440 ( .A1(n_1331), .A2(n_1441), .B1(n_1442), .B2(n_1443), .Y(n_1440) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_1340), .A2(n_1543), .B1(n_1566), .B2(n_1567), .Y(n_1565) );
XOR2x2_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1424), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1347), .B1(n_1388), .B2(n_1389), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
XNOR2xp5_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1349), .Y(n_1347) );
AOI21xp5_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1356), .B(n_1357), .Y(n_1354) );
AOI21xp5_ASAP7_75t_L g1398 ( .A1(n_1355), .A2(n_1399), .B(n_1400), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1375), .C(n_1380), .D(n_1385), .Y(n_1371) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NAND4xp25_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1415), .C(n_1418), .D(n_1421), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1466), .B1(n_1513), .B2(n_1514), .Y(n_1424) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1425), .Y(n_1513) );
NAND3xp33_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1453), .C(n_1461), .Y(n_1426) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1445), .Y(n_1427) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_1434), .A2(n_1437), .B1(n_1438), .B2(n_1439), .Y(n_1436) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_1434), .A2(n_1438), .B1(n_1471), .B2(n_1473), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_1438), .A2(n_1495), .B1(n_1496), .B2(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1466), .Y(n_1514) );
NAND3xp33_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1501), .C(n_1508), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1489), .Y(n_1468) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_1471), .A2(n_1472), .B1(n_1473), .B2(n_1474), .Y(n_1470) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_1476), .A2(n_1477), .B1(n_1479), .B2(n_1480), .Y(n_1475) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_1477), .A2(n_1480), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
INVx2_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
OAI21xp33_ASAP7_75t_L g1515 ( .A1(n_1516), .A2(n_1749), .B(n_1751), .Y(n_1515) );
NOR2x1_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1684), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1607), .Y(n_1517) );
A2O1A1Ixp33_ASAP7_75t_SL g1518 ( .A1(n_1519), .A2(n_1550), .B(n_1568), .C(n_1599), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1519), .B(n_1597), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1519), .B(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1519), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1539), .Y(n_1519) );
INVx2_ASAP7_75t_L g1584 ( .A(n_1520), .Y(n_1584) );
BUFx3_ASAP7_75t_L g1624 ( .A(n_1520), .Y(n_1624) );
OR2x2_ASAP7_75t_L g1672 ( .A(n_1520), .B(n_1620), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1520), .B(n_1676), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1520), .B(n_1640), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1520), .B(n_1602), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1533), .Y(n_1520) );
AND2x4_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1528), .Y(n_1522) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
OR2x2_ASAP7_75t_L g1544 ( .A(n_1524), .B(n_1529), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1527), .Y(n_1524) );
HB1xp67_ASAP7_75t_L g1904 ( .A(n_1525), .Y(n_1904) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1527), .Y(n_1536) );
AND2x4_ASAP7_75t_L g1530 ( .A(n_1528), .B(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1529), .B(n_1532), .Y(n_1546) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1534), .Y(n_1554) );
BUFx3_ASAP7_75t_L g1750 ( .A(n_1534), .Y(n_1750) );
AND2x4_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1537), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1535), .B(n_1537), .Y(n_1576) );
HB1xp67_ASAP7_75t_L g1905 ( .A(n_1535), .Y(n_1905) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
AND2x4_ASAP7_75t_L g1538 ( .A(n_1536), .B(n_1537), .Y(n_1538) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1538), .Y(n_1556) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1539), .B(n_1584), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1539), .B(n_1629), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1539), .B(n_1649), .Y(n_1648) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1539), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1547), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1540), .B(n_1591), .Y(n_1590) );
INVx2_ASAP7_75t_L g1603 ( .A(n_1540), .Y(n_1603) );
OAI22xp5_ASAP7_75t_L g1541 ( .A1(n_1542), .A2(n_1543), .B1(n_1545), .B2(n_1546), .Y(n_1541) );
BUFx3_ASAP7_75t_L g1559 ( .A(n_1543), .Y(n_1559) );
BUFx6f_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1546), .Y(n_1561) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_1546), .Y(n_1567) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1547), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1547), .B(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1547), .Y(n_1676) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
AOI211xp5_ASAP7_75t_SL g1674 ( .A1(n_1551), .A2(n_1597), .B(n_1675), .C(n_1677), .Y(n_1674) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1562), .Y(n_1551) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1552), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1552), .B(n_1563), .Y(n_1667) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1552), .B(n_1562), .Y(n_1673) );
BUFx3_ASAP7_75t_L g1691 ( .A(n_1552), .Y(n_1691) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx2_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
OAI211xp5_ASAP7_75t_L g1679 ( .A1(n_1562), .A2(n_1680), .B(n_1682), .C(n_1683), .Y(n_1679) );
OAI31xp33_ASAP7_75t_L g1726 ( .A1(n_1562), .A2(n_1631), .A3(n_1727), .B(n_1728), .Y(n_1726) );
NOR3xp33_ASAP7_75t_L g1745 ( .A(n_1562), .B(n_1677), .C(n_1687), .Y(n_1745) );
INVx2_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1563), .B(n_1604), .Y(n_1649) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1563), .Y(n_1664) );
INVx2_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx2_ASAP7_75t_SL g1613 ( .A(n_1564), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1564), .B(n_1606), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1564), .B(n_1580), .Y(n_1725) );
AOI22xp5_ASAP7_75t_L g1568 ( .A1(n_1569), .A2(n_1578), .B1(n_1592), .B2(n_1593), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1621 ( .A(n_1569), .B(n_1618), .Y(n_1621) );
O2A1O1Ixp33_ASAP7_75t_L g1661 ( .A1(n_1569), .A2(n_1618), .B(n_1662), .C(n_1665), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1574), .Y(n_1569) );
INVx1_ASAP7_75t_SL g1570 ( .A(n_1571), .Y(n_1570) );
CKINVDCx5p33_ASAP7_75t_R g1581 ( .A(n_1571), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1571), .B(n_1574), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1605 ( .A(n_1571), .B(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1571), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1571), .B(n_1618), .Y(n_1626) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1571), .Y(n_1678) );
OR2x2_ASAP7_75t_L g1687 ( .A(n_1571), .B(n_1587), .Y(n_1687) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1571), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1571), .B(n_1616), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
CKINVDCx5p33_ASAP7_75t_R g1592 ( .A(n_1574), .Y(n_1592) );
CKINVDCx6p67_ASAP7_75t_R g1606 ( .A(n_1574), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1574), .B(n_1613), .Y(n_1612) );
OAI32xp33_ASAP7_75t_L g1715 ( .A1(n_1574), .A2(n_1653), .A3(n_1691), .B1(n_1716), .B2(n_1717), .Y(n_1715) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1574), .B(n_1650), .Y(n_1717) );
OR2x6_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1577), .Y(n_1574) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
NOR2xp33_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1582), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1580), .B(n_1613), .Y(n_1647) );
NAND3xp33_ASAP7_75t_L g1660 ( .A(n_1580), .B(n_1628), .C(n_1637), .Y(n_1660) );
INVx3_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1581), .B(n_1595), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1581), .B(n_1606), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1581), .B(n_1637), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1692 ( .A(n_1581), .B(n_1693), .Y(n_1692) );
OAI211xp5_ASAP7_75t_L g1686 ( .A1(n_1582), .A2(n_1687), .B(n_1688), .C(n_1689), .Y(n_1686) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1585), .Y(n_1583) );
OR2x2_ASAP7_75t_L g1600 ( .A(n_1584), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1584), .B(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1584), .B(n_1676), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1584), .B(n_1640), .Y(n_1701) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1590), .Y(n_1586) );
INVx3_ASAP7_75t_L g1597 ( .A(n_1587), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1587), .B(n_1602), .Y(n_1609) );
INVx4_ASAP7_75t_L g1618 ( .A(n_1587), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1587), .B(n_1624), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1587), .B(n_1640), .Y(n_1639) );
NAND3xp33_ASAP7_75t_L g1666 ( .A(n_1587), .B(n_1605), .C(n_1667), .Y(n_1666) );
NOR2xp67_ASAP7_75t_SL g1740 ( .A(n_1587), .B(n_1623), .Y(n_1740) );
AND2x4_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1589), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1590), .B(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1590), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1590), .B(n_1618), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1590), .B(n_1629), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1591), .B(n_1603), .Y(n_1640) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
OAI21xp5_ASAP7_75t_SL g1706 ( .A1(n_1594), .A2(n_1707), .B(n_1718), .Y(n_1706) );
O2A1O1Ixp33_ASAP7_75t_L g1719 ( .A1(n_1595), .A2(n_1720), .B(n_1721), .C(n_1722), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1598), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1596), .B(n_1681), .Y(n_1695) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1597), .B(n_1602), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g1643 ( .A(n_1597), .B(n_1644), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_1597), .B(n_1701), .Y(n_1700) );
AOI21xp5_ASAP7_75t_L g1599 ( .A1(n_1600), .A2(n_1604), .B(n_1605), .Y(n_1599) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1600), .Y(n_1636) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1601), .Y(n_1716) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1602), .Y(n_1655) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1603), .B(n_1624), .Y(n_1623) );
INVx2_ASAP7_75t_L g1645 ( .A(n_1603), .Y(n_1645) );
NOR2xp33_ASAP7_75t_L g1658 ( .A(n_1603), .B(n_1624), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1604), .B(n_1714), .Y(n_1713) );
AOI211xp5_ASAP7_75t_L g1615 ( .A1(n_1605), .A2(n_1616), .B(n_1619), .C(n_1622), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1605), .B(n_1628), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1605), .B(n_1709), .Y(n_1708) );
AND2x4_ASAP7_75t_SL g1637 ( .A(n_1606), .B(n_1613), .Y(n_1637) );
NOR2xp33_ASAP7_75t_L g1689 ( .A(n_1606), .B(n_1690), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1606), .B(n_1691), .Y(n_1698) );
OR2x2_ASAP7_75t_L g1736 ( .A(n_1606), .B(n_1613), .Y(n_1736) );
O2A1O1Ixp33_ASAP7_75t_L g1607 ( .A1(n_1608), .A2(n_1630), .B(n_1650), .C(n_1651), .Y(n_1607) );
OAI211xp5_ASAP7_75t_SL g1608 ( .A1(n_1609), .A2(n_1610), .B(n_1615), .C(n_1627), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1693 ( .A(n_1609), .B(n_1624), .Y(n_1693) );
AOI21xp5_ASAP7_75t_L g1746 ( .A1(n_1609), .A2(n_1647), .B(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1612), .B(n_1614), .Y(n_1611) );
INVx2_ASAP7_75t_L g1668 ( .A(n_1612), .Y(n_1668) );
OAI221xp5_ASAP7_75t_L g1723 ( .A1(n_1616), .A2(n_1647), .B1(n_1724), .B2(n_1725), .C(n_1726), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1617), .B(n_1640), .Y(n_1669) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1618), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1621), .Y(n_1683) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1625), .Y(n_1622) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1624), .B(n_1645), .Y(n_1644) );
OR2x2_ASAP7_75t_L g1654 ( .A(n_1624), .B(n_1655), .Y(n_1654) );
OR2x2_ASAP7_75t_L g1681 ( .A(n_1624), .B(n_1676), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1624), .B(n_1705), .Y(n_1748) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1629), .Y(n_1727) );
OAI211xp5_ASAP7_75t_L g1630 ( .A1(n_1631), .A2(n_1633), .B(n_1635), .C(n_1648), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
OAI21xp5_ASAP7_75t_L g1703 ( .A1(n_1632), .A2(n_1704), .B(n_1705), .Y(n_1703) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
AOI222xp33_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1637), .B1(n_1638), .B2(n_1641), .C1(n_1643), .C2(n_1646), .Y(n_1635) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1637), .Y(n_1743) );
A2O1A1Ixp33_ASAP7_75t_L g1730 ( .A1(n_1638), .A2(n_1691), .B(n_1731), .C(n_1735), .Y(n_1730) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1640), .Y(n_1677) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
OAI22xp33_ASAP7_75t_L g1665 ( .A1(n_1645), .A2(n_1666), .B1(n_1668), .B2(n_1669), .Y(n_1665) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
O2A1O1Ixp33_ASAP7_75t_SL g1652 ( .A1(n_1649), .A2(n_1653), .B(n_1656), .C(n_1659), .Y(n_1652) );
NAND4xp25_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1661), .C(n_1670), .D(n_1679), .Y(n_1651) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1658), .Y(n_1656) );
INVxp67_ASAP7_75t_SL g1659 ( .A(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
OAI211xp5_ASAP7_75t_L g1738 ( .A1(n_1668), .A2(n_1739), .B(n_1741), .C(n_1744), .Y(n_1738) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1669), .Y(n_1724) );
A2O1A1Ixp33_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1673), .B(n_1674), .C(n_1678), .Y(n_1670) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1672), .B(n_1710), .Y(n_1709) );
INVxp67_ASAP7_75t_L g1718 ( .A(n_1673), .Y(n_1718) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1677), .B(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1678), .Y(n_1732) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
OAI211xp5_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1706), .B(n_1719), .C(n_1737), .Y(n_1684) );
O2A1O1Ixp33_ASAP7_75t_SL g1685 ( .A1(n_1686), .A2(n_1692), .B(n_1694), .C(n_1699), .Y(n_1685) );
INVx2_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
OAI21xp5_ASAP7_75t_L g1737 ( .A1(n_1691), .A2(n_1738), .B(n_1746), .Y(n_1737) );
OAI21xp33_ASAP7_75t_L g1694 ( .A1(n_1695), .A2(n_1696), .B(n_1697), .Y(n_1694) );
NOR2xp33_ASAP7_75t_L g1742 ( .A(n_1695), .B(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1696), .Y(n_1702) );
INVxp33_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
OAI21xp5_ASAP7_75t_L g1699 ( .A1(n_1700), .A2(n_1702), .B(n_1703), .Y(n_1699) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1701), .Y(n_1704) );
NAND4xp25_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1712), .C(n_1713), .D(n_1715), .Y(n_1707) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1712), .Y(n_1720) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1730), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1733), .Y(n_1731) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
INVxp67_ASAP7_75t_SL g1741 ( .A(n_1742), .Y(n_1741) );
INVxp67_ASAP7_75t_SL g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
CKINVDCx5p33_ASAP7_75t_R g1749 ( .A(n_1750), .Y(n_1749) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
XNOR2xp5_ASAP7_75t_L g1754 ( .A(n_1755), .B(n_1756), .Y(n_1754) );
AND4x1_ASAP7_75t_L g1756 ( .A(n_1757), .B(n_1772), .C(n_1800), .D(n_1842), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1758), .B(n_1759), .Y(n_1757) );
OR2x6_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1765), .Y(n_1759) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
NOR2xp67_ASAP7_75t_L g1765 ( .A(n_1766), .B(n_1767), .Y(n_1765) );
INVx2_ASAP7_75t_L g1841 ( .A(n_1766), .Y(n_1841) );
AND2x2_ASAP7_75t_L g1834 ( .A(n_1768), .B(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
OR2x6_ASAP7_75t_L g1838 ( .A(n_1769), .B(n_1839), .Y(n_1838) );
INVx2_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
NOR3xp33_ASAP7_75t_SL g1772 ( .A(n_1773), .B(n_1778), .C(n_1793), .Y(n_1772) );
BUFx2_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1776), .Y(n_1774) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
INVx2_ASAP7_75t_SL g1797 ( .A(n_1777), .Y(n_1797) );
OR2x2_ASAP7_75t_L g1798 ( .A(n_1777), .B(n_1799), .Y(n_1798) );
OAI221xp5_ASAP7_75t_L g1779 ( .A1(n_1780), .A2(n_1781), .B1(n_1782), .B2(n_1783), .C(n_1784), .Y(n_1779) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
OAI31xp33_ASAP7_75t_L g1800 ( .A1(n_1801), .A2(n_1809), .A3(n_1821), .B(n_1841), .Y(n_1800) );
INVx3_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVx2_ASAP7_75t_L g1808 ( .A(n_1804), .Y(n_1808) );
INVx3_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
CKINVDCx6p67_ASAP7_75t_R g1810 ( .A(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
INVx2_ASAP7_75t_L g1815 ( .A(n_1816), .Y(n_1815) );
INVx8_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
OAI221xp5_ASAP7_75t_L g1824 ( .A1(n_1825), .A2(n_1828), .B1(n_1829), .B2(n_1830), .C(n_1831), .Y(n_1824) );
INVx2_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
INVx2_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
AOI22xp33_ASAP7_75t_L g1833 ( .A1(n_1834), .A2(n_1836), .B1(n_1837), .B2(n_1840), .Y(n_1833) );
CKINVDCx11_ASAP7_75t_R g1837 ( .A(n_1838), .Y(n_1837) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1848), .Y(n_1842) );
OR2x2_ASAP7_75t_L g1849 ( .A(n_1845), .B(n_1850), .Y(n_1849) );
OR2x2_ASAP7_75t_L g1851 ( .A(n_1845), .B(n_1852), .Y(n_1851) );
BUFx2_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
INVxp67_ASAP7_75t_SL g1855 ( .A(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
HB1xp67_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1861), .Y(n_1860) );
NAND4xp25_ASAP7_75t_L g1882 ( .A(n_1883), .B(n_1886), .C(n_1891), .D(n_1894), .Y(n_1882) );
INVx2_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
INVx1_ASAP7_75t_L g1898 ( .A(n_1899), .Y(n_1898) );
CKINVDCx5p33_ASAP7_75t_R g1899 ( .A(n_1900), .Y(n_1899) );
A2O1A1Ixp33_ASAP7_75t_L g1902 ( .A1(n_1901), .A2(n_1903), .B(n_1905), .C(n_1906), .Y(n_1902) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1904), .Y(n_1903) );
endmodule