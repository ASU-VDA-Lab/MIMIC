module fake_jpeg_6501_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_15),
.B(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_19),
.B(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_13),
.B1(n_12),
.B2(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_24),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_28),
.B(n_10),
.Y(n_30)
);

OAI31xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_9),
.A3(n_7),
.B(n_8),
.Y(n_28)
);

AOI21x1_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_9),
.B(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

OAI31xp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_9),
.A3(n_12),
.B(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_12),
.B1(n_3),
.B2(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);


endmodule