module fake_jpeg_17832_n_98 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_1),
.Y(n_65)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_62),
.Y(n_69)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.C(n_52),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_53),
.B1(n_48),
.B2(n_40),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_71),
.B1(n_7),
.B2(n_8),
.Y(n_75)
);

OA22x2_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_49),
.B1(n_46),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_43),
.B1(n_14),
.B2(n_16),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_82),
.B(n_77),
.CON(n_85),
.SN(n_85)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_63),
.Y(n_87)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_88),
.B1(n_69),
.B2(n_67),
.C(n_76),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_74),
.B1(n_76),
.B2(n_18),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_37),
.C(n_17),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_10),
.B1(n_21),
.B2(n_23),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_25),
.C(n_26),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_27),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_30),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_31),
.C(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_34),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_36),
.Y(n_98)
);


endmodule