module real_jpeg_4588_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_300;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_299;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_244;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_1),
.A2(n_119),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_1),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_2),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_2),
.A2(n_61),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_94),
.B(n_97),
.C(n_100),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_61),
.B1(n_118),
.B2(n_123),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_61),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_72),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_2),
.B(n_130),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_156),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_2),
.B(n_247),
.C(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_2),
.B(n_244),
.C(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_26),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_26),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_26),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_6),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_7),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_10),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_205),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_203),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_174),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_126),
.C(n_167),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_17),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_65),
.B2(n_91),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_19),
.B(n_219),
.C(n_224),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_19),
.A2(n_20),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_20),
.B(n_65),
.C(n_92),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_30),
.B1(n_45),
.B2(n_57),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_30),
.B1(n_45),
.B2(n_57),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_22),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_72)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_24),
.Y(n_271)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_30),
.B(n_45),
.Y(n_199)
);

NAND2x1_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_45),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B1(n_40),
.B2(n_42),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_41),
.Y(n_276)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_45),
.Y(n_259)
);

AOI22x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_47),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_48),
.Y(n_155)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_49),
.Y(n_143)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_49),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_57),
.Y(n_198)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_86),
.B2(n_90),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_66),
.A2(n_71),
.B1(n_86),
.B2(n_90),
.Y(n_173)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_78)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_75),
.Y(n_98)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_93),
.A2(n_101),
.B1(n_102),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_93),
.Y(n_217)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_101),
.A2(n_102),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_102),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_102),
.B(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_102),
.B(n_191),
.C(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_111),
.B1(n_115),
.B2(n_117),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_103),
.A2(n_111),
.B1(n_117),
.B2(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_114),
.Y(n_236)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_117),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_139),
.B1(n_140),
.B2(n_166),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_140),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_131),
.B(n_136),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_181),
.B1(n_182),
.B2(n_189),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_137),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_139),
.A2(n_140),
.B1(n_243),
.B2(n_252),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_139),
.B(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_139),
.A2(n_140),
.B1(n_168),
.B2(n_213),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_139),
.B(n_213),
.C(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_161),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_173),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_169),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_172),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_200),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_194),
.B2(n_195),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_190),
.B2(n_191),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_190),
.A2(n_191),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_190),
.A2(n_191),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_191),
.B(n_287),
.C(n_289),
.Y(n_297)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_226),
.B(n_302),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_207),
.B(n_209),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.C(n_218),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_210),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_242),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_219),
.A2(n_220),
.B1(n_224),
.B2(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_296),
.B(n_301),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_284),
.B(n_295),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_263),
.B(n_283),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_254),
.B(n_262),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_241),
.B(n_253),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_238),
.B(n_240),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_265),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_282),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_277),
.B2(n_281),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_294),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_289),
.B1(n_290),
.B2(n_293),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);


endmodule