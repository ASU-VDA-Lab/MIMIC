module real_jpeg_3862_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_56),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_0),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_0),
.B(n_182),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_0),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_0),
.B(n_165),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_0),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_0),
.B(n_380),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_1),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_1),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_2),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_3),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_4),
.Y(n_182)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_5),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_5),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_7),
.Y(n_540)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_8),
.Y(n_380)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_10),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_10),
.B(n_38),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_10),
.B(n_108),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_10),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_10),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_10),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_10),
.B(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_10),
.B(n_421),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_11),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_54),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_12),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_12),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_12),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_12),
.B(n_187),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_12),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_13),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_13),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_13),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_13),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_13),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_14),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_14),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_14),
.B(n_56),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_14),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_14),
.B(n_222),
.Y(n_415)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_16),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_17),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_17),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_17),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_17),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_17),
.B(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_17),
.B(n_280),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_17),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_18),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_18),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_18),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_18),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_18),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_18),
.B(n_185),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_18),
.B(n_424),
.Y(n_423)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_538),
.B(n_541),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_49),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_30),
.B1(n_40),
.B2(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_27),
.B(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_53),
.C(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_34),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_34),
.Y(n_200)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_34),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_72),
.C(n_74),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_50),
.B(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_62),
.C(n_64),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_51),
.B(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_60),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_59),
.B1(n_67),
.B2(n_120),
.Y(n_124)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_57),
.Y(n_212)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_57),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_65),
.C(n_67),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_64),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_65),
.A2(n_66),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_67),
.A2(n_115),
.B1(n_116),
.B2(n_120),
.Y(n_514)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_70),
.Y(n_352)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_70),
.Y(n_364)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_71),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_131),
.B(n_537),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_128),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_79),
.B(n_128),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_125),
.C(n_126),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_80),
.A2(n_81),
.B1(n_533),
.B2(n_534),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_110),
.C(n_121),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_82),
.A2(n_83),
.B1(n_516),
.B2(n_518),
.Y(n_515)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_89),
.C(n_95),
.Y(n_125)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_88),
.Y(n_222)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_88),
.Y(n_273)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_94),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_106),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_96),
.B(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_100),
.A2(n_101),
.B1(n_106),
.B2(n_107),
.Y(n_507)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_110),
.A2(n_121),
.B1(n_122),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_110),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_120),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_111),
.B(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_115),
.A2(n_116),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_116),
.B(n_198),
.C(n_202),
.Y(n_511)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_118),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_125),
.B(n_126),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_531),
.B(n_536),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_500),
.B(n_528),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_305),
.B(n_499),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_253),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_135),
.B(n_253),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_195),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_136),
.B(n_196),
.C(n_231),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_166),
.C(n_179),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_137),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.C(n_154),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_138),
.B(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_142),
.C(n_143),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_144),
.A2(n_145),
.B1(n_154),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_146),
.B(n_153),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_148),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_154),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_164),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_158),
.B(n_163),
.C(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_164),
.B1(n_202),
.B2(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_163),
.B(n_202),
.C(n_235),
.Y(n_246)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_166),
.B(n_179),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_178),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_167)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_173),
.A2(n_177),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_176),
.C(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_173),
.B(n_245),
.C(n_249),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.C(n_191),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_186),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_181),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_186),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_188),
.B(n_191),
.Y(n_284)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_190),
.Y(n_327)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_231),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_197),
.B(n_209),
.C(n_230),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_200),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_220),
.B1(n_229),
.B2(n_230),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_216),
.Y(n_241)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_219),
.Y(n_395)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_243),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_232),
.B(n_244),
.C(n_251),
.Y(n_523)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.C(n_240),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_255),
.B(n_258),
.Y(n_495)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_260),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_282),
.C(n_285),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_262),
.B(n_488),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_270),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_263),
.A2(n_264),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_266),
.B(n_270),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_277),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_443)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_277),
.B(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_278),
.B(n_379),
.Y(n_378)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_285),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_299),
.C(n_303),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_287),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_288),
.B(n_455),
.Y(n_454)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_291),
.Y(n_456)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_299),
.B(n_303),
.Y(n_477)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_493),
.B(n_498),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_480),
.B(n_492),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_462),
.B(n_479),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_436),
.B(n_461),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_405),
.B(n_435),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_371),
.B(n_404),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_354),
.B(n_370),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_334),
.B(n_353),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_328),
.B(n_333),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_326),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_326),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_321),
.Y(n_335)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_336),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_345),
.B2(n_346),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_348),
.C(n_350),
.Y(n_369)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_342),
.Y(n_360)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_369),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_369),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_361),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_360),
.C(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_359),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_361),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_390),
.C(n_391),
.Y(n_389)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_364),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_374),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_388),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_389),
.C(n_392),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_378),
.C(n_381),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx4_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_387),
.Y(n_381)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_383),
.B(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_401),
.C(n_402),
.Y(n_433)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_396)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_397),
.Y(n_402)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_401),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_434),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_434),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_417),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_416),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_416),
.C(n_460),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_450),
.C(n_451),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_415),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_417),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_427),
.C(n_432),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_422),
.C(n_423),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_432),
.B2(n_433),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_430),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_459),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_459),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_448),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_440),
.C(n_448),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_442),
.B1(n_444),
.B2(n_445),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_471),
.C(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_453),
.C(n_458),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_478),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_478),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_469),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_468),
.C(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_474),
.C(n_476),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_490),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_490),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_487),
.C(n_497),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_496),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_524),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g528 ( 
.A1(n_501),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_520),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_520),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_509),
.B2(n_519),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_510),
.C(n_515),
.Y(n_535)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.C(n_508),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_522),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_508),
.Y(n_522)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_509),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_515),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_521),
.C(n_523),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_521),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_512),
.CI(n_513),
.CON(n_510),
.SN(n_510)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_516),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_525),
.B(n_527),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_527),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_535),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx13_ASAP7_75t_L g543 ( 
.A(n_540),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_544),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);


endmodule