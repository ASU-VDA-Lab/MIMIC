module fake_netlist_1_12492_n_733 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_733);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_733;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_52), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_51), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_64), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_77), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_0), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_68), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_63), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_41), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_83), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_47), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_23), .Y(n_120) );
BUFx5_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_58), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_20), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_11), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_69), .Y(n_128) );
INVx1_ASAP7_75t_SL g129 ( .A(n_84), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_26), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
BUFx10_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_11), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_25), .Y(n_135) );
INVx1_ASAP7_75t_SL g136 ( .A(n_39), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_18), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_10), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
INVxp33_ASAP7_75t_SL g140 ( .A(n_33), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_1), .Y(n_141) );
CKINVDCx14_ASAP7_75t_R g142 ( .A(n_85), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_0), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_50), .Y(n_145) );
INVx1_ASAP7_75t_SL g146 ( .A(n_18), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_44), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_92), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_24), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_7), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_3), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_87), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_121), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_110), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_108), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_109), .B(n_1), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_125), .B(n_2), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_122), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_137), .B(n_2), .Y(n_166) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_109), .A2(n_55), .B(n_105), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_148), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_116), .A2(n_131), .B(n_118), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_148), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_116), .B(n_57), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_114), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_143), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_163), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
NAND3xp33_ASAP7_75t_L g178 ( .A(n_159), .B(n_119), .C(n_128), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_155), .B(n_123), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_171), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_171), .Y(n_182) );
AND3x2_ASAP7_75t_L g183 ( .A(n_158), .B(n_111), .C(n_151), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
BUFx4f_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_154), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_157), .B(n_126), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_157), .B(n_146), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_155), .B(n_142), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
INVx6_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_155), .B(n_142), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_194), .B(n_155), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_193), .A2(n_154), .B1(n_168), .B2(n_170), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_194), .B(n_161), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_193), .A2(n_172), .B1(n_166), .B2(n_168), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_171), .B1(n_140), .B2(n_138), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_185), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_185), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_194), .B(n_112), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_177), .A2(n_167), .B(n_127), .C(n_134), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_199), .B(n_113), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_145), .B(n_130), .Y(n_212) );
NOR2xp67_ASAP7_75t_L g213 ( .A(n_188), .B(n_160), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_191), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_199), .B(n_115), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_193), .A2(n_172), .B1(n_173), .B2(n_141), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_199), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_179), .B(n_117), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_190), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_188), .B(n_120), .Y(n_220) );
NOR2x2_ASAP7_75t_L g221 ( .A(n_183), .B(n_132), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_188), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_178), .A2(n_133), .B1(n_150), .B2(n_152), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_179), .B(n_124), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_189), .B(n_144), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_196), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_196), .B(n_138), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g228 ( .A(n_196), .B(n_171), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_189), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_183), .B(n_129), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_177), .B(n_184), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_186), .A2(n_135), .B(n_136), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_177), .A2(n_138), .B1(n_149), .B2(n_153), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_177), .B(n_122), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_180), .B(n_121), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_226), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_229), .B(n_184), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_203), .B(n_184), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_231), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_214), .B(n_184), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_217), .B(n_192), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_210), .B(n_192), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_225), .B(n_192), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_226), .Y(n_244) );
OAI221xp5_ASAP7_75t_L g245 ( .A1(n_204), .A2(n_192), .B1(n_190), .B2(n_174), .C(n_175), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_216), .B(n_196), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_222), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_201), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_226), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_207), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_207), .B(n_180), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_206), .A2(n_186), .B(n_195), .Y(n_252) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_223), .A2(n_176), .B(n_175), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_206), .B(n_180), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_222), .B(n_196), .Y(n_255) );
AOI22x1_ASAP7_75t_L g256 ( .A1(n_212), .A2(n_180), .B1(n_182), .B2(n_195), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_186), .B(n_195), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_219), .A2(n_195), .B(n_182), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_202), .A2(n_174), .B1(n_176), .B2(n_181), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_226), .Y(n_260) );
NAND2x1_ASAP7_75t_L g261 ( .A(n_226), .B(n_182), .Y(n_261) );
NOR3xp33_ASAP7_75t_L g262 ( .A(n_230), .B(n_182), .C(n_181), .Y(n_262) );
INVx3_ASAP7_75t_SL g263 ( .A(n_221), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_235), .A2(n_195), .B(n_198), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_208), .A2(n_195), .B1(n_171), .B2(n_121), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_209), .A2(n_195), .B(n_160), .C(n_147), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_228), .A2(n_200), .B(n_198), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_266), .A2(n_234), .A3(n_232), .B(n_233), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_258), .A2(n_211), .B(n_215), .Y(n_269) );
NAND3xp33_ASAP7_75t_SL g270 ( .A(n_247), .B(n_224), .C(n_218), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_259), .B(n_220), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_227), .B(n_213), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_243), .A2(n_205), .B(n_213), .C(n_227), .Y(n_273) );
NOR4xp25_ASAP7_75t_L g274 ( .A(n_266), .B(n_160), .C(n_221), .D(n_121), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_257), .A2(n_171), .B(n_198), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_240), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_251), .A2(n_200), .B(n_197), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_242), .B(n_12), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_248), .A2(n_139), .B(n_147), .C(n_164), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_265), .B(n_164), .C(n_156), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_250), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_251), .A2(n_200), .B(n_197), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g283 ( .A1(n_247), .A2(n_139), .B1(n_147), .B2(n_14), .Y(n_283) );
AO32x2_ASAP7_75t_L g284 ( .A1(n_259), .A2(n_164), .A3(n_165), .B1(n_139), .B2(n_147), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_263), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_246), .B(n_12), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_264), .A2(n_197), .B(n_187), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_256), .A2(n_187), .B(n_139), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_245), .A2(n_187), .B(n_165), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_263), .B(n_13), .Y(n_290) );
INVx6_ASAP7_75t_L g291 ( .A(n_236), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_249), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_276), .A2(n_241), .B1(n_237), .B2(n_239), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_278), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_269), .A2(n_250), .B(n_254), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_281), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_278), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_276), .B(n_241), .Y(n_298) );
AO31x2_ASAP7_75t_L g299 ( .A1(n_279), .A2(n_238), .A3(n_267), .B(n_255), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_274), .A2(n_262), .B(n_253), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_275), .A2(n_254), .B(n_249), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_285), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_271), .A2(n_244), .B1(n_260), .B2(n_236), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_286), .B(n_244), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_270), .B(n_244), .Y(n_306) );
INVx6_ASAP7_75t_L g307 ( .A(n_292), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_290), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_288), .A2(n_261), .B(n_260), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_275), .A2(n_260), .B(n_236), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_272), .A2(n_260), .B(n_236), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_273), .A2(n_165), .B(n_164), .C(n_15), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_274), .A2(n_13), .B(n_14), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_305), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_314), .A2(n_289), .B(n_280), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_296), .B(n_284), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_309), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_310), .B(n_268), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_311), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_300), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_313), .A2(n_280), .B(n_287), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_294), .B(n_283), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_312), .A2(n_282), .B(n_277), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_293), .B(n_268), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_303), .B(n_165), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_299), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_299), .Y(n_340) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_268), .B(n_291), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_332), .B(n_301), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_325), .B(n_299), .Y(n_344) );
INVx4_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_325), .B(n_308), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_318), .B(n_164), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_315), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_322), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_318), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_319), .A2(n_298), .B1(n_307), .B2(n_302), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_340), .B(n_165), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_332), .B(n_15), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_326), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_16), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_339), .A2(n_291), .B(n_17), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_339), .B(n_16), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_321), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_339), .B(n_17), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_319), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_331), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_337), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_333), .B(n_19), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_333), .B(n_335), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_322), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_333), .B(n_19), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_368), .B(n_333), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_368), .B(n_333), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_347), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_346), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_371), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_369), .B(n_335), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_346), .B(n_302), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_371), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_380), .B(n_323), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_369), .B(n_335), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_380), .B(n_323), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_359), .B(n_335), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_345), .B(n_335), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_378), .B(n_329), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_379), .B(n_329), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_350), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_349), .B(n_334), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_349), .B(n_334), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_324), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_374), .B(n_324), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_344), .B(n_324), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_360), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_345), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_371), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_363), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_358), .B(n_334), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_324), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_367), .B(n_327), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_362), .A2(n_324), .B1(n_320), .B2(n_336), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_360), .B(n_341), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_358), .B(n_327), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_353), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
OAI21x1_ASAP7_75t_L g431 ( .A1(n_342), .A2(n_330), .B(n_336), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_367), .B(n_338), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_352), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_345), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_352), .Y(n_435) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_345), .B(n_322), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_360), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_362), .B(n_338), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_362), .B(n_338), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_373), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_373), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_375), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_344), .B(n_338), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_375), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_353), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_367), .B(n_338), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_354), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_354), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_382), .B(n_341), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_385), .B(n_338), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_381), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_418), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_418), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_415), .B(n_343), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_387), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_390), .B(n_381), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_387), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_392), .B(n_381), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
OAI211xp5_ASAP7_75t_L g462 ( .A1(n_406), .A2(n_355), .B(n_376), .C(n_385), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_385), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_434), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_389), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_437), .B(n_376), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_415), .B(n_343), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_395), .B(n_355), .C(n_366), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_423), .B(n_343), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_423), .B(n_343), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_405), .B(n_386), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_452), .B(n_376), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_386), .B(n_376), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_404), .B(n_382), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_434), .B(n_384), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_412), .B(n_343), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_412), .B(n_384), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_397), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_388), .B(n_348), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_393), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_393), .B(n_348), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_388), .B(n_348), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_389), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_391), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_413), .B(n_343), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_396), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_424), .B(n_366), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_394), .B(n_372), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_400), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_407), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_394), .B(n_372), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_403), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
INVx4_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_396), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_435), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_399), .B(n_372), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_413), .B(n_356), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_419), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_444), .B(n_356), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_448), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_444), .B(n_356), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_399), .B(n_361), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_426), .B(n_361), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_426), .B(n_361), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_448), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_449), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_426), .B(n_364), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_398), .B(n_372), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_450), .B(n_364), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_401), .B(n_342), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_449), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_419), .B(n_342), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_422), .B(n_342), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_430), .B(n_351), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_407), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_450), .B(n_364), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_450), .B(n_383), .Y(n_522) );
INVx3_ASAP7_75t_L g523 ( .A(n_436), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_440), .B(n_441), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_408), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_408), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_442), .B(n_383), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_443), .B(n_338), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_414), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_445), .B(n_338), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_414), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_422), .B(n_383), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_438), .B(n_370), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_428), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_417), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_432), .B(n_370), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_473), .B(n_409), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_486), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_453), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_534), .B(n_409), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_464), .B(n_438), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_460), .Y(n_543) );
OAI32xp33_ASAP7_75t_L g544 ( .A1(n_454), .A2(n_402), .A3(n_410), .B1(n_439), .B2(n_428), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_466), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_470), .A2(n_469), .B(n_455), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_455), .B(n_439), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_524), .B(n_410), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_462), .A2(n_425), .B1(n_447), .B2(n_451), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_469), .B(n_402), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_453), .A2(n_446), .B(n_429), .C(n_427), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_498), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_497), .B(n_351), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_529), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_491), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_482), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_494), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_503), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_461), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_465), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_524), .B(n_417), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_529), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_482), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_471), .B(n_427), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_488), .B(n_307), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_497), .B(n_357), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_471), .B(n_429), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_472), .B(n_446), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_499), .B(n_341), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_479), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_489), .B(n_370), .Y(n_577) );
NAND2xp33_ASAP7_75t_L g578 ( .A(n_483), .B(n_322), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_500), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_505), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_479), .B(n_357), .Y(n_581) );
NOR2xp33_ASAP7_75t_SL g582 ( .A(n_483), .B(n_357), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_502), .B(n_365), .Y(n_583) );
OAI32xp33_ASAP7_75t_L g584 ( .A1(n_468), .A2(n_357), .A3(n_351), .B1(n_365), .B2(n_320), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_472), .B(n_351), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_479), .B(n_365), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_R g587 ( .A1(n_478), .A2(n_307), .B(n_320), .C(n_431), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_523), .B(n_320), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_478), .B(n_431), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_514), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_510), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_507), .B(n_320), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_507), .B(n_320), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_511), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_504), .B(n_328), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_516), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_487), .B(n_330), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_513), .B(n_328), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_487), .B(n_330), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_532), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_504), .B(n_328), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_463), .A2(n_307), .B1(n_328), .B2(n_28), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_328), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_477), .A2(n_328), .B(n_22), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_506), .B(n_21), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_506), .B(n_29), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_527), .B(n_30), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_481), .B(n_31), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_484), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_536), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_521), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_536), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_456), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_474), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_554), .A2(n_475), .B1(n_457), .B2(n_476), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_549), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_554), .A2(n_476), .B1(n_523), .B2(n_508), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_549), .B(n_533), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_545), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_609), .B(n_515), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_556), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_582), .B(n_477), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_546), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_559), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g626 ( .A1(n_538), .A2(n_490), .A3(n_493), .B1(n_501), .B2(n_459), .C1(n_518), .C2(n_530), .Y(n_626) );
OAI211xp5_ASAP7_75t_SL g627 ( .A1(n_547), .A2(n_523), .B(n_528), .C(n_518), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_577), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_610), .B(n_521), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_612), .B(n_519), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_539), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_552), .A2(n_476), .B1(n_477), .B2(n_509), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_543), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_611), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_574), .B(n_600), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_553), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_599), .A2(n_512), .B1(n_508), .B2(n_509), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_601), .B(n_512), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_563), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_597), .A2(n_522), .B1(n_517), .B2(n_526), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_563), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_537), .B(n_540), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_553), .A2(n_522), .B1(n_531), .B2(n_526), .C1(n_525), .C2(n_535), .Y(n_644) );
AOI322xp5_ASAP7_75t_L g645 ( .A1(n_576), .A2(n_535), .A3(n_531), .B1(n_525), .B2(n_520), .C1(n_492), .C2(n_485), .Y(n_645) );
OAI22xp33_ASAP7_75t_SL g646 ( .A1(n_558), .A2(n_520), .B1(n_492), .B2(n_485), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_614), .B(n_458), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_562), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_572), .B(n_590), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_602), .A2(n_467), .B(n_458), .Y(n_650) );
AO22x1_ASAP7_75t_L g651 ( .A1(n_566), .A2(n_467), .B1(n_456), .B2(n_35), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_544), .A2(n_32), .B(n_34), .C(n_37), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_38), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_565), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_573), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_579), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_597), .B(n_106), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_550), .A2(n_40), .B1(n_42), .B2(n_43), .C(n_46), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_580), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_560), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_551), .B(n_48), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_592), .B(n_104), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_591), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_594), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_617), .A2(n_541), .B1(n_542), .B2(n_602), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_661), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_639), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_621), .Y(n_669) );
AOI221x1_ASAP7_75t_L g670 ( .A1(n_627), .A2(n_568), .B1(n_607), .B2(n_596), .C(n_604), .Y(n_670) );
OAI21xp33_ASAP7_75t_SL g671 ( .A1(n_622), .A2(n_587), .B(n_589), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_634), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_636), .B(n_564), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_637), .B(n_548), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g675 ( .A1(n_632), .A2(n_582), .A3(n_578), .B1(n_555), .B2(n_569), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_644), .A2(n_584), .B(n_607), .C(n_608), .Y(n_676) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_652), .B(n_555), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_659), .B(n_606), .C(n_605), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_635), .Y(n_680) );
OA21x2_ASAP7_75t_L g681 ( .A1(n_631), .A2(n_598), .B(n_603), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_616), .B(n_581), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_640), .B(n_567), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_618), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_643), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_615), .A2(n_585), .B1(n_593), .B2(n_570), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_632), .A2(n_569), .B(n_586), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_646), .A2(n_588), .B(n_598), .C(n_575), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_615), .A2(n_571), .B1(n_595), .B2(n_603), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_645), .B(n_575), .C(n_583), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_620), .B(n_588), .Y(n_691) );
A2O1A1O1Ixp25_ASAP7_75t_L g692 ( .A1(n_650), .A2(n_49), .B(n_53), .C(n_54), .D(n_56), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_651), .A2(n_59), .B(n_61), .Y(n_693) );
AOI33xp33_ASAP7_75t_L g694 ( .A1(n_619), .A2(n_62), .A3(n_65), .B1(n_66), .B2(n_67), .B3(n_70), .Y(n_694) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_650), .B(n_71), .Y(n_695) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_657), .B(n_72), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_657), .B(n_73), .C(n_74), .D(n_75), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_626), .A2(n_76), .B(n_78), .C(n_79), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_81), .B1(n_82), .B2(n_86), .C(n_88), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_653), .A2(n_89), .B(n_93), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_648), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_623), .A2(n_94), .B(n_95), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_642), .A2(n_96), .B(n_97), .C(n_99), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_624), .B(n_101), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_662), .B(n_103), .C(n_663), .D(n_625), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_633), .A2(n_654), .B1(n_664), .B2(n_660), .C(n_656), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_655), .A2(n_665), .B1(n_630), .B2(n_629), .C(n_638), .Y(n_707) );
O2A1O1Ixp5_ASAP7_75t_L g708 ( .A1(n_658), .A2(n_647), .B(n_628), .C(n_649), .Y(n_708) );
OA22x2_ASAP7_75t_L g709 ( .A1(n_666), .A2(n_670), .B1(n_689), .B2(n_686), .Y(n_709) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_671), .A2(n_690), .B1(n_680), .B2(n_706), .C1(n_672), .C2(n_707), .Y(n_710) );
OAI21xp33_ASAP7_75t_SL g711 ( .A1(n_675), .A2(n_677), .B(n_695), .Y(n_711) );
O2A1O1Ixp5_ASAP7_75t_L g712 ( .A1(n_708), .A2(n_690), .B(n_687), .C(n_691), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_667), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_701), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_698), .A2(n_688), .B(n_699), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_692), .B(n_676), .C(n_694), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_710), .B(n_684), .Y(n_717) );
AND5x1_ASAP7_75t_L g718 ( .A(n_709), .B(n_696), .C(n_673), .D(n_693), .E(n_679), .Y(n_718) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_711), .B(n_705), .C(n_703), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_712), .B(n_697), .C(n_700), .D(n_702), .Y(n_720) );
OR2x6_ASAP7_75t_L g721 ( .A(n_717), .B(n_713), .Y(n_721) );
NOR2x1p5_ASAP7_75t_L g722 ( .A(n_720), .B(n_716), .Y(n_722) );
NOR2x1p5_ASAP7_75t_L g723 ( .A(n_718), .B(n_714), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_722), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_721), .B(n_719), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_724), .A2(n_723), .B1(n_669), .B2(n_715), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_725), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_727), .B(n_725), .Y(n_728) );
OAI21x1_ASAP7_75t_L g729 ( .A1(n_726), .A2(n_704), .B(n_685), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_728), .A2(n_681), .B1(n_682), .B2(n_678), .Y(n_730) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_730), .A2(n_729), .B(n_728), .Y(n_731) );
OA21x2_ASAP7_75t_L g732 ( .A1(n_731), .A2(n_668), .B(n_674), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_732), .A2(n_683), .B1(n_681), .B2(n_692), .Y(n_733) );
endmodule