module real_jpeg_24796_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_26),
.B1(n_127),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_127),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_127),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_10),
.B1(n_27),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_140),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_140),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_140),
.Y(n_235)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_6),
.A2(n_44),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_6),
.B(n_32),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_136),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_55),
.C(n_60),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_6),
.B(n_68),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_6),
.A2(n_110),
.B1(n_229),
.B2(n_235),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_75),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_75),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_8),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_8),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_9),
.A2(n_27),
.B1(n_63),
.B2(n_137),
.Y(n_296)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_129),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_129),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_129),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_28),
.B1(n_52),
.B2(n_53),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_28),
.B1(n_59),
.B2(n_60),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_14),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_299)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_15),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_86),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_86),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_80),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_20),
.A2(n_21),
.B1(n_76),
.B2(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_48),
.C(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_41),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_24),
.A2(n_31),
.B(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_27),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_41),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_30),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_30),
.A2(n_32),
.B1(n_139),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_30),
.A2(n_32),
.B1(n_147),
.B2(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_30),
.A2(n_271),
.B(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_30),
.A2(n_90),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_31),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_31),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_34),
.B1(n_69),
.B2(n_70),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_33),
.A2(n_37),
.B(n_135),
.C(n_153),
.Y(n_152)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_33),
.B(n_136),
.CON(n_181),
.SN(n_181)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_34),
.B(n_36),
.C(n_137),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_34),
.A2(n_53),
.A3(n_69),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_64),
.B2(n_65),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_76),
.C(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_47),
.A2(n_48),
.B1(n_81),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_58),
.B(n_61),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_62),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_50),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_50),
.A2(n_190),
.B(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_50),
.A2(n_189),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_50),
.A2(n_188),
.B1(n_189),
.B2(n_209),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_50),
.A2(n_189),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_50),
.A2(n_123),
.B(n_265),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_53),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_52),
.B(n_70),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_53),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_58),
.B(n_61),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_58),
.B(n_136),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_59),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_66),
.A2(n_125),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_68),
.B(n_72),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_67),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_68),
.A2(n_72),
.B1(n_172),
.B2(n_181),
.Y(n_186)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_71),
.A2(n_130),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_76),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_76),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_80),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_81),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_83),
.A2(n_125),
.B1(n_130),
.B2(n_299),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_85),
.A2(n_125),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_325),
.A3(n_335),
.B1(n_338),
.B2(n_339),
.C(n_342),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_304),
.B(n_324),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_279),
.B(n_303),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_173),
.B(n_255),
.C(n_278),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_158),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_158),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_143),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_120),
.B1(n_141),
.B2(n_142),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_103),
.B(n_142),
.C(n_143),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_104),
.B(n_109),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_105),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_106),
.B(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B(n_116),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_110),
.A2(n_116),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_110),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_110),
.A2(n_226),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_110),
.A2(n_184),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_111),
.B(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_111),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_113),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_131),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_136),
.B(n_166),
.Y(n_240)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_276)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_159),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_162),
.B(n_164),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_168),
.B1(n_169),
.B2(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_167),
.B(n_220),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_250),
.B(n_254),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_203),
.B(n_249),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_178),
.B(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.C(n_187),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_179),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_187),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_199),
.C(n_202),
.Y(n_251)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_201),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_244),
.B(n_248),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_222),
.B(n_243),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_206),
.B(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_216),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_219),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_242),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_230),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_237),
.B(n_241),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_276),
.B2(n_277),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_267),
.C(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_266),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_266),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_280),
.B(n_281),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_302),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_290),
.B1(n_300),
.B2(n_301),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_301),
.C(n_302),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_286),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_287),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_286),
.A2(n_318),
.B(n_319),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_294),
.C(n_297),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_297),
.B2(n_298),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_305),
.B(n_306),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_322),
.B2(n_323),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_320),
.B2(n_321),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_321),
.C(n_323),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_327),
.C(n_332),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g337 ( 
.A(n_313),
.B(n_327),
.CI(n_332),
.CON(n_337),
.SN(n_337)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_316),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_333),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_336),
.B(n_337),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_337),
.Y(n_340)
);


endmodule