module fake_jpeg_15029_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_14),
.B(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_19),
.B(n_17),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_10),
.B1(n_8),
.B2(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_18),
.B(n_16),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_9),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_16),
.B1(n_10),
.B2(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_40),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_29),
.B(n_9),
.C(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_45),
.B1(n_32),
.B2(n_39),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_32),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_4),
.Y(n_44)
);

AOI322xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_15),
.A3(n_9),
.B1(n_6),
.B2(n_7),
.C1(n_5),
.C2(n_4),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_38),
.B(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_50),
.C(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_53),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI31xp33_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.A3(n_50),
.B(n_48),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_46),
.C(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_5),
.Y(n_60)
);


endmodule