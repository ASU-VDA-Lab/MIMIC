module fake_jpeg_31639_n_543 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_543);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_57),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_71),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_66),
.Y(n_156)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_90),
.Y(n_128)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_15),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_17),
.B(n_14),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_107),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_111),
.B(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_20),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_126),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_20),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_25),
.B1(n_37),
.B2(n_32),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_153),
.B1(n_174),
.B2(n_177),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_107),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g135 ( 
.A(n_55),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_144),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_57),
.B(n_40),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_79),
.A2(n_25),
.B1(n_34),
.B2(n_45),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_70),
.A2(n_51),
.B1(n_27),
.B2(n_48),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_155),
.A2(n_161),
.B1(n_27),
.B2(n_68),
.Y(n_214)
);

BUFx4f_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_159),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_76),
.A2(n_51),
.B1(n_27),
.B2(n_48),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_18),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_72),
.B(n_22),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_97),
.A2(n_34),
.B1(n_48),
.B2(n_45),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_102),
.A2(n_34),
.B1(n_45),
.B2(n_51),
.Y(n_177)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_192),
.Y(n_233)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_92),
.B1(n_104),
.B2(n_101),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_184),
.A2(n_190),
.B1(n_129),
.B2(n_131),
.Y(n_244)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_185),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_86),
.B(n_46),
.C(n_43),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_186),
.A2(n_197),
.B(n_206),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_114),
.A2(n_108),
.B1(n_100),
.B2(n_95),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_187),
.A2(n_223),
.B1(n_36),
.B2(n_29),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_84),
.B1(n_80),
.B2(n_77),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

BUFx4f_ASAP7_75t_SL g239 ( 
.A(n_193),
.Y(n_239)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_22),
.B1(n_40),
.B2(n_52),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

NAND2x1p5_ASAP7_75t_L g197 ( 
.A(n_128),
.B(n_24),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_198),
.Y(n_270)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_139),
.B(n_18),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_218),
.Y(n_250)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_207),
.Y(n_237)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_27),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_115),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_209),
.Y(n_247)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_24),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_212),
.Y(n_261)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_137),
.B(n_24),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_215),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_154),
.B1(n_112),
.B2(n_148),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_138),
.B(n_24),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_150),
.B(n_16),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_220),
.Y(n_266)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_221),
.A2(n_228),
.B1(n_143),
.B2(n_166),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_73),
.B1(n_63),
.B2(n_53),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_150),
.B(n_53),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_50),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_156),
.A2(n_24),
.B(n_46),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_229),
.B(n_31),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_41),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_160),
.Y(n_258)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_130),
.A2(n_174),
.B(n_153),
.C(n_161),
.Y(n_229)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_146),
.Y(n_230)
);

CKINVDCx12_ASAP7_75t_R g274 ( 
.A(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_145),
.B(n_50),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_231),
.B(n_232),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_43),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_229),
.A2(n_142),
.B1(n_162),
.B2(n_158),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_184),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_165),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_236),
.B(n_256),
.CI(n_206),
.CON(n_278),
.SN(n_278)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_240),
.A2(n_213),
.B1(n_201),
.B2(n_203),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_200),
.B(n_113),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_242),
.B(n_267),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_251),
.B1(n_258),
.B2(n_262),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_258),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_191),
.A2(n_175),
.B1(n_122),
.B2(n_112),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

NOR4xp25_ASAP7_75t_SL g256 ( 
.A(n_197),
.B(n_151),
.C(n_133),
.D(n_149),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_120),
.B1(n_123),
.B2(n_221),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_211),
.A2(n_146),
.B1(n_122),
.B2(n_110),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_214),
.B1(n_227),
.B2(n_196),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_205),
.B(n_31),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_183),
.B1(n_180),
.B2(n_188),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_178),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_286),
.C(n_263),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_296),
.B1(n_240),
.B2(n_234),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_279),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_241),
.A2(n_194),
.B1(n_225),
.B2(n_206),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_289),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_251),
.A2(n_224),
.B1(n_218),
.B2(n_198),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_186),
.C(n_181),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_293),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_190),
.B1(n_189),
.B2(n_199),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_292),
.Y(n_323)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_227),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_253),
.B(n_195),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_304),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_255),
.B1(n_272),
.B2(n_257),
.Y(n_313)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_233),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_204),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_244),
.A2(n_226),
.B1(n_179),
.B2(n_209),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_306),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_250),
.B(n_29),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_250),
.B(n_185),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_247),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_308),
.A2(n_298),
.B1(n_278),
.B2(n_304),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_321),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_236),
.B(n_234),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_311),
.A2(n_294),
.B(n_286),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_289),
.B1(n_276),
.B2(n_285),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_261),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_324),
.C(n_325),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_279),
.A2(n_236),
.B1(n_234),
.B2(n_237),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_318),
.A2(n_319),
.B1(n_281),
.B2(n_280),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_238),
.B1(n_264),
.B2(n_271),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_287),
.B(n_273),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_261),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_237),
.C(n_273),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_242),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_333),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_292),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_334),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_335),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_248),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_337),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

AO22x1_ASAP7_75t_SL g340 ( 
.A1(n_332),
.A2(n_278),
.B1(n_305),
.B2(n_283),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_SL g374 ( 
.A1(n_340),
.A2(n_351),
.B(n_357),
.C(n_361),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_359),
.B(n_361),
.Y(n_369)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_343),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_344),
.A2(n_349),
.B1(n_320),
.B2(n_252),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_309),
.B(n_288),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_346),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_332),
.A2(n_301),
.B(n_291),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_347),
.A2(n_329),
.B(n_326),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_318),
.A2(n_278),
.B1(n_294),
.B2(n_300),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_355),
.B1(n_360),
.B2(n_366),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_332),
.A2(n_299),
.B(n_274),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_321),
.B(n_277),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_358),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_317),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_353),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_302),
.B1(n_295),
.B2(n_293),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_311),
.A2(n_274),
.B(n_247),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_335),
.A2(n_277),
.B(n_249),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_308),
.A2(n_238),
.B1(n_284),
.B2(n_257),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_335),
.A2(n_264),
.B(n_239),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_252),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_364),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_320),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_365),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_316),
.A2(n_238),
.B1(n_284),
.B2(n_257),
.Y(n_366)
);

XOR2x2_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_325),
.Y(n_367)
);

A2O1A1O1Ixp25_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_345),
.B(n_364),
.C(n_357),
.D(n_340),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_348),
.C(n_314),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_373),
.C(n_380),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_314),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_392),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_374),
.B(n_376),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_348),
.C(n_310),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_363),
.A2(n_332),
.B(n_329),
.Y(n_376)
);

AOI22x1_ASAP7_75t_L g377 ( 
.A1(n_363),
.A2(n_315),
.B1(n_309),
.B2(n_312),
.Y(n_377)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_310),
.C(n_324),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_324),
.C(n_325),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_381),
.B(n_390),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_363),
.A2(n_319),
.B(n_315),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_382),
.A2(n_362),
.B(n_339),
.Y(n_411)
);

OAI211xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_336),
.B(n_322),
.C(n_337),
.Y(n_385)
);

AOI322xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_334),
.A3(n_330),
.B1(n_323),
.B2(n_343),
.C1(n_265),
.C2(n_239),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_333),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_344),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_388),
.A2(n_356),
.B1(n_358),
.B2(n_350),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_346),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_354),
.B(n_313),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_266),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_395),
.B(n_396),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_312),
.C(n_272),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_408),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_399),
.A2(n_404),
.B1(n_374),
.B2(n_389),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_351),
.B(n_347),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_402),
.A2(n_369),
.B(n_374),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_387),
.A2(n_355),
.B1(n_360),
.B2(n_366),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_410),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_384),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_345),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_417),
.Y(n_445)
);

A2O1A1O1Ixp25_ASAP7_75t_L g410 ( 
.A1(n_367),
.A2(n_357),
.B(n_340),
.C(n_362),
.D(n_344),
.Y(n_410)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_371),
.B(n_340),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_413),
.B(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_266),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_379),
.Y(n_418)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_383),
.A2(n_340),
.B1(n_360),
.B2(n_366),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_419),
.A2(n_290),
.B1(n_327),
.B2(n_246),
.Y(n_442)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_420),
.Y(n_433)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_420),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_422),
.A2(n_424),
.B1(n_425),
.B2(n_391),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_328),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_423),
.B(n_412),
.C(n_413),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_382),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_381),
.B(n_323),
.Y(n_425)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_429),
.C(n_431),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_373),
.C(n_368),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_396),
.C(n_391),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_411),
.B(n_410),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_392),
.C(n_376),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_435),
.C(n_441),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_372),
.C(n_383),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_387),
.B1(n_375),
.B2(n_389),
.Y(n_436)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_438),
.A2(n_414),
.B1(n_219),
.B2(n_239),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_374),
.C(n_270),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_442),
.A2(n_448),
.B1(n_418),
.B2(n_414),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_415),
.C(n_401),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_447),
.C(n_193),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_270),
.C(n_265),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_290),
.B1(n_246),
.B2(n_220),
.Y(n_448)
);

XOR2x2_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_406),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_462),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_407),
.Y(n_451)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_437),
.A2(n_421),
.B1(n_403),
.B2(n_404),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_452),
.A2(n_455),
.B1(n_457),
.B2(n_461),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_442),
.A2(n_403),
.B1(n_424),
.B2(n_416),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_402),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_469),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_459),
.A2(n_9),
.B(n_42),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_460),
.A2(n_465),
.B1(n_443),
.B2(n_446),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_448),
.A2(n_239),
.B1(n_36),
.B2(n_230),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_427),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_440),
.A2(n_36),
.B1(n_230),
.B2(n_193),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_433),
.B1(n_426),
.B2(n_447),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_438),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_467),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_42),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_13),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_462),
.C(n_429),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_477),
.C(n_466),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_454),
.A2(n_433),
.B(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_472),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_475),
.Y(n_494)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_445),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_482),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_444),
.C(n_441),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_481),
.A2(n_471),
.B1(n_460),
.B2(n_465),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_468),
.A2(n_435),
.B1(n_426),
.B2(n_13),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_10),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_483),
.B(n_484),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_10),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_487),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_486),
.B(n_9),
.Y(n_502)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_469),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_458),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_495),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_456),
.C(n_450),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_498),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_467),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_0),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_457),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_42),
.C(n_1),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_500),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_42),
.C(n_1),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_42),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_497),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_473),
.A2(n_472),
.B(n_479),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_0),
.Y(n_507)
);

OA21x2_ASAP7_75t_SL g504 ( 
.A1(n_494),
.A2(n_486),
.B(n_2),
.Y(n_504)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_507),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g509 ( 
.A1(n_491),
.A2(n_0),
.B(n_2),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_509),
.A2(n_3),
.B(n_4),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_511),
.B(n_515),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_502),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_2),
.B(n_3),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_489),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_2),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_492),
.B(n_3),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_517),
.Y(n_523)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_518),
.A2(n_505),
.B1(n_517),
.B2(n_5),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_508),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_524),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_515),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_490),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_525),
.B(n_514),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_506),
.C(n_514),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_530),
.Y(n_536)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_528),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_523),
.A2(n_488),
.B(n_499),
.Y(n_530)
);

AOI21xp33_ASAP7_75t_L g535 ( 
.A1(n_531),
.A2(n_520),
.B(n_526),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_521),
.C(n_518),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_535),
.C(n_529),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_537),
.A2(n_538),
.B(n_534),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_536),
.B(n_531),
.C(n_4),
.Y(n_538)
);

AOI221xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_5),
.B(n_8),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_5),
.Y(n_542)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_8),
.C(n_397),
.Y(n_543)
);


endmodule