module fake_jpeg_6879_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_20),
.B(n_16),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_46),
.B(n_22),
.C(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_13),
.B1(n_22),
.B2(n_15),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_14),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_30),
.B(n_25),
.Y(n_53)
);

FAx1_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_56),
.CI(n_35),
.CON(n_64),
.SN(n_64)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_33),
.B1(n_27),
.B2(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_37),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_58),
.B(n_54),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_68),
.B(n_67),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_56),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_61),
.C(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_89),
.C(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_82),
.B1(n_50),
.B2(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_88),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_50),
.B1(n_64),
.B2(n_56),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_62),
.C(n_56),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_64),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_62),
.A3(n_49),
.B1(n_27),
.B2(n_33),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_52),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_34),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_49),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_73),
.B1(n_59),
.B2(n_39),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_85),
.B1(n_88),
.B2(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_97),
.B1(n_101),
.B2(n_93),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_112),
.B(n_11),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_113),
.B(n_18),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_19),
.B(n_1),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_59),
.B(n_11),
.C(n_10),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_55),
.B1(n_48),
.B2(n_19),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_44),
.C(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_121),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_120),
.B(n_0),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_0),
.B(n_2),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_14),
.B(n_44),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_118),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_122),
.B(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_2),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.C(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_114),
.B(n_3),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_133),
.B(n_6),
.C(n_4),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_55),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_4),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_5),
.Y(n_137)
);


endmodule