module fake_jpeg_7640_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_3),
.B(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_45),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_12),
.Y(n_83)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_61),
.B1(n_27),
.B2(n_32),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_18),
.B1(n_24),
.B2(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_33),
.B1(n_29),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_21),
.B1(n_31),
.B2(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_32),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_27),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_17),
.B1(n_16),
.B2(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_74),
.B1(n_89),
.B2(n_53),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_31),
.B1(n_38),
.B2(n_16),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_78),
.B1(n_48),
.B2(n_46),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_88),
.C(n_26),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_27),
.B1(n_32),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_84),
.B1(n_53),
.B2(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_16),
.B1(n_30),
.B2(n_19),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_51),
.B(n_46),
.Y(n_112)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_22),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_0),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_33),
.B1(n_28),
.B2(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_50),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_112),
.B1(n_114),
.B2(n_73),
.Y(n_129)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_101),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_14),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_105),
.A2(n_111),
.B1(n_118),
.B2(n_108),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_52),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_47),
.B1(n_46),
.B2(n_30),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_26),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_64),
.C(n_88),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_51),
.B1(n_25),
.B2(n_19),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_88),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_106),
.B(n_120),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_63),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_137),
.C(n_143),
.Y(n_177)
);

NOR4xp25_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_82),
.C(n_65),
.D(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_26),
.B(n_25),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_130),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_74),
.B(n_68),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_131),
.B(n_71),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_139),
.B1(n_118),
.B2(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_68),
.B(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_116),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_86),
.B1(n_71),
.B2(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_66),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_86),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_148),
.B(n_3),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_93),
.B1(n_108),
.B2(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_106),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_163),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_157),
.B(n_162),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_120),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_154),
.A2(n_156),
.B(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_170),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_112),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_128),
.B1(n_146),
.B2(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_71),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_117),
.B(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_19),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_90),
.B(n_1),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_10),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_3),
.B(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_171),
.C(n_157),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_193),
.C(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_126),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_126),
.C(n_138),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_138),
.C(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_203),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_122),
.A3(n_142),
.B1(n_135),
.B2(n_8),
.C1(n_9),
.C2(n_11),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_166),
.B1(n_163),
.B2(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_158),
.B1(n_181),
.B2(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_156),
.B(n_154),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_208),
.B(n_198),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_207),
.A2(n_173),
.B(n_162),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_223),
.B(n_230),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_158),
.B1(n_154),
.B2(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_221),
.B1(n_229),
.B2(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_175),
.B1(n_153),
.B2(n_174),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_151),
.C(n_178),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_225),
.C(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_168),
.C(n_153),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_180),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_196),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_172),
.B1(n_164),
.B2(n_176),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_235),
.C(n_237),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_187),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_218),
.B1(n_223),
.B2(n_215),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_250),
.B(n_221),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_232),
.B(n_230),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_246),
.C(n_247),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_191),
.C(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_186),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_217),
.C(n_210),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_249),
.C(n_232),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_191),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_220),
.B(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_257),
.B1(n_259),
.B2(n_263),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_249),
.B(n_235),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_202),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_237),
.C(n_245),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_264),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_238),
.B(n_224),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_234),
.B(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_271),
.B(n_256),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_276),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_253),
.A2(n_229),
.B(n_205),
.C(n_190),
.Y(n_271)
);

OAI321xp33_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_231),
.A3(n_190),
.B1(n_195),
.B2(n_247),
.C(n_233),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_275),
.Y(n_280)
);

OAI321xp33_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_195),
.A3(n_246),
.B1(n_182),
.B2(n_8),
.C(n_9),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_182),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_182),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_277),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_286),
.B1(n_271),
.B2(n_9),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_256),
.B1(n_255),
.B2(n_122),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_271),
.B1(n_5),
.B2(n_6),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.C(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_12),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_280),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_142),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_270),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_293),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_13),
.B(n_14),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_13),
.Y(n_293)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_278),
.B1(n_281),
.B2(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_297),
.B1(n_289),
.B2(n_15),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_291),
.B(n_290),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_301),
.C(n_299),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_295),
.B(n_298),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_283),
.C(n_15),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_4),
.Y(n_305)
);


endmodule