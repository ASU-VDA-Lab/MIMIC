module fake_jpeg_9214_n_27 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_27);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_27;

wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_17;
wire n_25;
wire n_15;

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_11),
.B1(n_1),
.B2(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_2),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_21),
.B1(n_16),
.B2(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_24),
.B1(n_19),
.B2(n_3),
.Y(n_25)
);

OAI21x1_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_22),
.B(n_23),
.Y(n_26)
);

NAND4xp25_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_8),
.C(n_12),
.D(n_13),
.Y(n_27)
);


endmodule