module fake_jpeg_12357_n_431 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_2),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_58),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_40),
.B(n_9),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_95),
.Y(n_117)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_9),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_83),
.B(n_87),
.Y(n_134)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

CKINVDCx9p33_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_26),
.B(n_10),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_88),
.B(n_89),
.Y(n_168)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_92),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_94),
.B(n_100),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_37),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_101),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_104),
.Y(n_126)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_20),
.B(n_0),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_32),
.B(n_11),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_7),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_44),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_35),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_30),
.B1(n_18),
.B2(n_49),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_112),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_49),
.B1(n_18),
.B2(n_54),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_114),
.A2(n_136),
.B1(n_167),
.B2(n_71),
.Y(n_184)
);

INVx2_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_76),
.A2(n_30),
.B1(n_18),
.B2(n_49),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_143),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_59),
.A2(n_29),
.B1(n_50),
.B2(n_34),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_69),
.Y(n_181)
);

CKINVDCx12_ASAP7_75t_R g140 ( 
.A(n_70),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_35),
.B1(n_50),
.B2(n_19),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_34),
.B1(n_29),
.B2(n_22),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_67),
.A2(n_51),
.B1(n_47),
.B2(n_43),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_148),
.A2(n_150),
.B1(n_161),
.B2(n_179),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_80),
.A2(n_22),
.B1(n_19),
.B2(n_51),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_47),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_43),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_27),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_0),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_25),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_68),
.A2(n_24),
.B1(n_45),
.B2(n_14),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_12),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_125),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_108),
.A2(n_12),
.B1(n_15),
.B2(n_45),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_179),
.B1(n_112),
.B2(n_129),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_110),
.A2(n_45),
.B1(n_3),
.B2(n_5),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_74),
.B1(n_98),
.B2(n_92),
.Y(n_180)
);

AOI22x1_ASAP7_75t_L g263 ( 
.A1(n_180),
.A2(n_236),
.B1(n_193),
.B2(n_181),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_181),
.B(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_225),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_183),
.B(n_186),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_184),
.A2(n_214),
.B1(n_223),
.B2(n_225),
.Y(n_269)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_0),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_194),
.C(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_190),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_136),
.A2(n_85),
.B(n_101),
.C(n_37),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_191),
.A2(n_180),
.B(n_222),
.C(n_188),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_3),
.B1(n_37),
.B2(n_169),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_3),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_125),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_197),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_199),
.B(n_220),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_200),
.A2(n_203),
.B1(n_207),
.B2(n_213),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_128),
.A2(n_117),
.B(n_153),
.C(n_134),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_201),
.A2(n_193),
.B(n_204),
.C(n_202),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_142),
.B1(n_141),
.B2(n_124),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_122),
.B1(n_146),
.B2(n_175),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_113),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_138),
.B1(n_164),
.B2(n_147),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_173),
.B1(n_155),
.B2(n_139),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_169),
.A2(n_171),
.B1(n_135),
.B2(n_158),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_218),
.B1(n_232),
.B2(n_227),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_178),
.C(n_135),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_145),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_219),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_171),
.A2(n_157),
.B1(n_158),
.B2(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_119),
.B(n_145),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_119),
.B(n_178),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_236),
.C(n_227),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_174),
.A2(n_173),
.B1(n_144),
.B2(n_147),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

INVx11_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_115),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_230),
.Y(n_256)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.Y(n_262)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_234),
.B(n_232),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_197),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_152),
.B(n_166),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_115),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_276),
.C(n_239),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_246),
.A2(n_254),
.B(n_255),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_229),
.B(n_216),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_278),
.B(n_272),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_256),
.B1(n_237),
.B2(n_271),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_195),
.B1(n_224),
.B2(n_230),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_258),
.B(n_273),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_269),
.B1(n_270),
.B2(n_266),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_184),
.A2(n_183),
.B1(n_189),
.B2(n_191),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_242),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_196),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_277),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_187),
.A2(n_194),
.B(n_181),
.C(n_201),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_221),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_194),
.C(n_185),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_205),
.A2(n_234),
.B(n_233),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_198),
.B(n_228),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_209),
.B1(n_231),
.B2(n_211),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_282),
.A2(n_292),
.B1(n_300),
.B2(n_302),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_284),
.A2(n_285),
.B(n_299),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_267),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_246),
.B1(n_255),
.B2(n_254),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_291),
.B(n_257),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_288),
.B(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_252),
.B(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_251),
.B1(n_261),
.B2(n_238),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_240),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_293),
.B(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_305),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_276),
.C(n_263),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_310),
.C(n_267),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_263),
.B(n_278),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_244),
.B1(n_275),
.B2(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_258),
.A2(n_262),
.B1(n_271),
.B2(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_313),
.B1(n_284),
.B2(n_285),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_237),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_237),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_259),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_288),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_245),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_311),
.B(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_259),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_323),
.C(n_332),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_301),
.B1(n_304),
.B2(n_290),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_273),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_327),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_338),
.B(n_330),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_257),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_330),
.B(n_309),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_311),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_295),
.B(n_266),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_293),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_280),
.C(n_286),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_280),
.C(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_315),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_307),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_297),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_280),
.B1(n_313),
.B2(n_302),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_337),
.A2(n_297),
.B1(n_305),
.B2(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_343),
.B1(n_340),
.B2(n_319),
.Y(n_377)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_329),
.A2(n_296),
.B(n_289),
.C(n_308),
.D(n_281),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_342),
.B(n_357),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_312),
.B1(n_306),
.B2(n_294),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_345),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_336),
.B1(n_328),
.B2(n_318),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_331),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_359),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_324),
.B(n_325),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_354),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_346),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_334),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_355),
.B(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_332),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_329),
.A2(n_319),
.B(n_337),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_361),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_375),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_371),
.A2(n_343),
.B1(n_341),
.B2(n_347),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_333),
.C(n_321),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_334),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_326),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_377),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_326),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_378),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_353),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_383),
.C(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_387),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_357),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_346),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_363),
.A2(n_348),
.B1(n_344),
.B2(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_359),
.C(n_321),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_322),
.B1(n_354),
.B2(n_342),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_391),
.B(n_392),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_366),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_398),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_365),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_396),
.A2(n_402),
.B(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_380),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_400),
.Y(n_407)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_387),
.A2(n_362),
.B(n_371),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_397),
.B(n_374),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_405),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_393),
.A2(n_391),
.B(n_390),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_385),
.B(n_383),
.Y(n_417)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_396),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_408),
.Y(n_412)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_409),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_402),
.A2(n_388),
.B1(n_368),
.B2(n_386),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_410),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_379),
.C(n_401),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_415),
.B(n_417),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_407),
.A2(n_369),
.B1(n_378),
.B2(n_375),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_416),
.A2(n_369),
.B1(n_340),
.B2(n_368),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_406),
.B1(n_373),
.B2(n_370),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_370),
.Y(n_421)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_421),
.A2(n_413),
.B(n_411),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_373),
.B1(n_389),
.B2(n_401),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_422),
.A2(n_415),
.B(n_414),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_424),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_425),
.B(n_420),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_421),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_426),
.C(n_318),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_331),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_320),
.Y(n_431)
);


endmodule