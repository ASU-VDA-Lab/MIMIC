module fake_jpeg_9290_n_235 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_24),
.CON(n_41),
.SN(n_41)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_58),
.B1(n_60),
.B2(n_14),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_20),
.B1(n_26),
.B2(n_24),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_52),
.B1(n_56),
.B2(n_27),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_29),
.B1(n_20),
.B2(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_1),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_21),
.B(n_19),
.C(n_15),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_29),
.B1(n_18),
.B2(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_17),
.B1(n_27),
.B2(n_14),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

FAx1_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_39),
.CI(n_21),
.CON(n_64),
.SN(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_11),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_78),
.B1(n_43),
.B2(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_15),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_59),
.C(n_47),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_44),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_64),
.B(n_73),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_95),
.B(n_97),
.Y(n_110)
);

AOI211xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_49),
.B(n_55),
.C(n_52),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_75),
.B(n_70),
.C(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_96),
.B1(n_53),
.B2(n_77),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_46),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_47),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_43),
.B1(n_53),
.B2(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_55),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_13),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_78),
.B1(n_67),
.B2(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_53),
.B1(n_77),
.B2(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_81),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_131),
.B1(n_134),
.B2(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_134),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_80),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_132),
.C(n_141),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_85),
.B1(n_95),
.B2(n_98),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_110),
.C(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_91),
.B1(n_98),
.B2(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_129),
.B1(n_106),
.B2(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_84),
.B1(n_90),
.B2(n_68),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_9),
.Y(n_161)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_90),
.B1(n_88),
.B2(n_86),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_104),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_39),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_159),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_154),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_107),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_112),
.A3(n_116),
.B1(n_103),
.B2(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_69),
.B1(n_94),
.B2(n_42),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_160),
.Y(n_164)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND5xp2_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_21),
.C(n_19),
.D(n_14),
.E(n_50),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_135),
.B(n_140),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_50),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_10),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_131),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_168),
.C(n_158),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_170),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_176),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_182),
.Y(n_193)
);

BUFx12f_ASAP7_75t_SL g181 ( 
.A(n_172),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_190),
.B(n_65),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_148),
.C(n_146),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_150),
.B1(n_149),
.B2(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_155),
.B1(n_145),
.B2(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_161),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_162),
.C(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_152),
.B1(n_157),
.B2(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_177),
.B1(n_170),
.B2(n_128),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_164),
.B1(n_185),
.B2(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_184),
.C(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_166),
.B1(n_173),
.B2(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_162),
.B(n_9),
.C(n_11),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_65),
.B1(n_42),
.B2(n_4),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_211),
.Y(n_221)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_195),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_213),
.B1(n_201),
.B2(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_217),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_193),
.Y(n_217)
);

OAI321xp33_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_202),
.A3(n_194),
.B1(n_7),
.B2(n_5),
.C(n_6),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_218),
.A2(n_7),
.B(n_8),
.C(n_12),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_208),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_226),
.A3(n_221),
.B1(n_12),
.B2(n_8),
.C1(n_4),
.C2(n_2),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_217),
.C(n_219),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_230),
.B(n_229),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_232),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_234),
.Y(n_235)
);


endmodule