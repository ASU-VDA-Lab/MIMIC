module fake_ibex_1369_n_1026 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1026);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1026;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_972;
wire n_845;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_375;
wire n_317;
wire n_340;
wire n_280;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_580;
wire n_483;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_506;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_951;
wire n_272;
wire n_881;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_955;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_984;
wire n_1000;
wire n_394;
wire n_807;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g186 ( 
.A(n_43),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_13),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_80),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_146),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_34),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_43),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_55),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_137),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVxp67_ASAP7_75t_R g208 ( 
.A(n_79),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_62),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_29),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_97),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_87),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_22),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_1),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_64),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_26),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_154),
.B(n_33),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_95),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_129),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_132),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_94),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_85),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_L g243 ( 
.A(n_48),
.B(n_134),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_140),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_88),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_158),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_66),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_127),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_49),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_143),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_35),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_28),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_116),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_115),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_81),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_125),
.Y(n_260)
);

INVxp33_ASAP7_75t_SL g261 ( 
.A(n_102),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_96),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_32),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_92),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_89),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_126),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_7),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_83),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_111),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_37),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_114),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_82),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_27),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_148),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_84),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_182),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_152),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_14),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_19),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_73),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_106),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_34),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_48),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_173),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_39),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_86),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_170),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_71),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_165),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_98),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_41),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_159),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_153),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_113),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_118),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_15),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_100),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_54),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_42),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_104),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_142),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_59),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_136),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_56),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_14),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_63),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_197),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_197),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_266),
.B(n_0),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_202),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_202),
.B(n_0),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_203),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_203),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_267),
.B(n_1),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_209),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_212),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_189),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_209),
.B(n_2),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_189),
.Y(n_341)
);

CKINVDCx6p67_ASAP7_75t_R g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_210),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_265),
.B(n_67),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_3),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_210),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_261),
.A2(n_314),
.B1(n_305),
.B2(n_192),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_224),
.B(n_3),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_224),
.B(n_4),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_197),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_191),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_270),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_199),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_305),
.B(n_5),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_186),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g359 ( 
.A1(n_196),
.A2(n_90),
.B(n_184),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_200),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_188),
.B(n_8),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_196),
.A2(n_99),
.B(n_180),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_199),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_199),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_261),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_199),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_244),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_190),
.Y(n_369)
);

OAI22x1_ASAP7_75t_R g370 ( 
.A1(n_271),
.A2(n_289),
.B1(n_192),
.B2(n_222),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_205),
.Y(n_371)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_231),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_215),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_195),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_216),
.B(n_12),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_218),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_270),
.B(n_279),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_204),
.B(n_68),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_204),
.B(n_16),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_221),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_279),
.B(n_18),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_221),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_279),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_242),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_208),
.B(n_18),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_226),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_206),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_226),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_272),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_227),
.B(n_240),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_242),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_211),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_299),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_242),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_193),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_272),
.A2(n_105),
.B(n_179),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_213),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_242),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_278),
.A2(n_309),
.B(n_284),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_252),
.B(n_20),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_278),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_254),
.B(n_22),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_255),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_263),
.B(n_23),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_400),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_274),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_207),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_344),
.A2(n_201),
.B1(n_239),
.B2(n_233),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_356),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_198),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_325),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_L g426 ( 
.A(n_325),
.B(n_287),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_380),
.B(n_369),
.Y(n_428)
);

NOR2x1p5_ASAP7_75t_L g429 ( 
.A(n_342),
.B(n_277),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_349),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_282),
.B1(n_285),
.B2(n_281),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_347),
.A2(n_239),
.B1(n_273),
.B2(n_259),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_369),
.B(n_311),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_344),
.A2(n_273),
.B1(n_259),
.B2(n_303),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_386),
.B(n_311),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_326),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_194),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_326),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_327),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_327),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_384),
.B(n_338),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_384),
.B(n_245),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g450 ( 
.A1(n_360),
.A2(n_286),
.B1(n_323),
.B2(n_292),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_374),
.B(n_257),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_333),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_374),
.B(n_269),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_333),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_319),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_342),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_333),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_327),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_328),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_328),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_394),
.B(n_313),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_328),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_373),
.B(n_269),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_388),
.B(n_319),
.Y(n_467)
);

AO21x2_ASAP7_75t_L g468 ( 
.A1(n_329),
.A2(n_217),
.B(n_214),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_337),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_275),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_328),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_328),
.Y(n_472)
);

INVx8_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_393),
.B(n_219),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_345),
.Y(n_475)
);

AND2x2_ASAP7_75t_SL g476 ( 
.A(n_386),
.B(n_324),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_304),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_398),
.B(n_295),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_398),
.B(n_371),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_377),
.B(n_220),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_404),
.B(n_310),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_350),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_312),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_350),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_391),
.B(n_223),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_350),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_339),
.A2(n_317),
.B1(n_318),
.B2(n_320),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_346),
.B(n_225),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_352),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_382),
.Y(n_491)
);

INVx4_ASAP7_75t_SL g492 ( 
.A(n_379),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_352),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_357),
.B(n_228),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_341),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_341),
.B(n_229),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_365),
.A2(n_307),
.B1(n_303),
.B2(n_201),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_351),
.B(n_232),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_331),
.B(n_234),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_354),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_331),
.B(n_235),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_335),
.B(n_283),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_354),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_354),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_381),
.A2(n_324),
.B1(n_193),
.B2(n_230),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_335),
.B(n_297),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_370),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_355),
.B(n_193),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_343),
.B(n_297),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_383),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_343),
.B(n_193),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_387),
.B(n_236),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_387),
.B(n_237),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_389),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_389),
.B(n_390),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_390),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_402),
.B(n_238),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_376),
.B(n_230),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_402),
.B(n_241),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_361),
.B(n_247),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_401),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_363),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx4_ASAP7_75t_SL g527 ( 
.A(n_399),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_436),
.B(n_524),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_513),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_423),
.B(n_302),
.Y(n_530)
);

AO22x1_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_434),
.B1(n_456),
.B2(n_432),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_476),
.A2(n_308),
.B1(n_316),
.B2(n_248),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_308),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_465),
.B(n_470),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_476),
.A2(n_290),
.B1(n_280),
.B2(n_249),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_187),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_250),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_448),
.B(n_253),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_246),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_486),
.B(n_251),
.Y(n_541)
);

AND2x6_ASAP7_75t_SL g542 ( 
.A(n_409),
.B(n_256),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_438),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_409),
.A2(n_300),
.B1(n_258),
.B2(n_260),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_420),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_440),
.B(n_262),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_518),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_442),
.B(n_264),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_478),
.B(n_268),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_410),
.B(n_276),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_409),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_473),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_454),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_498),
.B(n_416),
.C(n_475),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_449),
.B(n_288),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_435),
.B(n_291),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_435),
.B(n_294),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_424),
.B(n_324),
.Y(n_560)
);

CKINVDCx6p67_ASAP7_75t_R g561 ( 
.A(n_479),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_435),
.B(n_306),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_415),
.A2(n_422),
.B1(n_430),
.B2(n_419),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_456),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_435),
.B(n_315),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_406),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_422),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_495),
.Y(n_569)
);

INVxp33_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

OAI22x1_ASAP7_75t_L g571 ( 
.A1(n_429),
.A2(n_509),
.B1(n_439),
.B2(n_450),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_457),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_430),
.A2(n_411),
.B1(n_412),
.B2(n_407),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_322),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_451),
.B(n_359),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_480),
.B(n_503),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_469),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_511),
.B(n_362),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_424),
.B(n_324),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_491),
.A2(n_243),
.B1(n_397),
.B2(n_362),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_491),
.B(n_397),
.Y(n_581)
);

NOR3x1_ASAP7_75t_L g582 ( 
.A(n_484),
.B(n_23),
.C(n_24),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_453),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_441),
.B(n_396),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_444),
.B(n_396),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_399),
.Y(n_587)
);

OA22x2_ASAP7_75t_L g588 ( 
.A1(n_413),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_417),
.B(n_364),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_463),
.B(n_28),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_SL g592 ( 
.A1(n_500),
.A2(n_502),
.B(n_520),
.C(n_516),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_463),
.B(n_31),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_431),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_521),
.B(n_399),
.Y(n_595)
);

NAND2xp33_ASAP7_75t_L g596 ( 
.A(n_458),
.B(n_364),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_418),
.A2(n_395),
.B1(n_392),
.B2(n_385),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_523),
.B(n_367),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_421),
.B(n_367),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_490),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_493),
.Y(n_601)
);

AND2x6_ASAP7_75t_SL g602 ( 
.A(n_489),
.B(n_36),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_428),
.A2(n_395),
.B1(n_392),
.B2(n_385),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

OR2x2_ASAP7_75t_SL g605 ( 
.A(n_450),
.B(n_37),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_473),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_481),
.B(n_395),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_463),
.B(n_38),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_473),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_482),
.B(n_38),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_474),
.B(n_39),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_468),
.B(n_40),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_488),
.B(n_40),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_450),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_425),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_489),
.B(n_47),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_49),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_494),
.B(n_50),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_426),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_512),
.B(n_51),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_528),
.B(n_583),
.Y(n_622)
);

NOR2x1_ASAP7_75t_L g623 ( 
.A(n_545),
.B(n_497),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_613),
.A2(n_488),
.B1(n_517),
.B2(n_519),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_547),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_583),
.B(n_589),
.Y(n_626)
);

AO32x1_ASAP7_75t_L g627 ( 
.A1(n_591),
.A2(n_408),
.A3(n_593),
.B1(n_608),
.B2(n_592),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_589),
.B(n_500),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_570),
.B(n_504),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_578),
.A2(n_575),
.B(n_581),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_534),
.B(n_504),
.Y(n_631)
);

OR2x6_ASAP7_75t_SL g632 ( 
.A(n_564),
.B(n_606),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_615),
.Y(n_633)
);

BUFx8_ASAP7_75t_L g634 ( 
.A(n_609),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_553),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_543),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_433),
.B(n_455),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_573),
.A2(n_520),
.B1(n_455),
.B2(n_467),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_529),
.B(n_497),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_569),
.B(n_499),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_571),
.B(n_515),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_531),
.B(n_522),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_553),
.B(n_492),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_576),
.B(n_530),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_537),
.A2(n_466),
.B(n_507),
.C(n_492),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_561),
.B(n_52),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_533),
.B(n_53),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_610),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_555),
.A2(n_507),
.B1(n_527),
.B2(n_525),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_560),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_585),
.Y(n_653)
);

OR2x6_ASAP7_75t_SL g654 ( 
.A(n_542),
.B(n_54),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_573),
.A2(n_506),
.B1(n_505),
.B2(n_501),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_579),
.B(n_567),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_SL g658 ( 
.A1(n_563),
.A2(n_487),
.B(n_485),
.Y(n_658)
);

AOI33xp33_ASAP7_75t_L g659 ( 
.A1(n_614),
.A2(n_483),
.A3(n_471),
.B1(n_464),
.B2(n_461),
.B3(n_460),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_544),
.B(n_58),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_585),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_605),
.A2(n_414),
.B1(n_459),
.B2(n_427),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_594),
.B(n_614),
.C(n_541),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_535),
.A2(n_446),
.B1(n_437),
.B2(n_472),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_538),
.A2(n_437),
.B(n_447),
.C(n_445),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_539),
.B(n_61),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_568),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_540),
.Y(n_670)
);

AO21x1_ASAP7_75t_L g671 ( 
.A1(n_612),
.A2(n_74),
.B(n_75),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_563),
.B(n_76),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_554),
.B(n_77),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_574),
.A2(n_532),
.B1(n_617),
.B2(n_616),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_590),
.Y(n_675)
);

OR2x2_ASAP7_75t_SL g676 ( 
.A(n_602),
.B(n_101),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_618),
.A2(n_443),
.B1(n_108),
.B2(n_110),
.Y(n_677)
);

XOR2xp5_ASAP7_75t_L g678 ( 
.A(n_588),
.B(n_112),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_551),
.A2(n_443),
.B1(n_117),
.B2(n_119),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_550),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_549),
.A2(n_588),
.B1(n_611),
.B2(n_556),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_566),
.B(n_572),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_620),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_546),
.A2(n_149),
.B(n_150),
.Y(n_685)
);

CKINVDCx6p67_ASAP7_75t_R g686 ( 
.A(n_557),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_619),
.Y(n_687)
);

AO32x2_ASAP7_75t_L g688 ( 
.A1(n_582),
.A2(n_155),
.A3(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_600),
.B(n_174),
.Y(n_689)
);

NOR3xp33_ASAP7_75t_L g690 ( 
.A(n_604),
.B(n_548),
.C(n_565),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_598),
.A2(n_587),
.B(n_599),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_558),
.A2(n_562),
.B1(n_621),
.B2(n_607),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_595),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_603),
.A2(n_597),
.B1(n_590),
.B2(n_596),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_590),
.B(n_570),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_622),
.B(n_590),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_671),
.A2(n_681),
.A3(n_666),
.B(n_662),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_634),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_634),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_626),
.B(n_625),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_636),
.B(n_635),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_648),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_624),
.A2(n_674),
.B1(n_628),
.B2(n_650),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_SL g705 ( 
.A1(n_678),
.A2(n_654),
.B1(n_660),
.B2(n_641),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_632),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_670),
.B(n_642),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_687),
.B(n_674),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_681),
.A2(n_662),
.B1(n_643),
.B2(n_629),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_643),
.A2(n_640),
.B1(n_624),
.B2(n_656),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_661),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_669),
.B(n_652),
.Y(n_713)
);

AO31x2_ASAP7_75t_L g714 ( 
.A1(n_677),
.A2(n_679),
.A3(n_693),
.B(n_665),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_638),
.A2(n_691),
.B(n_658),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_656),
.B(n_692),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_696),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_643),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_686),
.B(n_664),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_668),
.Y(n_720)
);

NOR2x1_ASAP7_75t_SL g721 ( 
.A(n_675),
.B(n_694),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_677),
.A2(n_679),
.A3(n_693),
.B(n_665),
.Y(n_722)
);

BUFx8_ASAP7_75t_L g723 ( 
.A(n_688),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_694),
.A2(n_673),
.B1(n_639),
.B2(n_667),
.Y(n_724)
);

AO31x2_ASAP7_75t_L g725 ( 
.A1(n_684),
.A2(n_655),
.A3(n_647),
.B(n_685),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_659),
.B(n_690),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_684),
.A2(n_672),
.B(n_689),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_644),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_633),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_637),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_SL g731 ( 
.A1(n_651),
.A2(n_695),
.B(n_653),
.C(n_644),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_633),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_627),
.A2(n_680),
.B(n_683),
.Y(n_733)
);

AO31x2_ASAP7_75t_L g734 ( 
.A1(n_688),
.A2(n_671),
.A3(n_630),
.B(n_681),
.Y(n_734)
);

OAI21xp33_ASAP7_75t_SL g735 ( 
.A1(n_682),
.A2(n_688),
.B(n_676),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_682),
.A2(n_622),
.B1(n_646),
.B2(n_625),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_646),
.A2(n_674),
.B(n_681),
.C(n_592),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_634),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_622),
.A2(n_434),
.B1(n_545),
.B2(n_416),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_646),
.A2(n_575),
.B(n_649),
.C(n_631),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_626),
.B(n_545),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_622),
.B(n_626),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_632),
.Y(n_743)
);

AOI211x1_ASAP7_75t_L g744 ( 
.A1(n_662),
.A2(n_646),
.B(n_681),
.C(n_674),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_646),
.A2(n_575),
.B(n_649),
.C(n_631),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_622),
.B(n_626),
.Y(n_746)
);

INVxp67_ASAP7_75t_SL g747 ( 
.A(n_622),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_622),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_634),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_622),
.Y(n_751)
);

AO31x2_ASAP7_75t_L g752 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_622),
.A2(n_646),
.B1(n_625),
.B2(n_626),
.Y(n_753)
);

AO31x2_ASAP7_75t_L g754 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_622),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_622),
.B(n_570),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_626),
.B(n_545),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_634),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_673),
.B(n_645),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_622),
.B(n_528),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_622),
.Y(n_761)
);

AO31x2_ASAP7_75t_L g762 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_622),
.B(n_528),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_622),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_528),
.Y(n_765)
);

AOI221x1_ASAP7_75t_L g766 ( 
.A1(n_681),
.A2(n_630),
.B1(n_662),
.B2(n_663),
.C(n_684),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

AO31x2_ASAP7_75t_L g768 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_622),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_622),
.B(n_528),
.Y(n_770)
);

CKINVDCx11_ASAP7_75t_R g771 ( 
.A(n_632),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_622),
.B(n_570),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_622),
.B(n_626),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_646),
.A2(n_575),
.B(n_649),
.C(n_631),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_622),
.A2(n_646),
.B1(n_625),
.B2(n_626),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_622),
.B(n_528),
.Y(n_779)
);

AO31x2_ASAP7_75t_L g780 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_780)
);

NAND3x1_ASAP7_75t_L g781 ( 
.A(n_648),
.B(n_555),
.C(n_365),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_622),
.B(n_570),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_622),
.B(n_625),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_622),
.B(n_528),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_785)
);

BUFx2_ASAP7_75t_R g786 ( 
.A(n_632),
.Y(n_786)
);

AOI211x1_ASAP7_75t_L g787 ( 
.A1(n_662),
.A2(n_646),
.B(n_681),
.C(n_674),
.Y(n_787)
);

AO31x2_ASAP7_75t_L g788 ( 
.A1(n_671),
.A2(n_630),
.A3(n_681),
.B(n_575),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_675),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_L g790 ( 
.A1(n_622),
.A2(n_570),
.B(n_646),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_646),
.A2(n_674),
.B(n_681),
.C(n_592),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_622),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_622),
.B(n_528),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_661),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_622),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_622),
.B(n_552),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_626),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_622),
.B(n_528),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_760),
.B(n_763),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_704),
.A2(n_777),
.B1(n_753),
.B2(n_747),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_737),
.A2(n_791),
.B(n_745),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_765),
.B(n_770),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_SL g804 ( 
.A1(n_724),
.A2(n_736),
.B(n_709),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_779),
.B(n_784),
.Y(n_805)
);

OA21x2_ASAP7_75t_L g806 ( 
.A1(n_715),
.A2(n_733),
.B(n_766),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_761),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_771),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_767),
.Y(n_809)
);

AO21x2_ASAP7_75t_L g810 ( 
.A1(n_731),
.A2(n_710),
.B(n_726),
.Y(n_810)
);

INVx3_ASAP7_75t_SL g811 ( 
.A(n_738),
.Y(n_811)
);

NAND2x1_ASAP7_75t_L g812 ( 
.A(n_759),
.B(n_728),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_727),
.A2(n_740),
.B(n_776),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_793),
.B(n_798),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_775),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_742),
.B(n_746),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_778),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_773),
.B(n_797),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_741),
.B(n_757),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_792),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_750),
.B(n_751),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_711),
.A2(n_744),
.B1(n_787),
.B2(n_755),
.Y(n_822)
);

OA21x2_ASAP7_75t_L g823 ( 
.A1(n_718),
.A2(n_734),
.B(n_697),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_749),
.B(n_774),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_699),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_781),
.A2(n_764),
.B(n_795),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_739),
.B(n_769),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_786),
.B(n_758),
.Y(n_828)
);

OAI21x1_ASAP7_75t_SL g829 ( 
.A1(n_721),
.A2(n_728),
.B(n_701),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_756),
.B(n_772),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_783),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_720),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_789),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_782),
.B(n_790),
.Y(n_834)
);

AO31x2_ASAP7_75t_L g835 ( 
.A1(n_734),
.A2(n_780),
.A3(n_752),
.B(n_788),
.Y(n_835)
);

AO31x2_ASAP7_75t_L g836 ( 
.A1(n_752),
.A2(n_768),
.A3(n_754),
.B(n_788),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_713),
.A2(n_723),
.B1(n_707),
.B2(n_705),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_789),
.B(n_700),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_752),
.A2(n_754),
.B(n_762),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_730),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_707),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_716),
.A2(n_759),
.B(n_719),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_729),
.A2(n_732),
.B(n_785),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_759),
.B(n_702),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_789),
.B(n_712),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_796),
.B(n_706),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_796),
.A2(n_703),
.B1(n_708),
.B2(n_723),
.Y(n_847)
);

BUFx8_ASAP7_75t_L g848 ( 
.A(n_743),
.Y(n_848)
);

AO31x2_ASAP7_75t_L g849 ( 
.A1(n_698),
.A2(n_725),
.A3(n_714),
.B(n_722),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_729),
.A2(n_732),
.B(n_714),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_722),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_794),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_698),
.A2(n_725),
.B(n_722),
.Y(n_853)
);

AOI21xp33_ASAP7_75t_SL g854 ( 
.A1(n_717),
.A2(n_509),
.B(n_743),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_748),
.B(n_761),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_747),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_747),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_748),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_738),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_771),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_738),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_748),
.Y(n_862)
);

OAI211xp5_ASAP7_75t_L g863 ( 
.A1(n_735),
.A2(n_416),
.B(n_614),
.C(n_747),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_760),
.B(n_763),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_748),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_748),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

BUFx12f_ASAP7_75t_L g868 ( 
.A(n_771),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_748),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_822),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_856),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_804),
.B(n_813),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_856),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_829),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_857),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_816),
.B(n_799),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_800),
.B(n_827),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_832),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_801),
.B(n_800),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_849),
.B(n_853),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_827),
.B(n_799),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_812),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_840),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_849),
.B(n_803),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_849),
.B(n_803),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_816),
.B(n_805),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_805),
.B(n_814),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_850),
.B(n_843),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_849),
.B(n_814),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_851),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_865),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_864),
.B(n_839),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_864),
.B(n_810),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_874),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_874),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_871),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_879),
.B(n_836),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_892),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_892),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_884),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_871),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_873),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_884),
.B(n_823),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_874),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_882),
.B(n_837),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_879),
.A2(n_837),
.B1(n_834),
.B2(n_826),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_875),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_874),
.B(n_847),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_884),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_879),
.B(n_885),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_875),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_835),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_870),
.B(n_844),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_891),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_889),
.B(n_819),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_806),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_872),
.B(n_835),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_890),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_887),
.B(n_876),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_870),
.B(n_806),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_900),
.B(n_880),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_900),
.B(n_880),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_914),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_918),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_909),
.B(n_880),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_915),
.B(n_893),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_915),
.B(n_877),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_910),
.B(n_897),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_911),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_907),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_917),
.B(n_888),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_895),
.B(n_846),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_898),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_910),
.B(n_877),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_899),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_929),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_924),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_926),
.B(n_899),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_931),
.B(n_888),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_921),
.B(n_916),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_921),
.B(n_916),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_930),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_922),
.B(n_920),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_922),
.B(n_920),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_925),
.B(n_903),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_926),
.B(n_912),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_935),
.B(n_933),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_925),
.B(n_903),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_936),
.B(n_923),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_947),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_936),
.B(n_928),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_942),
.B(n_932),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_939),
.B(n_931),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_937),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_L g955 ( 
.A1(n_942),
.A2(n_932),
.B(n_908),
.Y(n_955)
);

AND2x2_ASAP7_75t_SL g956 ( 
.A(n_939),
.B(n_895),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_938),
.Y(n_957)
);

OAI32xp33_ASAP7_75t_L g958 ( 
.A1(n_938),
.A2(n_895),
.A3(n_808),
.B1(n_891),
.B2(n_894),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_946),
.B(n_934),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_946),
.A2(n_905),
.B1(n_906),
.B2(n_919),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_947),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_940),
.B(n_928),
.Y(n_962)
);

NAND4xp25_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_828),
.C(n_905),
.D(n_863),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_949),
.B(n_868),
.Y(n_964)
);

OAI211xp5_ASAP7_75t_SL g965 ( 
.A1(n_952),
.A2(n_863),
.B(n_859),
.C(n_861),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_951),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_957),
.B(n_945),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_954),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_959),
.B(n_945),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_956),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_956),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_SL g973 ( 
.A1(n_952),
.A2(n_808),
.B(n_904),
.C(n_901),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_SL g974 ( 
.A1(n_955),
.A2(n_945),
.B(n_948),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_959),
.B(n_948),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_962),
.B(n_940),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_958),
.A2(n_907),
.B(n_939),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_SL g978 ( 
.A1(n_960),
.A2(n_913),
.B1(n_895),
.B2(n_931),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_974),
.A2(n_963),
.B1(n_953),
.B2(n_913),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_974),
.A2(n_953),
.B1(n_913),
.B2(n_950),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_972),
.A2(n_913),
.B1(n_961),
.B2(n_931),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_978),
.A2(n_913),
.B1(n_934),
.B2(n_927),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_972),
.A2(n_913),
.B1(n_940),
.B2(n_944),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_L g984 ( 
.A1(n_973),
.A2(n_860),
.B(n_854),
.C(n_826),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_971),
.A2(n_913),
.B1(n_944),
.B2(n_943),
.Y(n_985)
);

OAI22xp33_ASAP7_75t_L g986 ( 
.A1(n_977),
.A2(n_904),
.B1(n_894),
.B2(n_872),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_941),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_964),
.A2(n_970),
.B(n_967),
.C(n_975),
.Y(n_988)
);

OAI211xp5_ASAP7_75t_SL g989 ( 
.A1(n_979),
.A2(n_966),
.B(n_842),
.C(n_881),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_988),
.A2(n_965),
.B1(n_967),
.B2(n_976),
.C(n_968),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_987),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_980),
.B(n_941),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_982),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_983),
.A2(n_904),
.B1(n_894),
.B2(n_872),
.Y(n_994)
);

AOI21xp33_ASAP7_75t_SL g995 ( 
.A1(n_986),
.A2(n_811),
.B(n_824),
.Y(n_995)
);

AOI221x1_ASAP7_75t_L g996 ( 
.A1(n_984),
.A2(n_968),
.B1(n_969),
.B2(n_883),
.C(n_878),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_981),
.A2(n_896),
.B(n_902),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_991),
.B(n_825),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_995),
.B(n_969),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_825),
.C(n_820),
.Y(n_1000)
);

NAND4xp25_ASAP7_75t_SL g1001 ( 
.A(n_996),
.B(n_870),
.C(n_848),
.D(n_919),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_993),
.Y(n_1002)
);

OA211x2_ASAP7_75t_L g1003 ( 
.A1(n_990),
.A2(n_848),
.B(n_842),
.C(n_811),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_997),
.B(n_838),
.C(n_845),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_833),
.Y(n_1005)
);

NAND2x1_ASAP7_75t_L g1006 ( 
.A(n_1004),
.B(n_992),
.Y(n_1006)
);

NOR4xp75_ASAP7_75t_L g1007 ( 
.A(n_1002),
.B(n_881),
.C(n_994),
.D(n_824),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_998),
.Y(n_1008)
);

NOR2x1_ASAP7_75t_L g1009 ( 
.A(n_1001),
.B(n_824),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1000),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_SL g1011 ( 
.A1(n_1003),
.A2(n_943),
.B(n_882),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_SL g1012 ( 
.A(n_1001),
.B(n_841),
.C(n_802),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_1009),
.B(n_833),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1008),
.A2(n_1006),
.B1(n_1010),
.B2(n_1005),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1012),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_1011),
.B(n_830),
.C(n_867),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_1007),
.B(n_867),
.C(n_809),
.Y(n_1017)
);

NAND4xp25_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_855),
.C(n_876),
.D(n_886),
.Y(n_1018)
);

XNOR2x1_ASAP7_75t_L g1019 ( 
.A(n_1015),
.B(n_838),
.Y(n_1019)
);

OR3x2_ASAP7_75t_L g1020 ( 
.A(n_1018),
.B(n_815),
.C(n_807),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_1019),
.A2(n_1013),
.B1(n_1020),
.B2(n_1014),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1021),
.B(n_1016),
.Y(n_1022)
);

AOI222xp33_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_1017),
.B1(n_866),
.B2(n_869),
.C1(n_862),
.C2(n_858),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1023),
.A2(n_846),
.B1(n_845),
.B2(n_817),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_1024),
.B(n_846),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_1025),
.A2(n_831),
.B1(n_821),
.B2(n_852),
.Y(n_1026)
);


endmodule