module fake_aes_8527_n_729 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_729);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_729;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_135;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_716;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g80 ( .A(n_42), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_25), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_74), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_24), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_61), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_40), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_51), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_68), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_78), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_41), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_5), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_23), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_4), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_14), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_75), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_12), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_44), .Y(n_102) );
XNOR2xp5_ASAP7_75t_L g103 ( .A(n_10), .B(n_53), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_37), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_21), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_5), .B(n_15), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_56), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_3), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_9), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_22), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_26), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_71), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_6), .Y(n_120) );
INVx2_ASAP7_75t_SL g121 ( .A(n_69), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_27), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_18), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_6), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_17), .Y(n_127) );
INVxp33_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_3), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_115), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_121), .B(n_0), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_116), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_110), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_110), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_87), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_117), .Y(n_145) );
AND3x1_ASAP7_75t_L g146 ( .A(n_106), .B(n_1), .C(n_2), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_95), .B(n_1), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_85), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_85), .A2(n_4), .B(n_7), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
NAND2xp33_ASAP7_75t_L g152 ( .A(n_116), .B(n_35), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_117), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_117), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_117), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_116), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_86), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_95), .B(n_7), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_88), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_89), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_106), .B(n_8), .Y(n_168) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_89), .A2(n_38), .B(n_70), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_87), .B(n_9), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g171 ( .A(n_119), .B(n_76), .Y(n_171) );
CKINVDCx8_ASAP7_75t_R g172 ( .A(n_119), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_116), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_132), .B(n_97), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_170), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_132), .B(n_94), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_170), .B(n_98), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_140), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_168), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_172), .A2(n_129), .B1(n_98), .B2(n_101), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_134), .B(n_128), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_132), .B(n_101), .Y(n_187) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_170), .B(n_129), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_168), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_168), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_134), .B(n_120), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_136), .B(n_114), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_147), .B(n_80), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_147), .B(n_122), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx4_ASAP7_75t_L g204 ( .A(n_150), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_144), .B(n_127), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
AND3x4_ASAP7_75t_L g207 ( .A(n_172), .B(n_103), .C(n_111), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_130), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_130), .B(n_92), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_133), .Y(n_213) );
INVxp67_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_138), .B(n_113), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_138), .B(n_113), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_142), .B(n_105), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g220 ( .A(n_171), .B(n_105), .C(n_125), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_149), .B(n_107), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_149), .B(n_99), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_154), .B(n_166), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_140), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_154), .B(n_91), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_155), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_166), .B(n_125), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_140), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_155), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_167), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_172), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_140), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_167), .B(n_107), .Y(n_236) );
INVxp67_ASAP7_75t_L g237 ( .A(n_148), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_160), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_146), .B(n_114), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_159), .Y(n_240) );
AND2x6_ASAP7_75t_L g241 ( .A(n_159), .B(n_99), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_239), .A2(n_171), .B1(n_150), .B2(n_164), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_225), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_204), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_237), .B(n_146), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_225), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_225), .B(n_91), .Y(n_249) );
INVx4_ASAP7_75t_L g250 ( .A(n_193), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_233), .B(n_148), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_214), .B(n_164), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_193), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_178), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_185), .B(n_83), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_234), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_176), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_177), .B(n_84), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_185), .B(n_102), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_187), .B(n_123), .Y(n_262) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_198), .B(n_100), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_187), .B(n_159), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_224), .Y(n_266) );
AO22x1_ASAP7_75t_L g267 ( .A1(n_207), .A2(n_126), .B1(n_103), .B2(n_109), .Y(n_267) );
INVx5_ASAP7_75t_L g268 ( .A(n_241), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_174), .B(n_118), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_224), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_230), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_230), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_188), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_188), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_230), .Y(n_277) );
AND2x6_ASAP7_75t_L g278 ( .A(n_195), .B(n_100), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_219), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_174), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_187), .B(n_165), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_239), .A2(n_150), .B1(n_118), .B2(n_165), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_200), .B(n_112), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_234), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_241), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_197), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_239), .B(n_169), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_210), .B(n_162), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_196), .B(n_124), .Y(n_292) );
NAND2x1p5_ASAP7_75t_L g293 ( .A(n_219), .B(n_150), .Y(n_293) );
OR2x6_ASAP7_75t_L g294 ( .A(n_197), .B(n_169), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_222), .B(n_165), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_205), .Y(n_296) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_205), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_222), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_184), .A2(n_108), .B1(n_111), .B2(n_93), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_236), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_229), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_241), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_208), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_180), .A2(n_162), .B(n_163), .C(n_165), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_236), .B(n_96), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_229), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_199), .B(n_162), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_208), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_201), .A2(n_169), .B(n_152), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_241), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_244), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_258), .B(n_197), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_302), .B(n_209), .Y(n_316) );
NOR2xp33_ASAP7_75t_SL g317 ( .A(n_246), .B(n_207), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_309), .B(n_220), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_309), .A2(n_190), .B(n_189), .C(n_183), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
BUFx5_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_263), .A2(n_203), .B(n_218), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_250), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_283), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_250), .Y(n_327) );
INVx5_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_244), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_266), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_245), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_296), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_247), .A2(n_202), .B1(n_199), .B2(n_213), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_266), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_251), .B(n_221), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_255), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_251), .B(n_202), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_307), .A2(n_215), .B(n_223), .C(n_227), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_252), .B(n_215), .Y(n_342) );
OR2x2_ASAP7_75t_SL g343 ( .A(n_275), .B(n_112), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_276), .Y(n_344) );
BUFx8_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_242), .B(n_223), .C(n_218), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_255), .B(n_208), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_260), .B(n_240), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_300), .Y(n_349) );
NOR2x1_ASAP7_75t_R g350 ( .A(n_257), .B(n_104), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_297), .B(n_162), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_266), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_247), .A2(n_241), .B1(n_124), .B2(n_163), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_262), .B(n_163), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_247), .A2(n_163), .B1(n_160), .B2(n_152), .Y(n_357) );
INVx6_ASAP7_75t_SL g358 ( .A(n_290), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_297), .B(n_10), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_267), .B(n_160), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_243), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_292), .B(n_11), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_245), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_270), .A2(n_292), .B(n_265), .C(n_284), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_289), .B(n_11), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_263), .A2(n_238), .B(n_232), .Y(n_366) );
NAND3xp33_ASAP7_75t_L g367 ( .A(n_260), .B(n_238), .C(n_232), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_256), .B(n_13), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_261), .B(n_13), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_333), .B(n_262), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_328), .B(n_289), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_326), .A2(n_257), .B1(n_287), .B2(n_278), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_248), .B1(n_278), .B2(n_290), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_278), .B1(n_290), .B2(n_249), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_324), .Y(n_375) );
AO21x1_ASAP7_75t_L g376 ( .A1(n_364), .A2(n_293), .B(n_312), .Y(n_376) );
CKINVDCx11_ASAP7_75t_R g377 ( .A(n_337), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_344), .B(n_299), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_365), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_365), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_316), .A2(n_295), .B1(n_253), .B2(n_285), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_342), .B(n_278), .Y(n_382) );
INVx6_ASAP7_75t_L g383 ( .A(n_328), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_253), .B1(n_249), .B2(n_250), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_360), .A2(n_286), .B1(n_269), .B2(n_259), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_287), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_320), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_317), .A2(n_259), .B1(n_269), .B2(n_286), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_310), .B1(n_291), .B2(n_269), .C(n_259), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_360), .A2(n_264), .B1(n_279), .B2(n_280), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_336), .B(n_305), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_348), .A2(n_293), .B1(n_264), .B2(n_294), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
OR2x6_ASAP7_75t_L g395 ( .A(n_360), .B(n_288), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_356), .A2(n_160), .B(n_305), .C(n_145), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
AOI221xp5_ASAP7_75t_SL g398 ( .A1(n_341), .A2(n_280), .B1(n_279), .B2(n_274), .C(n_254), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_348), .A2(n_294), .B1(n_277), .B2(n_271), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_330), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_334), .A2(n_294), .B1(n_277), .B2(n_271), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_358), .A2(n_294), .B1(n_277), .B2(n_271), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_321), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_388), .B(n_403), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_400), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_395), .Y(n_406) );
AOI21xp33_ASAP7_75t_SL g407 ( .A1(n_372), .A2(n_369), .B(n_368), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_393), .A2(n_373), .B1(n_401), .B2(n_374), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_392), .Y(n_409) );
AO31x2_ASAP7_75t_L g410 ( .A1(n_376), .A2(n_131), .A3(n_145), .B(n_369), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_400), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_315), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_375), .A2(n_345), .B1(n_368), .B2(n_359), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_379), .A2(n_345), .B1(n_380), .B2(n_399), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_370), .B(n_343), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_351), .B1(n_362), .B2(n_367), .Y(n_417) );
AOI332xp33_ASAP7_75t_L g418 ( .A1(n_374), .A2(n_354), .A3(n_357), .B1(n_352), .B2(n_349), .B3(n_339), .C1(n_361), .C2(n_131), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_397), .A2(n_356), .B1(n_319), .B2(n_346), .C(n_357), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_373), .B(n_347), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_384), .A2(n_318), .B1(n_325), .B2(n_327), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_381), .A2(n_323), .B(n_319), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_323), .B1(n_325), .B2(n_327), .C(n_305), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_402), .A2(n_322), .B1(n_353), .B2(n_335), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_395), .A2(n_322), .B1(n_353), .B2(n_335), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_396), .A2(n_322), .B1(n_271), .B2(n_277), .Y(n_426) );
OAI22xp33_ASAP7_75t_SL g427 ( .A1(n_395), .A2(n_350), .B1(n_328), .B2(n_314), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_398), .A2(n_366), .B1(n_254), .B2(n_272), .C(n_273), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_385), .B(n_272), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_395), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_377), .A2(n_322), .B1(n_274), .B2(n_273), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_407), .A2(n_385), .B1(n_391), .B2(n_389), .C(n_366), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_413), .B(n_377), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_416), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_416), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_413), .A2(n_391), .B1(n_383), .B2(n_322), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_420), .B(n_371), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_420), .B(n_371), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_404), .B(n_409), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_408), .A2(n_383), .B1(n_322), .B2(n_386), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_408), .A2(n_383), .B1(n_330), .B2(n_353), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_407), .B(n_329), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_422), .A2(n_363), .B(n_331), .Y(n_444) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_414), .A2(n_145), .B(n_131), .C(n_160), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_415), .A2(n_394), .B1(n_353), .B2(n_335), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_409), .A2(n_335), .B1(n_332), .B2(n_400), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_412), .B(n_288), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_406), .B(n_394), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_419), .A2(n_332), .B1(n_400), .B2(n_131), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_332), .B1(n_328), .B2(n_313), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_429), .B(n_412), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_427), .A2(n_145), .A3(n_139), .B1(n_143), .B2(n_135), .B3(n_153), .Y(n_454) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_430), .A2(n_135), .B(n_139), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_425), .A2(n_332), .B1(n_15), .B2(n_16), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_427), .A2(n_423), .B1(n_417), .B2(n_431), .C(n_432), .Y(n_457) );
CKINVDCx10_ASAP7_75t_R g458 ( .A(n_418), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_429), .B(n_14), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_405), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_421), .B(n_135), .C(n_139), .D(n_143), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_405), .B(n_313), .Y(n_462) );
OAI21xp33_ASAP7_75t_SL g463 ( .A1(n_426), .A2(n_311), .B(n_153), .Y(n_463) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_424), .B(n_173), .C(n_161), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_405), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_428), .B(n_143), .C(n_153), .D(n_157), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_410), .B(n_311), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_418), .A2(n_173), .B1(n_161), .B2(n_157), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_411), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_460), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_446), .B(n_410), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_435), .B(n_410), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_440), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_457), .B(n_157), .C(n_158), .D(n_19), .Y(n_474) );
NOR3xp33_ASAP7_75t_SL g475 ( .A(n_434), .B(n_16), .C(n_17), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_438), .B(n_410), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_453), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_436), .B(n_410), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_438), .B(n_410), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_439), .B(n_411), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_467), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_469), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_439), .B(n_411), .Y(n_483) );
INVxp67_ASAP7_75t_R g484 ( .A(n_456), .Y(n_484) );
OAI33xp33_ASAP7_75t_L g485 ( .A1(n_442), .A2(n_158), .A3(n_20), .B1(n_21), .B2(n_23), .B3(n_19), .Y(n_485) );
OAI211xp5_ASAP7_75t_SL g486 ( .A1(n_447), .A2(n_158), .B(n_228), .C(n_216), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_465), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_450), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_450), .B(n_20), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_468), .B(n_173), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_173), .Y(n_492) );
OAI31xp33_ASAP7_75t_L g493 ( .A1(n_468), .A2(n_192), .A3(n_186), .B(n_194), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g494 ( .A1(n_461), .A2(n_173), .A3(n_161), .B1(n_216), .B2(n_212), .B3(n_206), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_455), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_455), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_443), .A2(n_268), .B(n_304), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_458), .B(n_303), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_443), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_441), .B(n_173), .Y(n_501) );
OAI222xp33_ASAP7_75t_L g502 ( .A1(n_447), .A2(n_268), .B1(n_304), .B2(n_30), .C1(n_32), .C2(n_33), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_454), .A2(n_161), .B1(n_173), .B2(n_140), .C(n_141), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_462), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_445), .B(n_161), .C(n_173), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_448), .B(n_313), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_433), .A2(n_161), .B1(n_141), .B2(n_151), .C(n_156), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_437), .B(n_449), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_437), .B(n_161), .Y(n_509) );
NAND5xp2_ASAP7_75t_L g510 ( .A(n_451), .B(n_268), .C(n_304), .D(n_34), .E(n_36), .Y(n_510) );
OAI221xp5_ASAP7_75t_L g511 ( .A1(n_451), .A2(n_161), .B1(n_313), .B2(n_303), .C(n_288), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_466), .B(n_192), .C(n_228), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_463), .B(n_141), .C(n_156), .Y(n_513) );
AND2x4_ASAP7_75t_SL g514 ( .A(n_449), .B(n_303), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_141), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_456), .A2(n_186), .A3(n_179), .B(n_175), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_446), .B(n_141), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_448), .A2(n_303), .B(n_304), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_446), .B(n_156), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_460), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_446), .B(n_156), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_453), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_477), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_521), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_484), .A2(n_304), .B1(n_268), .B2(n_141), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_470), .Y(n_527) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_474), .B(n_156), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_473), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_523), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_471), .B(n_156), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_523), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_472), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_478), .Y(n_536) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_474), .B(n_156), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_521), .B(n_156), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_484), .A2(n_268), .B1(n_141), .B2(n_151), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_498), .A2(n_151), .B(n_141), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_490), .B(n_151), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_489), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_489), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_518), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_500), .B(n_151), .Y(n_545) );
NAND2xp33_ASAP7_75t_L g546 ( .A(n_475), .B(n_151), .Y(n_546) );
INVxp33_ASAP7_75t_L g547 ( .A(n_470), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_470), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_518), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_476), .B(n_151), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_481), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_476), .B(n_151), .Y(n_552) );
NOR3xp33_ASAP7_75t_SL g553 ( .A(n_510), .B(n_28), .C(n_29), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_479), .B(n_45), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_483), .B(n_46), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_483), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_481), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_479), .B(n_47), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_522), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_471), .B(n_48), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_500), .B(n_49), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_488), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_522), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_487), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_485), .B(n_175), .C(n_212), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_494), .B(n_206), .C(n_194), .Y(n_568) );
XNOR2xp5_ASAP7_75t_L g569 ( .A(n_480), .B(n_50), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_487), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_480), .B(n_52), .Y(n_571) );
HB1xp67_ASAP7_75t_SL g572 ( .A(n_488), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_482), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_508), .A2(n_235), .B1(n_231), .B2(n_226), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_514), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_500), .B(n_54), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_55), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_509), .A2(n_58), .B(n_59), .Y(n_578) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_486), .A2(n_516), .A3(n_501), .B1(n_492), .B2(n_514), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_482), .B(n_60), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_482), .B(n_62), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_514), .B(n_65), .Y(n_582) );
AOI31xp67_ASAP7_75t_L g583 ( .A1(n_504), .A2(n_179), .A3(n_66), .B(n_67), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_499), .B(n_235), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_525), .B(n_501), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_529), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_579), .B(n_517), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_540), .A2(n_517), .B(n_493), .C(n_513), .Y(n_588) );
INVxp33_ASAP7_75t_L g589 ( .A(n_572), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_524), .B(n_499), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_527), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_530), .B(n_499), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_532), .B(n_492), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_557), .B(n_496), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_533), .B(n_495), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_550), .B(n_496), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_534), .B(n_495), .Y(n_598) );
CKINVDCx16_ASAP7_75t_R g599 ( .A(n_569), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_570), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_535), .Y(n_601) );
NOR3xp33_ASAP7_75t_SL g602 ( .A(n_539), .B(n_502), .C(n_513), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_548), .B(n_495), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_548), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_542), .B(n_516), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_552), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_546), .A2(n_516), .B1(n_493), .B2(n_497), .C(n_507), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_543), .B(n_504), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_552), .B(n_504), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g612 ( .A1(n_537), .A2(n_505), .B(n_506), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_564), .B(n_495), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_551), .B(n_491), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_541), .B(n_505), .C(n_503), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_531), .B(n_515), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_551), .B(n_511), .Y(n_617) );
AND3x2_ASAP7_75t_L g618 ( .A(n_554), .B(n_512), .C(n_519), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_547), .B(n_181), .Y(n_619) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_563), .B(n_181), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_546), .B(n_181), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_544), .B(n_235), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_558), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_545), .B(n_553), .C(n_531), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_554), .B(n_181), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_558), .B(n_191), .Y(n_626) );
AOI33xp33_ASAP7_75t_L g627 ( .A1(n_577), .A2(n_191), .A3(n_211), .B1(n_217), .B2(n_226), .B3(n_231), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_560), .B(n_191), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_573), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_560), .B(n_191), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_575), .Y(n_631) );
OR2x6_ASAP7_75t_L g632 ( .A(n_562), .B(n_211), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_555), .B(n_235), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_559), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_561), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_599), .B(n_528), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_601), .B(n_531), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_587), .A2(n_526), .B(n_577), .C(n_571), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_589), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_586), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_632), .B(n_538), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_597), .B(n_573), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_629), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_603), .B(n_565), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_589), .B(n_562), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_591), .B(n_562), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_631), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_597), .B(n_545), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_610), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_594), .B(n_556), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_596), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_600), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_633), .B(n_576), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_588), .A2(n_582), .B(n_563), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_587), .A2(n_563), .B1(n_567), .B2(n_576), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_585), .Y(n_659) );
XNOR2x1_ASAP7_75t_L g660 ( .A(n_632), .B(n_581), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_629), .B(n_581), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_590), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_635), .Y(n_663) );
AOI321xp33_ASAP7_75t_L g664 ( .A1(n_605), .A2(n_580), .A3(n_574), .B1(n_568), .B2(n_578), .C(n_584), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_611), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_636), .B(n_580), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_608), .B(n_584), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_592), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_607), .B(n_583), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_595), .B(n_211), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_632), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_623), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_616), .Y(n_673) );
AO22x2_ASAP7_75t_L g674 ( .A1(n_595), .A2(n_211), .B1(n_217), .B2(n_226), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_598), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_588), .A2(n_231), .B(n_217), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_593), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g678 ( .A1(n_627), .A2(n_226), .B1(n_231), .B2(n_609), .C(n_624), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_613), .B(n_616), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_614), .Y(n_680) );
AOI211x1_ASAP7_75t_L g681 ( .A1(n_612), .A2(n_615), .B(n_614), .C(n_630), .Y(n_681) );
XOR2x2_ASAP7_75t_L g682 ( .A(n_618), .B(n_620), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_617), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_602), .B(n_627), .C(n_604), .Y(n_684) );
NAND2xp33_ASAP7_75t_SL g685 ( .A(n_602), .B(n_616), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_625), .Y(n_686) );
AOI211xp5_ASAP7_75t_SL g687 ( .A1(n_621), .A2(n_628), .B(n_595), .C(n_619), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_626), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_622), .B(n_634), .C(n_621), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_618), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_601), .B(n_529), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_587), .A2(n_484), .B1(n_528), .B2(n_546), .Y(n_692) );
AOI221x1_ASAP7_75t_L g693 ( .A1(n_685), .A2(n_690), .B1(n_676), .B2(n_684), .C(n_683), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_681), .B(n_662), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_685), .A2(n_648), .B(n_678), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_641), .A2(n_655), .B1(n_654), .B2(n_677), .C(n_676), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_691), .A2(n_642), .B1(n_652), .B2(n_668), .C(n_650), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_646), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_637), .A2(n_692), .A3(n_648), .B(n_687), .Y(n_699) );
AO22x2_ASAP7_75t_L g700 ( .A1(n_637), .A2(n_646), .B1(n_660), .B2(n_663), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_645), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_675), .A2(n_665), .B1(n_678), .B2(n_659), .C(n_680), .Y(n_702) );
AOI221xp5_ASAP7_75t_SL g703 ( .A1(n_657), .A2(n_658), .B1(n_649), .B2(n_644), .C(n_639), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_682), .B(n_671), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_644), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_640), .A2(n_660), .B(n_643), .Y(n_706) );
OAI211xp5_ASAP7_75t_SL g707 ( .A1(n_706), .A2(n_664), .B(n_669), .C(n_679), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_701), .Y(n_708) );
OAI21xp33_ASAP7_75t_SL g709 ( .A1(n_699), .A2(n_673), .B(n_638), .Y(n_709) );
OAI21x1_ASAP7_75t_SL g710 ( .A1(n_695), .A2(n_667), .B(n_647), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_703), .B(n_651), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_700), .A2(n_666), .B1(n_651), .B2(n_686), .C(n_667), .Y(n_712) );
AOI21xp33_ASAP7_75t_SL g713 ( .A1(n_700), .A2(n_674), .B(n_689), .Y(n_713) );
OA22x2_ASAP7_75t_L g714 ( .A1(n_693), .A2(n_656), .B1(n_688), .B2(n_672), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_709), .B(n_702), .C(n_694), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_711), .B(n_704), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_708), .B(n_697), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_714), .Y(n_718) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_713), .B(n_696), .C(n_698), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_719), .B(n_712), .C(n_707), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_717), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_720), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_722), .Y(n_724) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_721), .B(n_716), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_724), .A2(n_715), .B1(n_710), .B2(n_705), .C(n_689), .Y(n_726) );
NOR2x1p5_ASAP7_75t_L g727 ( .A(n_725), .B(n_723), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_726), .B1(n_653), .B2(n_661), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_670), .B(n_674), .Y(n_729) );
endmodule