module real_aes_4672_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
HB1xp67_ASAP7_75t_L g175 ( .A(n_0), .Y(n_175) );
INVx1_ASAP7_75t_L g365 ( .A(n_1), .Y(n_365) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_1), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_2), .A2(n_13), .B1(n_207), .B2(n_267), .Y(n_275) );
INVx2_ASAP7_75t_L g246 ( .A(n_3), .Y(n_246) );
INVx1_ASAP7_75t_SL g322 ( .A(n_4), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_5), .A2(n_48), .B1(n_113), .B2(n_119), .Y(n_112) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_6), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_7), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_8), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_9), .B(n_55), .Y(n_147) );
INVxp67_ASAP7_75t_L g160 ( .A(n_9), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_10), .A2(n_41), .B1(n_336), .B2(n_337), .Y(n_335) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_11), .A2(n_53), .B(n_228), .Y(n_227) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_11), .A2(n_53), .B(n_228), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_12), .B(n_91), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_14), .B(n_242), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_15), .A2(n_61), .B1(n_231), .B2(n_234), .Y(n_230) );
INVx2_ASAP7_75t_L g271 ( .A(n_16), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_17), .A2(n_21), .B1(n_277), .B2(n_279), .Y(n_276) );
BUFx3_ASAP7_75t_L g184 ( .A(n_18), .Y(n_184) );
O2A1O1Ixp5_ASAP7_75t_L g264 ( .A1(n_19), .A2(n_203), .B(n_265), .C(n_266), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_20), .A2(n_49), .B1(n_239), .B2(n_241), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_22), .Y(n_308) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_24), .A2(n_62), .B1(n_344), .B2(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g258 ( .A(n_25), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_26), .A2(n_66), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g92 ( .A(n_27), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_27), .B(n_54), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_28), .B(n_254), .Y(n_360) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_28), .Y(n_635) );
INVx2_ASAP7_75t_L g268 ( .A(n_29), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g86 ( .A1(n_30), .A2(n_75), .B1(n_87), .B2(n_109), .Y(n_86) );
AOI221xp5_ASAP7_75t_SL g136 ( .A1(n_31), .A2(n_68), .B1(n_137), .B2(n_140), .C(n_141), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_32), .Y(n_310) );
INVx2_ASAP7_75t_L g388 ( .A(n_33), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_34), .Y(n_151) );
AOI221xp5_ASAP7_75t_L g152 ( .A1(n_35), .A2(n_50), .B1(n_153), .B2(n_154), .C(n_161), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_36), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g326 ( .A(n_37), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_38), .A2(n_47), .B1(n_127), .B2(n_135), .Y(n_126) );
INVx1_ASAP7_75t_L g304 ( .A(n_39), .Y(n_304) );
INVx1_ASAP7_75t_L g228 ( .A(n_40), .Y(n_228) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_42), .Y(n_195) );
AND2x4_ASAP7_75t_L g199 ( .A(n_42), .B(n_193), .Y(n_199) );
AND2x4_ASAP7_75t_L g262 ( .A(n_42), .B(n_193), .Y(n_262) );
INVx1_ASAP7_75t_L g331 ( .A(n_43), .Y(n_331) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_44), .Y(n_204) );
INVx2_ASAP7_75t_L g81 ( .A(n_45), .Y(n_81) );
AO22x1_ASAP7_75t_L g161 ( .A1(n_46), .A2(n_64), .B1(n_162), .B2(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_51), .B(n_324), .Y(n_392) );
OA22x2_ASAP7_75t_L g96 ( .A1(n_52), .A2(n_55), .B1(n_91), .B2(n_95), .Y(n_96) );
INVx1_ASAP7_75t_L g132 ( .A(n_52), .Y(n_132) );
INVx1_ASAP7_75t_L g108 ( .A(n_54), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_54), .B(n_130), .Y(n_150) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_54), .Y(n_187) );
OAI21xp33_ASAP7_75t_L g133 ( .A1(n_55), .A2(n_60), .B(n_134), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_56), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_57), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_58), .B(n_235), .Y(n_328) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_59), .Y(n_174) );
INVx1_ASAP7_75t_L g94 ( .A(n_60), .Y(n_94) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_60), .B(n_73), .Y(n_148) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_63), .Y(n_208) );
INVx1_ASAP7_75t_L g233 ( .A(n_63), .Y(n_233) );
BUFx5_ASAP7_75t_L g278 ( .A(n_63), .Y(n_278) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_65), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_65), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g391 ( .A(n_67), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_69), .Y(n_395) );
INVx2_ASAP7_75t_L g314 ( .A(n_70), .Y(n_314) );
INVx2_ASAP7_75t_SL g193 ( .A(n_71), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_72), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_73), .B(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_74), .A2(n_82), .B1(n_165), .B2(n_626), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_74), .Y(n_626) );
AO32x2_ASAP7_75t_L g273 ( .A1(n_76), .A2(n_198), .A3(n_269), .B1(n_274), .B2(n_281), .Y(n_273) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_76), .A2(n_274), .B1(n_415), .B2(n_417), .Y(n_414) );
AOI221xp5_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_179), .B1(n_196), .B2(n_209), .C(n_618), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_166), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_82), .B1(n_164), .B2(n_165), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_80), .Y(n_164) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g165 ( .A(n_82), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_82), .A2(n_165), .B1(n_620), .B2(n_621), .Y(n_619) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND3xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_136), .C(n_152), .Y(n_84) );
AND4x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_112), .C(n_122), .D(n_126), .Y(n_85) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x4_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g153 ( .A(n_88), .B(n_117), .Y(n_153) );
AND2x2_ASAP7_75t_L g162 ( .A(n_88), .B(n_120), .Y(n_162) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
INVx1_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
NAND2xp33_ASAP7_75t_L g90 ( .A(n_91), .B(n_92), .Y(n_90) );
INVx2_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx3_ASAP7_75t_L g100 ( .A(n_91), .Y(n_100) );
NAND2xp33_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_92), .B(n_132), .Y(n_131) );
INVxp67_ASAP7_75t_L g188 ( .A(n_92), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_94), .B(n_95), .Y(n_93) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_94), .A2(n_134), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g116 ( .A(n_96), .Y(n_116) );
AND2x2_ASAP7_75t_L g139 ( .A(n_96), .B(n_115), .Y(n_139) );
AND2x2_ASAP7_75t_L g158 ( .A(n_96), .B(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g123 ( .A(n_97), .B(n_114), .Y(n_123) );
AND2x4_ASAP7_75t_L g127 ( .A(n_97), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_102), .Y(n_97) );
OR2x2_ASAP7_75t_L g111 ( .A(n_98), .B(n_103), .Y(n_111) );
AND2x4_ASAP7_75t_L g117 ( .A(n_98), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g121 ( .A(n_98), .Y(n_121) );
AND2x2_ASAP7_75t_L g155 ( .A(n_98), .B(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_101), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_100), .B(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g130 ( .A(n_100), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g149 ( .A(n_101), .B(n_129), .C(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g118 ( .A(n_104), .Y(n_118) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AND2x4_ASAP7_75t_L g135 ( .A(n_110), .B(n_128), .Y(n_135) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g125 ( .A(n_111), .Y(n_125) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
AND2x4_ASAP7_75t_L g119 ( .A(n_114), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g124 ( .A(n_114), .B(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x4_ASAP7_75t_L g140 ( .A(n_117), .B(n_139), .Y(n_140) );
AND2x4_ASAP7_75t_L g120 ( .A(n_118), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g138 ( .A(n_120), .B(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g163 ( .A(n_120), .B(n_128), .Y(n_163) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_151), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_145), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_158), .Y(n_154) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_172), .B1(n_177), .B2(n_178), .Y(n_166) );
INVx1_ASAP7_75t_L g177 ( .A(n_167), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_168), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_172), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B1(n_175), .B2(n_176), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g176 ( .A(n_175), .Y(n_176) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_190), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g623 ( .A(n_183), .B(n_190), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .C(n_189), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_194), .Y(n_190) );
OR2x2_ASAP7_75t_L g628 ( .A(n_191), .B(n_195), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_191), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_191), .B(n_194), .Y(n_632) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g223 ( .A(n_199), .B(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g319 ( .A(n_199), .Y(n_319) );
AND2x2_ASAP7_75t_L g415 ( .A(n_199), .B(n_416), .Y(n_415) );
OA21x2_ASAP7_75t_L g630 ( .A1(n_200), .A2(n_631), .B(n_632), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_205), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_202), .B(n_261), .Y(n_306) );
INVx4_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_203), .A2(n_275), .B1(n_276), .B2(n_280), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_203), .A2(n_355), .B(n_357), .Y(n_354) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
INVx3_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
INVx4_ASAP7_75t_L g255 ( .A(n_204), .Y(n_255) );
INVx1_ASAP7_75t_L g348 ( .A(n_204), .Y(n_348) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
INVxp67_ASAP7_75t_SL g346 ( .A(n_207), .Y(n_346) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g235 ( .A(n_208), .Y(n_235) );
INVx6_ASAP7_75t_L g242 ( .A(n_208), .Y(n_242) );
INVx2_ASAP7_75t_L g302 ( .A(n_208), .Y(n_302) );
INVxp33_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_512), .Y(n_213) );
NAND3xp33_ASAP7_75t_L g214 ( .A(n_215), .B(n_409), .C(n_464), .Y(n_214) );
AOI211xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_288), .B(n_377), .C(n_407), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_284), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_272), .Y(n_218) );
AND2x4_ASAP7_75t_L g470 ( .A(n_219), .B(n_434), .Y(n_470) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g412 ( .A(n_220), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_248), .Y(n_220) );
OR2x2_ASAP7_75t_L g286 ( .A(n_221), .B(n_248), .Y(n_286) );
AND2x2_ASAP7_75t_L g463 ( .A(n_221), .B(n_414), .Y(n_463) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g382 ( .A(n_222), .Y(n_382) );
INVx1_ASAP7_75t_L g439 ( .A(n_222), .Y(n_439) );
AOI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_245), .Y(n_222) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_225), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
BUFx3_ASAP7_75t_L g312 ( .A(n_227), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B1(n_238), .B2(n_243), .Y(n_229) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g298 ( .A(n_232), .Y(n_298) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g240 ( .A(n_233), .Y(n_240) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g279 ( .A(n_235), .Y(n_279) );
INVx1_ASAP7_75t_L g337 ( .A(n_235), .Y(n_337) );
INVx1_ASAP7_75t_L g356 ( .A(n_235), .Y(n_356) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_237), .A2(n_321), .B(n_322), .C(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_237), .B(n_339), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_237), .A2(n_298), .B(n_391), .C(n_392), .Y(n_390) );
INVx3_ASAP7_75t_L g265 ( .A(n_239), .Y(n_265) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g324 ( .A(n_240), .Y(n_324) );
INVx1_ASAP7_75t_L g387 ( .A(n_241), .Y(n_387) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g252 ( .A(n_242), .Y(n_252) );
INVx2_ASAP7_75t_SL g267 ( .A(n_242), .Y(n_267) );
INVx2_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_243), .B(n_261), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_243), .B(n_261), .C(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_244), .A2(n_326), .B(n_327), .C(n_328), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_244), .A2(n_387), .B(n_388), .C(n_389), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
BUFx3_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_247), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g352 ( .A(n_247), .Y(n_352) );
INVx1_ASAP7_75t_L g396 ( .A(n_248), .Y(n_396) );
INVx2_ASAP7_75t_L g402 ( .A(n_248), .Y(n_402) );
AND2x2_ASAP7_75t_L g424 ( .A(n_248), .B(n_418), .Y(n_424) );
AND2x2_ASAP7_75t_L g433 ( .A(n_248), .B(n_384), .Y(n_433) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_263), .A3(n_269), .B(n_270), .Y(n_248) );
AOI221x1_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B1(n_257), .B2(n_259), .C(n_261), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g257 ( .A(n_254), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_255), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g417 ( .A(n_269), .Y(n_417) );
INVx2_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
AND2x2_ASAP7_75t_L g423 ( .A(n_272), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g457 ( .A(n_272), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g535 ( .A(n_272), .B(n_438), .Y(n_535) );
AND2x2_ASAP7_75t_L g588 ( .A(n_272), .B(n_433), .Y(n_588) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_272), .B(n_383), .Y(n_604) );
BUFx3_ASAP7_75t_L g614 ( .A(n_272), .Y(n_614) );
BUFx8_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g400 ( .A(n_273), .Y(n_400) );
AND2x2_ASAP7_75t_L g504 ( .A(n_273), .B(n_505), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_277), .A2(n_308), .B1(n_309), .B2(n_310), .Y(n_307) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g327 ( .A(n_278), .Y(n_327) );
INVx2_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
INVx2_ASAP7_75t_L g358 ( .A(n_278), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_278), .Y(n_362) );
INVx1_ASAP7_75t_L g321 ( .A(n_279), .Y(n_321) );
INVxp67_ASAP7_75t_L g376 ( .A(n_281), .Y(n_376) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_282), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g330 ( .A(n_283), .Y(n_330) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_283), .B(n_319), .Y(n_339) );
BUFx3_ASAP7_75t_L g341 ( .A(n_283), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_283), .B(n_319), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_283), .B(n_319), .Y(n_393) );
INVx1_ASAP7_75t_L g416 ( .A(n_283), .Y(n_416) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND3xp33_ASAP7_75t_SL g599 ( .A(n_285), .B(n_600), .C(n_603), .Y(n_599) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g478 ( .A(n_286), .Y(n_478) );
NAND2x1_ASAP7_75t_L g288 ( .A(n_289), .B(n_367), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_289), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_332), .Y(n_290) );
INVx1_ASAP7_75t_L g425 ( .A(n_291), .Y(n_425) );
AND2x2_ASAP7_75t_L g555 ( .A(n_291), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g593 ( .A(n_291), .B(n_446), .Y(n_593) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_315), .Y(n_291) );
OR2x2_ASAP7_75t_L g460 ( .A(n_292), .B(n_374), .Y(n_460) );
AND2x2_ASAP7_75t_L g547 ( .A(n_292), .B(n_421), .Y(n_547) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g448 ( .A(n_293), .B(n_406), .Y(n_448) );
BUFx2_ASAP7_75t_L g452 ( .A(n_293), .Y(n_452) );
OR2x2_ASAP7_75t_L g469 ( .A(n_293), .B(n_317), .Y(n_469) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_311), .B(n_313), .Y(n_293) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_294), .A2(n_313), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_305), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_300), .B2(n_303), .Y(n_295) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_309), .B(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g499 ( .A(n_316), .B(n_350), .Y(n_499) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
INVx2_ASAP7_75t_L g406 ( .A(n_317), .Y(n_406) );
AND2x2_ASAP7_75t_L g480 ( .A(n_317), .B(n_375), .Y(n_480) );
INVx1_ASAP7_75t_L g532 ( .A(n_317), .Y(n_532) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_317), .Y(n_566) );
AO31x2_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .A3(n_325), .B(n_329), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_330), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_332), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g484 ( .A(n_332), .B(n_480), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_332), .B(n_452), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_332), .B(n_451), .Y(n_615) );
NAND2xp67_ASAP7_75t_L g616 ( .A(n_332), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_349), .Y(n_332) );
INVx1_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
INVx2_ASAP7_75t_L g421 ( .A(n_333), .Y(n_421) );
INVx1_ASAP7_75t_L g429 ( .A(n_333), .Y(n_429) );
AND2x2_ASAP7_75t_L g491 ( .A(n_333), .B(n_350), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_334), .B(n_342), .Y(n_333) );
AND2x2_ASAP7_75t_SL g528 ( .A(n_334), .B(n_342), .Y(n_528) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .B(n_340), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_339), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_347), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g431 ( .A(n_349), .B(n_375), .Y(n_431) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g374 ( .A(n_350), .Y(n_374) );
INVx1_ASAP7_75t_L g455 ( .A(n_350), .Y(n_455) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_350), .Y(n_523) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_359), .B(n_366), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B(n_363), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_368), .A2(n_561), .B1(n_563), .B2(n_565), .Y(n_560) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_373), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
BUFx3_ASAP7_75t_L g475 ( .A(n_370), .Y(n_475) );
AND2x2_ASAP7_75t_L g522 ( .A(n_371), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AND2x2_ASAP7_75t_L g531 ( .A(n_374), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_397), .B(n_403), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_378), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
AND2x4_ASAP7_75t_L g398 ( .A(n_380), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_380), .B(n_413), .Y(n_533) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g489 ( .A(n_381), .B(n_383), .Y(n_489) );
INVx2_ASAP7_75t_L g540 ( .A(n_381), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_381), .B(n_424), .Y(n_594) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g505 ( .A(n_382), .Y(n_505) );
INVx2_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx2_ASAP7_75t_L g458 ( .A(n_383), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_383), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_383), .B(n_448), .Y(n_551) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_396), .Y(n_383) );
INVx2_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
INVx1_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
BUFx3_ASAP7_75t_L g472 ( .A(n_384), .Y(n_472) );
AND2x4_ASAP7_75t_L g542 ( .A(n_384), .B(n_400), .Y(n_542) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AO31x2_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_390), .A3(n_393), .B(n_394), .Y(n_385) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g488 ( .A(n_399), .Y(n_488) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_400), .B(n_505), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_401), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g438 ( .A(n_402), .B(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
INVx1_ASAP7_75t_L g564 ( .A(n_402), .Y(n_564) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp67_ASAP7_75t_L g494 ( .A(n_405), .B(n_460), .Y(n_494) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g510 ( .A(n_406), .B(n_497), .Y(n_510) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_406), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_426), .C(n_435), .Y(n_409) );
OAI22xp33_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_419), .B1(n_422), .B2(n_425), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx2_ASAP7_75t_L g585 ( .A(n_412), .Y(n_585) );
AND2x4_ASAP7_75t_L g477 ( .A(n_413), .B(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g493 ( .A(n_413), .Y(n_493) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
INVx1_ASAP7_75t_L g442 ( .A(n_414), .Y(n_442) );
AND2x4_ASAP7_75t_L g471 ( .A(n_414), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g483 ( .A(n_418), .B(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_420), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g583 ( .A(n_420), .B(n_499), .Y(n_583) );
BUFx2_ASAP7_75t_L g446 ( .A(n_421), .Y(n_446) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_421), .Y(n_572) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_423), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g503 ( .A(n_424), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g543 ( .A(n_424), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g578 ( .A(n_424), .B(n_497), .Y(n_578) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .Y(n_426) );
INVx3_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
AND2x2_ASAP7_75t_L g525 ( .A(n_428), .B(n_480), .Y(n_525) );
INVx1_ASAP7_75t_L g607 ( .A(n_428), .Y(n_607) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g498 ( .A(n_429), .B(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g508 ( .A(n_431), .Y(n_508) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_431), .Y(n_573) );
OR2x6_ASAP7_75t_L g609 ( .A(n_431), .B(n_610), .Y(n_609) );
OAI31xp33_ASAP7_75t_L g524 ( .A1(n_432), .A2(n_444), .A3(n_525), .B(n_526), .Y(n_524) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_L g519 ( .A(n_433), .Y(n_519) );
INVx2_ASAP7_75t_L g602 ( .A(n_433), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_443), .B(n_449), .Y(n_435) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_438), .Y(n_612) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_439), .Y(n_474) );
INVx2_ASAP7_75t_L g497 ( .A(n_439), .Y(n_497) );
AOI33xp33_ASAP7_75t_L g492 ( .A1(n_440), .A2(n_493), .A3(n_494), .B1(n_495), .B2(n_496), .B3(n_498), .Y(n_492) );
AND2x2_ASAP7_75t_L g559 ( .A(n_440), .B(n_497), .Y(n_559) );
AND2x2_ASAP7_75t_L g561 ( .A(n_440), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
NOR2x1p5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g479 ( .A(n_446), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g473 ( .A(n_448), .B(n_474), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_448), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g597 ( .A(n_448), .B(n_491), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_456), .B1(n_459), .B2(n_461), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g517 ( .A(n_452), .B(n_491), .Y(n_517) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_454), .B(n_475), .Y(n_549) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g556 ( .A(n_455), .B(n_528), .Y(n_556) );
AND2x2_ASAP7_75t_L g590 ( .A(n_455), .B(n_528), .Y(n_590) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp67_ASAP7_75t_SL g526 ( .A(n_460), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_L g550 ( .A(n_463), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_485), .C(n_500), .Y(n_464) );
OAI21xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_475), .B(n_476), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_470), .B1(n_471), .B2(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g617 ( .A(n_469), .Y(n_617) );
INVx2_ASAP7_75t_L g568 ( .A(n_471), .Y(n_568) );
INVx1_ASAP7_75t_L g601 ( .A(n_474), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_479), .B1(n_481), .B2(n_484), .Y(n_476) );
AND2x2_ASAP7_75t_L g490 ( .A(n_480), .B(n_491), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_481), .A2(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g511 ( .A(n_491), .Y(n_511) );
AND2x2_ASAP7_75t_L g565 ( .A(n_491), .B(n_566), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_493), .B(n_510), .C(n_511), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_493), .A2(n_554), .B1(n_557), .B2(n_558), .C(n_560), .Y(n_553) );
INVx2_ASAP7_75t_L g515 ( .A(n_495), .Y(n_515) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
BUFx3_ASAP7_75t_L g587 ( .A(n_497), .Y(n_587) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_547), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_506), .B(n_509), .Y(n_502) );
AND2x4_ASAP7_75t_SL g563 ( .A(n_504), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_513), .B(n_552), .C(n_580), .D(n_598), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_529), .Y(n_513) );
OAI221xp5_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_516), .B1(n_518), .B2(n_521), .C(n_524), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g544 ( .A(n_520), .Y(n_544) );
INVx1_ASAP7_75t_L g575 ( .A(n_520), .Y(n_575) );
INVxp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g546 ( .A(n_523), .Y(n_546) );
INVx1_ASAP7_75t_SL g557 ( .A(n_525), .Y(n_557) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g537 ( .A(n_528), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_533), .B1(n_534), .B2(n_536), .C(n_538), .Y(n_529) );
AND2x2_ASAP7_75t_L g589 ( .A(n_532), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g579 ( .A(n_536), .Y(n_579) );
O2A1O1Ixp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_543), .B(n_545), .C(n_548), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B(n_551), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_567), .Y(n_552) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_574), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_578), .B2(n_579), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B1(n_586), .B2(n_589), .C(n_591), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_594), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_605), .B1(n_611), .B2(n_613), .Y(n_598) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_616), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B1(n_624), .B2(n_627), .C1(n_629), .C2(n_633), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_620), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
endmodule