module fake_netlist_6_4802_n_1233 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1233);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1233;

wire n_992;
wire n_801;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_653;
wire n_236;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;

INVx1_ASAP7_75t_L g175 ( 
.A(n_16),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_34),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_29),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_67),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_25),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_38),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_42),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_38),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_39),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_20),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_40),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_86),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_158),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_87),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_50),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_99),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_48),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_57),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_152),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_151),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_25),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_15),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_97),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_64),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_62),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_50),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_149),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_14),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_144),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_154),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_102),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_164),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_168),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_153),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_103),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_163),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_66),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_10),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_55),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_43),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_116),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_112),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_84),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_59),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_65),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_123),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_26),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_76),
.Y(n_265)
);

BUFx2_ASAP7_75t_R g266 ( 
.A(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_174),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_117),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_166),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_150),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_52),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_169),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_171),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_119),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_19),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_98),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_18),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_45),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_165),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_139),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_159),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_104),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_56),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_130),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_71),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_20),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_37),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_46),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_17),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_213),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_189),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_176),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_213),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_191),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_180),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_197),
.B(n_0),
.Y(n_305)
);

INVx4_ASAP7_75t_R g306 ( 
.A(n_238),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_281),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_183),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_190),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_244),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_175),
.Y(n_317)
);

BUFx6f_ASAP7_75t_SL g318 ( 
.A(n_238),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_195),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_204),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_190),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_198),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_192),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_217),
.B(n_0),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_205),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_252),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_211),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_251),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_216),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_252),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_219),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_197),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_249),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_1),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_249),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_221),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_278),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_222),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_227),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_237),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_264),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_273),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_273),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_209),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_274),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_274),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_287),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_295),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_182),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_289),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_177),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_184),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_251),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_178),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_187),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_196),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_255),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_214),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_223),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_255),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_224),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_225),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_181),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_292),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_185),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_226),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_206),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_234),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_240),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_247),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_250),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_188),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_257),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_276),
.B(n_179),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_229),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_186),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_199),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_209),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_325),
.A2(n_229),
.B1(n_232),
.B2(n_231),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_188),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_193),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_303),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_193),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_338),
.B(n_209),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_306),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_194),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_179),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_243),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_265),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_299),
.B(n_194),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_235),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_332),
.B(n_265),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_296),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_298),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_307),
.B(n_266),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_305),
.B(n_260),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_335),
.B(n_302),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_324),
.Y(n_435)
);

AND2x4_ASAP7_75t_SL g436 ( 
.A(n_358),
.B(n_232),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_300),
.B(n_209),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_304),
.B(n_270),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_381),
.B(n_235),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_321),
.B(n_275),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_361),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_300),
.B(n_209),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_318),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_381),
.B(n_312),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_311),
.B(n_242),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_299),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_311),
.B(n_242),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_371),
.B(n_282),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_318),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_330),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_320),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_320),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_329),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_329),
.B(n_200),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_331),
.B(n_291),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_394),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_402),
.B(n_432),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_331),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_426),
.A2(n_312),
.B1(n_215),
.B2(n_230),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_261),
.B1(n_215),
.B2(n_230),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_402),
.B(n_333),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_402),
.A2(n_453),
.B1(n_452),
.B2(n_439),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_445),
.B(n_333),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_370),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_443),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_L g482 ( 
.A1(n_389),
.A2(n_434),
.B1(n_454),
.B2(n_450),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_389),
.B(n_342),
.C(n_340),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

NOR2x1p5_ASAP7_75t_L g486 ( 
.A(n_449),
.B(n_360),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_426),
.A2(n_215),
.B1(n_230),
.B2(n_261),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_447),
.B(n_340),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_452),
.A2(n_386),
.B1(n_385),
.B2(n_373),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_441),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_426),
.B(n_342),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_436),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_447),
.B(n_344),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_398),
.A2(n_375),
.B1(n_286),
.B2(n_284),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_416),
.B(n_344),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_416),
.B(n_345),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_453),
.B(n_345),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_387),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_444),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_416),
.B(n_346),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_393),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_454),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_439),
.B(n_455),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_346),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_451),
.A2(n_364),
.B1(n_367),
.B2(n_372),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_444),
.B(n_384),
.C(n_380),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

AND3x1_ASAP7_75t_L g522 ( 
.A(n_454),
.B(n_432),
.C(n_440),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_393),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_398),
.A2(n_261),
.B1(n_215),
.B2(n_230),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_494),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_527),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_514),
.B(n_451),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_457),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_500),
.A2(n_448),
.B1(n_440),
.B2(n_425),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_492),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_451),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_476),
.B(n_425),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_476),
.B(n_440),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_467),
.A2(n_442),
.B(n_437),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_522),
.A2(n_434),
.B1(n_451),
.B2(n_442),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_483),
.B(n_513),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_483),
.B(n_455),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_503),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_513),
.B(n_456),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_446),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_483),
.B(n_448),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_474),
.A2(n_456),
.B1(n_448),
.B2(n_437),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_477),
.B(n_423),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_477),
.B(n_480),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_502),
.B(n_446),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_462),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_466),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_423),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_480),
.B(n_438),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_485),
.B(n_438),
.Y(n_560)
);

BUFx5_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_503),
.B(n_449),
.Y(n_562)
);

O2A1O1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_482),
.A2(n_390),
.B(n_392),
.C(n_396),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_466),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_485),
.B(n_438),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_527),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_516),
.B(n_411),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_490),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_493),
.B(n_435),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_522),
.B(n_411),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_411),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_493),
.B(n_435),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_478),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_518),
.A2(n_424),
.B(n_392),
.C(n_396),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_518),
.B(n_408),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_472),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_525),
.B(n_215),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_500),
.A2(n_433),
.B1(n_415),
.B2(n_408),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_488),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_500),
.B(n_408),
.Y(n_583)
);

BUFx8_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_459),
.B(n_411),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_470),
.B(n_436),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_413),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_500),
.A2(n_433),
.B1(n_415),
.B2(n_413),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_517),
.B(n_411),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_488),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_470),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_469),
.B(n_411),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_489),
.B(n_347),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_495),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_498),
.A2(n_417),
.B1(n_433),
.B2(n_406),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_463),
.A2(n_433),
.B1(n_415),
.B2(n_413),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_471),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_465),
.B(n_347),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_506),
.B(n_353),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_524),
.B(n_421),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_478),
.A2(n_390),
.B(n_406),
.C(n_424),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_520),
.B(n_354),
.C(n_353),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_464),
.B(n_354),
.C(n_364),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_527),
.B(n_411),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_471),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_487),
.A2(n_367),
.B1(n_372),
.B2(n_297),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_486),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_497),
.B(n_301),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_486),
.B(n_436),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_499),
.B(n_308),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_499),
.B(n_315),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_495),
.B(n_310),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_509),
.B(n_323),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_521),
.A2(n_433),
.B1(n_246),
.B2(n_263),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_521),
.B(n_337),
.Y(n_623)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_509),
.B(n_411),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_509),
.B(n_415),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_537),
.A2(n_515),
.B(n_512),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_574),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_430),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_578),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_537),
.A2(n_515),
.B(n_512),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_552),
.A2(n_339),
.B1(n_357),
.B2(n_355),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_532),
.B(n_521),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_546),
.A2(n_515),
.B(n_512),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_543),
.A2(n_351),
.B1(n_352),
.B2(n_526),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_593),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_536),
.B(n_283),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_575),
.A2(n_523),
.B(n_496),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_543),
.B(n_547),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_528),
.A2(n_526),
.B(n_519),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_545),
.A2(n_526),
.B(n_519),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_539),
.A2(n_290),
.B1(n_523),
.B2(n_473),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_554),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_554),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_620),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_533),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_574),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_558),
.A2(n_519),
.B(n_501),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_539),
.A2(n_523),
.B1(n_473),
.B2(n_496),
.Y(n_649)
);

AOI21x1_ASAP7_75t_L g650 ( 
.A1(n_567),
.A2(n_481),
.B(n_415),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_540),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_544),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_551),
.B(n_473),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_473),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_548),
.A2(n_519),
.B(n_501),
.Y(n_656)
);

AOI211xp5_ASAP7_75t_L g657 ( 
.A1(n_614),
.A2(n_429),
.B(n_427),
.C(n_405),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_607),
.B(n_407),
.C(n_405),
.Y(n_658)
);

AOI22x1_ASAP7_75t_L g659 ( 
.A1(n_549),
.A2(n_496),
.B1(n_505),
.B2(n_481),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_579),
.B(n_430),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_625),
.A2(n_505),
.B(n_496),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_550),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_563),
.B(n_505),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_603),
.B(n_407),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_531),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_538),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_556),
.B(n_557),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_542),
.A2(n_597),
.B1(n_562),
.B2(n_595),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_606),
.A2(n_505),
.B(n_481),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_564),
.Y(n_670)
);

OAI321xp33_ASAP7_75t_L g671 ( 
.A1(n_614),
.A2(n_427),
.A3(n_414),
.B1(n_429),
.B2(n_412),
.C(n_422),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_621),
.B(n_430),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_553),
.A2(n_501),
.B(n_475),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_625),
.A2(n_501),
.B(n_475),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_573),
.B(n_421),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_577),
.B(n_421),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_541),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_559),
.B(n_421),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_618),
.B(n_619),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_559),
.B(n_458),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_553),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_574),
.B(n_475),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_576),
.A2(n_475),
.B(n_458),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_602),
.A2(n_272),
.B1(n_202),
.B2(n_203),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_560),
.B(n_458),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_576),
.A2(n_475),
.B(n_458),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_560),
.A2(n_475),
.B(n_458),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_600),
.Y(n_688)
);

NOR2x1p5_ASAP7_75t_SL g689 ( 
.A(n_561),
.B(n_610),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_550),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_568),
.B(n_623),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_565),
.A2(n_507),
.B(n_504),
.Y(n_692)
);

BUFx4f_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_565),
.A2(n_409),
.B(n_403),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_616),
.B(n_412),
.Y(n_695)
);

AOI21xp33_ASAP7_75t_L g696 ( 
.A1(n_583),
.A2(n_589),
.B(n_534),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_583),
.A2(n_261),
.B1(n_230),
.B2(n_403),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_605),
.A2(n_507),
.B(n_504),
.Y(n_698)
);

AO21x1_ASAP7_75t_L g699 ( 
.A1(n_589),
.A2(n_422),
.B(n_414),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_569),
.B(n_572),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_570),
.A2(n_591),
.B(n_594),
.C(n_585),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_572),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_608),
.B(n_431),
.Y(n_703)
);

O2A1O1Ixp5_ASAP7_75t_L g704 ( 
.A1(n_611),
.A2(n_431),
.B(n_418),
.C(n_403),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_601),
.B(n_587),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_622),
.A2(n_590),
.B(n_581),
.C(n_609),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_615),
.B(n_588),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_598),
.B(n_504),
.Y(n_709)
);

NOR2x1p5_ASAP7_75t_SL g710 ( 
.A(n_561),
.B(n_409),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_538),
.B(n_504),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_584),
.Y(n_712)
);

CKINVDCx10_ASAP7_75t_R g713 ( 
.A(n_529),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_586),
.A2(n_507),
.B(n_504),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_592),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_596),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_599),
.A2(n_507),
.B(n_504),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_617),
.A2(n_587),
.B1(n_604),
.B2(n_601),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_538),
.B(n_507),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_612),
.A2(n_418),
.B(n_409),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_604),
.B(n_561),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_646),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_628),
.B(n_631),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_679),
.B(n_535),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_664),
.A2(n_571),
.B(n_431),
.C(n_419),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_699),
.A2(n_419),
.B(n_420),
.C(n_418),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_665),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_627),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_670),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_691),
.A2(n_566),
.B1(n_529),
.B2(n_201),
.Y(n_732)
);

AOI21x1_ASAP7_75t_L g733 ( 
.A1(n_663),
.A2(n_624),
.B(n_401),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_666),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_695),
.B(n_566),
.Y(n_735)
);

NAND2x1p5_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_627),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_677),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_635),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_666),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_707),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_700),
.B(n_566),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_636),
.A2(n_419),
.B(n_420),
.C(n_428),
.Y(n_742)
);

O2A1O1Ixp5_ASAP7_75t_L g743 ( 
.A1(n_638),
.A2(n_637),
.B(n_669),
.C(n_701),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_652),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_702),
.A2(n_685),
.B(n_680),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_713),
.B(n_693),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_688),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_SL g748 ( 
.A1(n_706),
.A2(n_420),
.B(n_401),
.C(n_428),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_642),
.A2(n_428),
.B(n_561),
.C(n_580),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_645),
.B(n_584),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_716),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_634),
.B(n_561),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_671),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_643),
.B(n_613),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_641),
.B(n_613),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_668),
.A2(n_708),
.B1(n_672),
.B2(n_718),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_627),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_673),
.A2(n_613),
.B(n_561),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_678),
.A2(n_511),
.B(n_507),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_660),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_709),
.A2(n_511),
.B(n_261),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_644),
.B(n_207),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_696),
.A2(n_580),
.B1(n_259),
.B2(n_258),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_681),
.B(n_208),
.Y(n_765)
);

AO32x1_ASAP7_75t_L g766 ( 
.A1(n_649),
.A2(n_580),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_629),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_667),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_657),
.B(n_210),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_697),
.A2(n_580),
.B1(n_267),
.B2(n_262),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_654),
.A2(n_511),
.B(n_268),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_647),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_703),
.B(n_212),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_662),
.A2(n_218),
.B1(n_220),
.B2(n_228),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_658),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_647),
.B(n_233),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_641),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_690),
.B(n_236),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_711),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_R g781 ( 
.A(n_641),
.B(n_239),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_684),
.B(n_241),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_655),
.B(n_245),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_659),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_662),
.B(n_705),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_648),
.A2(n_511),
.B(n_288),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_725),
.A2(n_692),
.A3(n_698),
.B(n_639),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_761),
.B(n_712),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_745),
.A2(n_721),
.B(n_692),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_738),
.Y(n_790)
);

AOI221x1_ASAP7_75t_L g791 ( 
.A1(n_762),
.A2(n_633),
.B1(n_698),
.B2(n_630),
.C(n_626),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_741),
.A2(n_656),
.B(n_640),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_759),
.A2(n_694),
.B(n_633),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_743),
.A2(n_719),
.B(n_683),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_735),
.A2(n_682),
.B1(n_632),
.B2(n_277),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_733),
.A2(n_753),
.B(n_760),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_743),
.A2(n_626),
.B(n_630),
.Y(n_797)
);

AO22x2_ASAP7_75t_L g798 ( 
.A1(n_723),
.A2(n_661),
.B1(n_717),
.B2(n_714),
.Y(n_798)
);

BUFx12f_ASAP7_75t_L g799 ( 
.A(n_744),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_750),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_735),
.A2(n_683),
.B(n_686),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_722),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_730),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_769),
.A2(n_757),
.B1(n_764),
.B2(n_771),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_786),
.A2(n_686),
.B(n_674),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_761),
.B(n_661),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_731),
.Y(n_807)
);

AO31x2_ASAP7_75t_L g808 ( 
.A1(n_784),
.A2(n_717),
.A3(n_714),
.B(n_676),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_750),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_755),
.A2(n_674),
.B(n_687),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_778),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_724),
.B(n_768),
.Y(n_812)
);

OAI22x1_ASAP7_75t_L g813 ( 
.A1(n_785),
.A2(n_650),
.B1(n_269),
.B2(n_279),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_727),
.A2(n_704),
.B(n_687),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_755),
.A2(n_675),
.B(n_720),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_727),
.A2(n_689),
.B(n_710),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_782),
.A2(n_256),
.B1(n_285),
.B2(n_511),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_749),
.A2(n_580),
.B(n_388),
.Y(n_818)
);

NOR2x1_ASAP7_75t_SL g819 ( 
.A(n_756),
.B(n_729),
.Y(n_819)
);

AO22x2_ASAP7_75t_L g820 ( 
.A1(n_740),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_779),
.B(n_8),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_751),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_729),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_729),
.Y(n_824)
);

AOI21x1_ASAP7_75t_L g825 ( 
.A1(n_772),
.A2(n_783),
.B(n_765),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_763),
.A2(n_511),
.B1(n_393),
.B2(n_397),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_779),
.A2(n_388),
.B1(n_397),
.B2(n_399),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_749),
.A2(n_388),
.B(n_393),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_748),
.A2(n_742),
.B(n_764),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_777),
.A2(n_393),
.B(n_397),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_774),
.B(n_9),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_10),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_754),
.A2(n_393),
.B(n_399),
.C(n_397),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_726),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_770),
.A2(n_399),
.B(n_397),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_773),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_729),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_732),
.A2(n_399),
.B1(n_12),
.B2(n_13),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_SL g839 ( 
.A1(n_776),
.A2(n_11),
.B(n_12),
.Y(n_839)
);

NAND2x1_ASAP7_75t_L g840 ( 
.A(n_767),
.B(n_399),
.Y(n_840)
);

OA21x2_ASAP7_75t_L g841 ( 
.A1(n_728),
.A2(n_399),
.B(n_388),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_804),
.A2(n_775),
.B1(n_747),
.B2(n_737),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_806),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_802),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_808),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_804),
.A2(n_771),
.B1(n_736),
.B2(n_756),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_838),
.A2(n_775),
.B1(n_781),
.B2(n_780),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_821),
.A2(n_831),
.B1(n_812),
.B2(n_788),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_839),
.A2(n_820),
.B1(n_832),
.B2(n_834),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_824),
.Y(n_850)
);

CKINVDCx16_ASAP7_75t_R g851 ( 
.A(n_799),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_820),
.A2(n_781),
.B1(n_780),
.B2(n_734),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_800),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_808),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_837),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_836),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_803),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_808),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_790),
.A2(n_780),
.B1(n_734),
.B2(n_739),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_811),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_816),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_807),
.B(n_780),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_816),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_798),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_SL g866 ( 
.A1(n_839),
.A2(n_736),
.B(n_746),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_800),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_795),
.A2(n_756),
.B1(n_767),
.B2(n_739),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_817),
.A2(n_809),
.B1(n_813),
.B2(n_829),
.Y(n_869)
);

CKINVDCx11_ASAP7_75t_R g870 ( 
.A(n_809),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_798),
.B(n_758),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_827),
.A2(n_758),
.B1(n_746),
.B2(n_766),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_819),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_841),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_787),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_758),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_823),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_SL g878 ( 
.A1(n_829),
.A2(n_758),
.B1(n_766),
.B2(n_14),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_801),
.B(n_11),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_SL g880 ( 
.A1(n_818),
.A2(n_766),
.B(n_15),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_797),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_810),
.A2(n_399),
.B1(n_388),
.B2(n_18),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_840),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_787),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_797),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_787),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_825),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_796),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_794),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_830),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_833),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_791),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_835),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_789),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_814),
.B(n_51),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_L g896 ( 
.A1(n_815),
.A2(n_13),
.B(n_17),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_826),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_805),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_845),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_865),
.Y(n_900)
);

INVx6_ASAP7_75t_L g901 ( 
.A(n_873),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_874),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_845),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_845),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_865),
.B(n_793),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_854),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_870),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_854),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_881),
.B(n_814),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_853),
.B(n_792),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_854),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_866),
.B(n_19),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_874),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_858),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_828),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_858),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_858),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_855),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_871),
.B(n_828),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_886),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_886),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_871),
.B(n_818),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_889),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_874),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_843),
.B(n_849),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_874),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_843),
.B(n_21),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_889),
.Y(n_929)
);

OA21x2_ASAP7_75t_L g930 ( 
.A1(n_892),
.A2(n_388),
.B(n_22),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_888),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_888),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_887),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_867),
.B(n_53),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_861),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_849),
.B(n_21),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_909),
.B(n_884),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_909),
.B(n_884),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_912),
.A2(n_896),
.B(n_847),
.C(n_869),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_936),
.A2(n_896),
.B(n_879),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_921),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_910),
.A2(n_894),
.B(n_891),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_935),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_931),
.Y(n_944)
);

AO22x2_ASAP7_75t_L g945 ( 
.A1(n_926),
.A2(n_892),
.B1(n_885),
.B2(n_881),
.Y(n_945)
);

INVx5_ASAP7_75t_SL g946 ( 
.A(n_915),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_875),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_909),
.B(n_919),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_935),
.B(n_875),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_933),
.B(n_935),
.Y(n_950)
);

OA21x2_ASAP7_75t_L g951 ( 
.A1(n_920),
.A2(n_885),
.B(n_898),
.Y(n_951)
);

OA21x2_ASAP7_75t_L g952 ( 
.A1(n_920),
.A2(n_893),
.B(n_895),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_912),
.A2(n_852),
.B(n_880),
.C(n_846),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_926),
.B(n_844),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_919),
.B(n_875),
.Y(n_955)
);

OA21x2_ASAP7_75t_L g956 ( 
.A1(n_922),
.A2(n_895),
.B(n_844),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_936),
.A2(n_872),
.B(n_891),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_933),
.B(n_875),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_901),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_934),
.A2(n_880),
.B(n_848),
.C(n_878),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_919),
.B(n_861),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_905),
.B(n_891),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_928),
.A2(n_882),
.B(n_856),
.C(n_842),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_928),
.A2(n_891),
.B1(n_897),
.B2(n_868),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_SL g965 ( 
.A1(n_930),
.A2(n_887),
.B1(n_873),
.B2(n_850),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_902),
.B(n_861),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_919),
.B(n_861),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_921),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_919),
.B(n_864),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_905),
.B(n_857),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_923),
.B(n_864),
.Y(n_971)
);

OA21x2_ASAP7_75t_L g972 ( 
.A1(n_922),
.A2(n_857),
.B(n_863),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_923),
.B(n_864),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_902),
.B(n_863),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_923),
.B(n_864),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_902),
.B(n_864),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_940),
.A2(n_905),
.B1(n_900),
.B2(n_923),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_972),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_941),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_SL g980 ( 
.A(n_957),
.B(n_924),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_941),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_972),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_954),
.B(n_931),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_954),
.B(n_932),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_941),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_972),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_972),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_948),
.B(n_921),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_948),
.B(n_904),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_961),
.B(n_904),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_961),
.B(n_904),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_939),
.A2(n_930),
.B1(n_918),
.B2(n_923),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_950),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_966),
.B(n_902),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_967),
.B(n_917),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_972),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_964),
.B(n_918),
.Y(n_997)
);

OAI222xp33_ASAP7_75t_L g998 ( 
.A1(n_964),
.A2(n_900),
.B1(n_915),
.B2(n_862),
.C1(n_853),
.C2(n_855),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_967),
.B(n_971),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_971),
.B(n_917),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_968),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_992),
.A2(n_940),
.B1(n_945),
.B2(n_946),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_982),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_979),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_992),
.A2(n_945),
.B1(n_953),
.B2(n_960),
.C(n_957),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_SL g1006 ( 
.A(n_997),
.B(n_963),
.C(n_965),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_979),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_979),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_946),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_988),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_997),
.A2(n_962),
.B1(n_887),
.B2(n_946),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_982),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_981),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_981),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_994),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_986),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_981),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_985),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_977),
.A2(n_962),
.B1(n_887),
.B2(n_946),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_985),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_977),
.A2(n_962),
.B1(n_946),
.B2(n_959),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_985),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1003),
.Y(n_1023)
);

INVxp33_ASAP7_75t_L g1024 ( 
.A(n_1009),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_1009),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1003),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1015),
.B(n_999),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1010),
.B(n_999),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1003),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1012),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_1006),
.B(n_907),
.Y(n_1031)
);

AND2x4_ASAP7_75t_SL g1032 ( 
.A(n_1011),
.B(n_974),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1012),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_994),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1031),
.A2(n_1005),
.B1(n_1002),
.B2(n_1019),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_1028),
.B(n_980),
.Y(n_1036)
);

OAI211xp5_ASAP7_75t_L g1037 ( 
.A1(n_1025),
.A2(n_965),
.B(n_1021),
.C(n_978),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_959),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1023),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_1027),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1035),
.B(n_1028),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_1040),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1039),
.Y(n_1043)
);

NAND4xp25_ASAP7_75t_L g1044 ( 
.A(n_1037),
.B(n_860),
.C(n_959),
.D(n_942),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1044),
.A2(n_1024),
.B1(n_1036),
.B2(n_1037),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1041),
.A2(n_851),
.B(n_1032),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1042),
.A2(n_1032),
.B1(n_1038),
.B2(n_1034),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1038),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1043),
.Y(n_1049)
);

OAI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_1044),
.A2(n_962),
.B1(n_987),
.B2(n_978),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1043),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1044),
.A2(n_945),
.B1(n_901),
.B2(n_962),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1043),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1043),
.Y(n_1054)
);

OAI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_1041),
.A2(n_901),
.B1(n_1030),
.B2(n_1026),
.C(n_1023),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1048),
.B(n_980),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1049),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_1045),
.B(n_851),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1051),
.Y(n_1059)
);

OAI221xp5_ASAP7_75t_L g1060 ( 
.A1(n_1046),
.A2(n_901),
.B1(n_1030),
.B2(n_1026),
.C(n_1033),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1053),
.B(n_853),
.C(n_1033),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1054),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1052),
.B(n_1029),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1052),
.B(n_1029),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1047),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1050),
.A2(n_998),
.B(n_860),
.C(n_987),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_1055),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1045),
.B(n_860),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1049),
.Y(n_1069)
);

OAI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1052),
.A2(n_996),
.B1(n_986),
.B2(n_993),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1048),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1057),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1059),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1058),
.A2(n_998),
.B(n_945),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1069),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1071),
.B(n_980),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1071),
.B(n_1065),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1062),
.B(n_1012),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1056),
.Y(n_1079)
);

AOI322xp5_ASAP7_75t_L g1080 ( 
.A1(n_1068),
.A2(n_996),
.A3(n_1016),
.B1(n_937),
.B2(n_993),
.C1(n_988),
.C2(n_989),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1063),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1067),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1067),
.B(n_994),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1070),
.B(n_853),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_SL g1085 ( 
.A1(n_1060),
.A2(n_1016),
.B(n_983),
.C(n_984),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_1061),
.B(n_22),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1064),
.B(n_994),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1066),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1057),
.B(n_1016),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1057),
.Y(n_1090)
);

NOR4xp25_ASAP7_75t_L g1091 ( 
.A(n_1082),
.B(n_1077),
.C(n_1073),
.D(n_1075),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1083),
.B(n_1081),
.Y(n_1092)
);

OAI221xp5_ASAP7_75t_L g1093 ( 
.A1(n_1074),
.A2(n_1088),
.B1(n_1079),
.B2(n_1086),
.C(n_1072),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_1076),
.B(n_23),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1090),
.B(n_859),
.C(n_942),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1089),
.B(n_23),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_1080),
.B(n_853),
.C(n_930),
.Y(n_1097)
);

AOI211xp5_ASAP7_75t_L g1098 ( 
.A1(n_1084),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1098)
);

OAI211xp5_ASAP7_75t_L g1099 ( 
.A1(n_1085),
.A2(n_853),
.B(n_930),
.C(n_983),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1089),
.A2(n_945),
.B(n_984),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1087),
.B(n_1004),
.Y(n_1101)
);

OAI211xp5_ASAP7_75t_L g1102 ( 
.A1(n_1078),
.A2(n_930),
.B(n_29),
.C(n_30),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1078),
.B(n_901),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1077),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1083),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1077),
.Y(n_1106)
);

AND4x1_ASAP7_75t_L g1107 ( 
.A(n_1077),
.B(n_28),
.C(n_30),
.D(n_31),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_1104),
.B(n_28),
.C(n_32),
.Y(n_1108)
);

OAI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1091),
.A2(n_958),
.B1(n_970),
.B2(n_1018),
.C(n_1017),
.Y(n_1109)
);

NOR3xp33_ASAP7_75t_SL g1110 ( 
.A(n_1093),
.B(n_32),
.C(n_33),
.Y(n_1110)
);

OAI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1091),
.A2(n_1022),
.B1(n_1020),
.B2(n_1018),
.C(n_1017),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1092),
.A2(n_33),
.B(n_35),
.Y(n_1112)
);

OAI211xp5_ASAP7_75t_L g1113 ( 
.A1(n_1098),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1113)
);

OAI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1106),
.A2(n_36),
.B(n_41),
.C(n_43),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1094),
.B(n_1004),
.Y(n_1115)
);

AOI321xp33_ASAP7_75t_L g1116 ( 
.A1(n_1105),
.A2(n_41),
.A3(n_44),
.B1(n_45),
.B2(n_46),
.C(n_47),
.Y(n_1116)
);

OAI211xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1103),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1097),
.A2(n_1022),
.B1(n_1020),
.B2(n_1013),
.C(n_1014),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1096),
.Y(n_1119)
);

AOI221xp5_ASAP7_75t_L g1120 ( 
.A1(n_1099),
.A2(n_1013),
.B1(n_1014),
.B2(n_1008),
.C(n_1007),
.Y(n_1120)
);

NOR4xp75_ASAP7_75t_L g1121 ( 
.A(n_1101),
.B(n_49),
.C(n_876),
.D(n_877),
.Y(n_1121)
);

NAND4xp25_ASAP7_75t_L g1122 ( 
.A(n_1100),
.B(n_910),
.C(n_850),
.D(n_876),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_1095),
.B(n_1102),
.C(n_1107),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1093),
.A2(n_1008),
.B1(n_1007),
.B2(n_49),
.C(n_944),
.Y(n_1124)
);

NOR4xp25_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_877),
.C(n_944),
.D(n_1001),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1091),
.A2(n_994),
.B(n_974),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1091),
.A2(n_974),
.B1(n_950),
.B2(n_1001),
.C(n_932),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1091),
.A2(n_974),
.B1(n_950),
.B2(n_1001),
.C(n_966),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1091),
.A2(n_952),
.B(n_970),
.C(n_956),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_1104),
.B(n_60),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1107),
.B(n_950),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1123),
.A2(n_1108),
.B(n_1119),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1115),
.Y(n_1133)
);

BUFx2_ASAP7_75t_R g1134 ( 
.A(n_1116),
.Y(n_1134)
);

AOI311xp33_ASAP7_75t_L g1135 ( 
.A1(n_1126),
.A2(n_911),
.A3(n_903),
.B(n_906),
.C(n_916),
.Y(n_1135)
);

NOR2x1_ASAP7_75t_L g1136 ( 
.A(n_1114),
.B(n_883),
.Y(n_1136)
);

OAI211xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1110),
.A2(n_63),
.B(n_68),
.C(n_70),
.Y(n_1137)
);

OAI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1124),
.A2(n_952),
.B1(n_958),
.B2(n_883),
.C(n_943),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_SL g1139 ( 
.A(n_1131),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1113),
.Y(n_1140)
);

AO21x1_ASAP7_75t_L g1141 ( 
.A1(n_1112),
.A2(n_947),
.B(n_976),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1121),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1109),
.A2(n_958),
.B1(n_947),
.B2(n_952),
.Y(n_1143)
);

NAND2x1_ASAP7_75t_SL g1144 ( 
.A(n_1117),
.B(n_952),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1130),
.B(n_988),
.Y(n_1145)
);

OAI221xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1129),
.A2(n_1127),
.B1(n_1118),
.B2(n_1128),
.C(n_1125),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1111),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1122),
.B(n_952),
.C(n_883),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1120),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1119),
.Y(n_1150)
);

AOI222xp33_ASAP7_75t_L g1151 ( 
.A1(n_1127),
.A2(n_989),
.B1(n_1000),
.B2(n_973),
.C1(n_975),
.C2(n_969),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1110),
.B(n_989),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1123),
.A2(n_966),
.B1(n_1000),
.B2(n_991),
.C(n_990),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1123),
.A2(n_966),
.B1(n_1000),
.B2(n_991),
.C(n_990),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_1119),
.B(n_73),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_L g1156 ( 
.A(n_1150),
.B(n_74),
.Y(n_1156)
);

XNOR2x1_ASAP7_75t_L g1157 ( 
.A(n_1140),
.B(n_75),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1152),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1133),
.B(n_990),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_L g1160 ( 
.A(n_1132),
.B(n_973),
.C(n_975),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1137),
.B(n_78),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1138),
.B(n_79),
.C(n_83),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1139),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1136),
.Y(n_1164)
);

NAND4xp75_ASAP7_75t_L g1165 ( 
.A(n_1142),
.B(n_956),
.C(n_991),
.D(n_995),
.Y(n_1165)
);

NAND4xp75_ASAP7_75t_L g1166 ( 
.A(n_1141),
.B(n_956),
.C(n_995),
.D(n_937),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1155),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1147),
.B(n_995),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1134),
.B(n_85),
.Y(n_1169)
);

OAI211xp5_ASAP7_75t_L g1170 ( 
.A1(n_1144),
.A2(n_956),
.B(n_969),
.C(n_937),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1147),
.B(n_947),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1145),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1147),
.Y(n_1173)
);

AO22x2_ASAP7_75t_L g1174 ( 
.A1(n_1149),
.A2(n_1148),
.B1(n_1143),
.B2(n_1146),
.Y(n_1174)
);

NAND4xp25_ASAP7_75t_L g1175 ( 
.A(n_1135),
.B(n_938),
.C(n_955),
.D(n_947),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1154),
.B(n_938),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1153),
.B(n_88),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1163),
.B(n_1151),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1173),
.A2(n_958),
.B1(n_943),
.B2(n_976),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1169),
.B(n_956),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1164),
.A2(n_976),
.B(n_924),
.Y(n_1181)
);

NOR2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1158),
.B(n_89),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1167),
.B(n_90),
.C(n_93),
.Y(n_1183)
);

OAI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1162),
.A2(n_958),
.B1(n_943),
.B2(n_924),
.C(n_929),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1174),
.A2(n_976),
.B1(n_929),
.B2(n_955),
.C(n_927),
.Y(n_1185)
);

XOR2xp5_ASAP7_75t_L g1186 ( 
.A(n_1157),
.B(n_94),
.Y(n_1186)
);

NOR3xp33_ASAP7_75t_L g1187 ( 
.A(n_1172),
.B(n_95),
.C(n_96),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_1156),
.B(n_1171),
.C(n_1168),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1174),
.A2(n_929),
.B(n_890),
.Y(n_1189)
);

AND3x4_ASAP7_75t_L g1190 ( 
.A(n_1161),
.B(n_968),
.C(n_106),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1159),
.A2(n_913),
.B1(n_925),
.B2(n_927),
.C(n_968),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_SL g1192 ( 
.A(n_1177),
.B(n_949),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1188),
.B(n_1159),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1192),
.A2(n_1160),
.B1(n_1176),
.B2(n_1170),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1182),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1178),
.A2(n_1166),
.B(n_1165),
.C(n_1175),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1189),
.B(n_105),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1186),
.B(n_949),
.Y(n_1198)
);

AOI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1181),
.A2(n_1190),
.B1(n_1183),
.B2(n_1185),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1184),
.A2(n_951),
.B1(n_915),
.B2(n_114),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1180),
.Y(n_1201)
);

AO21x1_ASAP7_75t_L g1202 ( 
.A1(n_1187),
.A2(n_110),
.B(n_111),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1179),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1191),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1188),
.A2(n_913),
.B1(n_927),
.B2(n_925),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1190),
.Y(n_1206)
);

AOI21xp33_ASAP7_75t_L g1207 ( 
.A1(n_1178),
.A2(n_115),
.B(n_118),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1195),
.A2(n_951),
.B1(n_915),
.B2(n_124),
.Y(n_1208)
);

OAI22x1_ASAP7_75t_L g1209 ( 
.A1(n_1199),
.A2(n_927),
.B1(n_925),
.B2(n_913),
.Y(n_1209)
);

AO22x2_ASAP7_75t_L g1210 ( 
.A1(n_1193),
.A2(n_913),
.B1(n_925),
.B2(n_916),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1197),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1206),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1193),
.A2(n_1194),
.B1(n_1203),
.B2(n_1200),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1201),
.A2(n_914),
.B1(n_911),
.B2(n_908),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1204),
.A2(n_951),
.B1(n_949),
.B2(n_125),
.Y(n_1215)
);

OAI22x1_ASAP7_75t_L g1216 ( 
.A1(n_1198),
.A2(n_951),
.B1(n_122),
.B2(n_127),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1202),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1217),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1211),
.B(n_1196),
.Y(n_1219)
);

AOI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1212),
.A2(n_1207),
.B1(n_1205),
.B2(n_132),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1213),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1216),
.Y(n_1222)
);

NOR3xp33_ASAP7_75t_L g1223 ( 
.A(n_1208),
.B(n_1209),
.C(n_1215),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1221),
.B(n_120),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1218),
.Y(n_1225)
);

BUFx4f_ASAP7_75t_SL g1226 ( 
.A(n_1222),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1223),
.B(n_1210),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1225),
.A2(n_1219),
.B(n_1220),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_1226),
.B1(n_1227),
.B2(n_1214),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1229),
.B(n_1224),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1230),
.A2(n_908),
.B1(n_899),
.B2(n_914),
.Y(n_1231)
);

OAI221xp5_ASAP7_75t_R g1232 ( 
.A1(n_1231),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.C(n_138),
.Y(n_1232)
);

AOI211xp5_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_142),
.B(n_143),
.C(n_145),
.Y(n_1233)
);


endmodule