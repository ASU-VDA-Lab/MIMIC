module fake_jpeg_20397_n_18 (n_0, n_3, n_2, n_1, n_18);

input n_0;
input n_3;
input n_2;
input n_1;

output n_18;

wire n_13;
wire n_11;
wire n_14;
wire n_17;
wire n_16;
wire n_10;
wire n_12;
wire n_4;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

INVx5_ASAP7_75t_L g4 ( 
.A(n_2),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_3),
.Y(n_5)
);

INVx6_ASAP7_75t_SL g6 ( 
.A(n_2),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_SL g8 ( 
.A1(n_5),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_8)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_6),
.B(n_1),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_0),
.C(n_1),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_4),
.C(n_5),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_7),
.B(n_6),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_13),
.Y(n_15)
);

AOI321xp33_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_7),
.A3(n_6),
.B1(n_0),
.B2(n_9),
.C(n_4),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_6),
.B(n_4),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_16),
.A2(n_15),
.B(n_7),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_7),
.C(n_0),
.Y(n_18)
);


endmodule