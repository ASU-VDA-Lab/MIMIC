module fake_jpeg_14954_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_40),
.B(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_23),
.B(n_3),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_16),
.B(n_30),
.C(n_29),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_24),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_37),
.C(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_53),
.C(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_28),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_56),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_32),
.B1(n_38),
.B2(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_33),
.B1(n_53),
.B2(n_5),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_32),
.B1(n_38),
.B2(n_28),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_55),
.B1(n_51),
.B2(n_57),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_17),
.B1(n_22),
.B2(n_21),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_57),
.A3(n_45),
.B1(n_37),
.B2(n_54),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_94),
.B(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_91),
.B1(n_65),
.B2(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_101),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_44),
.C(n_46),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_99),
.C(n_64),
.Y(n_107)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_100),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_33),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_79),
.B(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_33),
.B1(n_59),
.B2(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_18),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_77),
.C(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_122),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_115),
.B1(n_123),
.B2(n_109),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_83),
.B(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_67),
.B(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_63),
.Y(n_128)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_63),
.B1(n_65),
.B2(n_5),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_2),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_123),
.B1(n_112),
.B2(n_111),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_135),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_83),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_115),
.C(n_91),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_90),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_160),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_110),
.A3(n_114),
.B1(n_118),
.B2(n_104),
.C1(n_108),
.C2(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_141),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_132),
.C(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_159),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_118),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_96),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_84),
.B1(n_104),
.B2(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_97),
.C(n_94),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_88),
.B1(n_94),
.B2(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_153),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_172),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_142),
.B(n_138),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_148),
.B(n_147),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.C(n_173),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_132),
.C(n_127),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_174),
.B(n_98),
.Y(n_185)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_137),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_181),
.B1(n_164),
.B2(n_170),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_160),
.B1(n_145),
.B2(n_158),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_185),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_157),
.B1(n_144),
.B2(n_127),
.Y(n_181)
);

FAx1_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_159),
.CI(n_134),
.CON(n_183),
.SN(n_183)
);

OAI21x1_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_177),
.B(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_154),
.C(n_63),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_182),
.C(n_179),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_193),
.C(n_191),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_13),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_6),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_182),
.C(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_199),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_183),
.B(n_12),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_3),
.B(n_5),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_3),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_200),
.B(n_6),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_8),
.B(n_9),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_11),
.Y(n_205)
);

AOI21x1_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_198),
.B(n_8),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_9),
.B(n_10),
.Y(n_213)
);

OA21x2_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_207),
.B(n_208),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_10),
.B(n_212),
.Y(n_215)
);


endmodule