module fake_jpeg_19139_n_180 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_5),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_32)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_11),
.B1(n_14),
.B2(n_17),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_26),
.B1(n_28),
.B2(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_33),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_49),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_48),
.B1(n_39),
.B2(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_22),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_27),
.C(n_31),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_55),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_58),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_36),
.B(n_37),
.C(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_52),
.B1(n_51),
.B2(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_64),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_27),
.C(n_34),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_39),
.B1(n_13),
.B2(n_12),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_77),
.B(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_40),
.B1(n_45),
.B2(n_49),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_41),
.B(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_81),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2x1_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_55),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_86),
.B(n_72),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_93),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_61),
.C(n_60),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.C(n_71),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_63),
.C(n_54),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_59),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_74),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_57),
.B(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_102),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_74),
.B1(n_64),
.B2(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_91),
.B1(n_89),
.B2(n_85),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_86),
.B(n_85),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_95),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_45),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_49),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_40),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_16),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_40),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_110),
.B1(n_113),
.B2(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_120),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_18),
.B(n_9),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_129),
.C(n_102),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_18),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_21),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_101),
.B1(n_99),
.B2(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_136),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_139),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_117),
.C(n_121),
.Y(n_147)
);

AOI31xp67_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_104),
.A3(n_16),
.B(n_21),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_16),
.B1(n_7),
.B2(n_10),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_116),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_150),
.Y(n_160)
);

XOR2x1_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_120),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_117),
.C(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_18),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_116),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_161),
.C(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_146),
.B(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_137),
.B1(n_127),
.B2(n_129),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_160),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_6),
.B1(n_10),
.B2(n_9),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_5),
.C(n_9),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_3),
.C(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_10),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_3),
.B1(n_4),
.B2(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.C(n_4),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_168),
.B(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_178),
.Y(n_180)
);


endmodule