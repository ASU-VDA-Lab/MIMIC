module fake_jpeg_30967_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_5),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_32),
.Y(n_47)
);

CKINVDCx9p33_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_12),
.B1(n_19),
.B2(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_53),
.B1(n_57),
.B2(n_37),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_19),
.B(n_12),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_43),
.B(n_47),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_30),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_22),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_23),
.B1(n_16),
.B2(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_42),
.B1(n_40),
.B2(n_31),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_77),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_73),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_14),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_14),
.B1(n_22),
.B2(n_13),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_13),
.B1(n_8),
.B2(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_62),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_8),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_81),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_65),
.B(n_44),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_67),
.B1(n_94),
.B2(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_83),
.B1(n_96),
.B2(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_107),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_68),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_84),
.C(n_95),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_67),
.B(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_77),
.B1(n_63),
.B2(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_98),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_85),
.A3(n_88),
.B1(n_83),
.B2(n_80),
.C1(n_69),
.C2(n_89),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_85),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_114),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_91),
.B(n_87),
.C(n_86),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_105),
.B1(n_100),
.B2(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.C(n_119),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_100),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_105),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_125),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_113),
.B1(n_97),
.B2(n_93),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_113),
.B1(n_76),
.B2(n_45),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_120),
.B(n_59),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_127),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_58),
.C(n_61),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_69),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_133),
.B(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_129),
.C(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_60),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_62),
.Y(n_136)
);


endmodule