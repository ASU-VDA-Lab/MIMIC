module fake_jpeg_1750_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_73),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_58),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_1),
.B(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_62),
.C(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_71),
.Y(n_105)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_57),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_90),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_103),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_76),
.B1(n_58),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_65),
.B1(n_53),
.B2(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_60),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_83),
.C(n_45),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_87),
.B1(n_63),
.B2(n_54),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_113),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_119),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_59),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_87),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_126),
.Y(n_128)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_49),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_29),
.B(n_26),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_104),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_136),
.C(n_140),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_100),
.B(n_108),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_131),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_1),
.B(n_2),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_147),
.B1(n_5),
.B2(n_8),
.C(n_9),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_137),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_43),
.C(n_39),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_36),
.C(n_35),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_32),
.C(n_30),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_145),
.C(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_24),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_3),
.CI(n_4),
.CON(n_147),
.SN(n_147)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_16),
.C(n_6),
.D(n_7),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_161),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

OR2x4_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_10),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_145),
.Y(n_171)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_130),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.C(n_162),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_163),
.B(n_154),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_132),
.B1(n_148),
.B2(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_172),
.A2(n_174),
.B1(n_150),
.B2(n_156),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_162),
.B(n_157),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_179),
.B1(n_173),
.B2(n_12),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_152),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_156),
.A3(n_164),
.B1(n_154),
.B2(n_141),
.C1(n_15),
.C2(n_11),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.C(n_178),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_11),
.B(n_12),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.C(n_183),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_181),
.C(n_14),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_13),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_15),
.Y(n_190)
);


endmodule