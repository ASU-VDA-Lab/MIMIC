module fake_jpeg_23808_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_31),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_26),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_53),
.Y(n_59)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_21),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_26),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_25),
.B(n_16),
.Y(n_86)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_40),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_37),
.C(n_41),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_53),
.C(n_56),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_71),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_86),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_41),
.B1(n_43),
.B2(n_50),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_41),
.B1(n_38),
.B2(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_32),
.B1(n_17),
.B2(n_27),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_77),
.B1(n_16),
.B2(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_38),
.B1(n_26),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_33),
.B1(n_25),
.B2(n_20),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_36),
.B(n_39),
.C(n_22),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_24),
.B(n_28),
.C(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_99),
.B1(n_111),
.B2(n_78),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_106),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_103),
.B(n_66),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_53),
.C(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_108),
.B1(n_88),
.B2(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_58),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_63),
.B(n_29),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_63),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_33),
.B1(n_20),
.B2(n_23),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_119),
.B1(n_97),
.B2(n_95),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_80),
.B1(n_76),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_133),
.B1(n_103),
.B2(n_97),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_120),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_125),
.B(n_136),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_126),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_70),
.B(n_75),
.C(n_65),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_131),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_70),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_68),
.B1(n_85),
.B2(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_155),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_97),
.CI(n_106),
.CON(n_151),
.SN(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_115),
.C(n_60),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_96),
.B1(n_93),
.B2(n_100),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_153),
.A2(n_121),
.B1(n_79),
.B2(n_24),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_157),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_92),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_93),
.B(n_62),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_144),
.B(n_154),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_167),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_115),
.B(n_132),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_168),
.B(n_149),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_177),
.B(n_139),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_124),
.C(n_114),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_174),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_153),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_120),
.B(n_117),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_62),
.C(n_60),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_172),
.C(n_1),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_67),
.C(n_81),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_0),
.B(n_1),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_176),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_158),
.B(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_121),
.B1(n_138),
.B2(n_137),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_187),
.B(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_192),
.C(n_166),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_147),
.C(n_151),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_184),
.C(n_162),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_147),
.C(n_151),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_157),
.A3(n_141),
.B1(n_149),
.B2(n_146),
.C(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_137),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_0),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_195),
.Y(n_206)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_194),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_199),
.C(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_172),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_161),
.C(n_175),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_180),
.B(n_177),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_209),
.B(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_205),
.C(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_164),
.B1(n_184),
.B2(n_160),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_167),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_164),
.B1(n_170),
.B2(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_209),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_191),
.B1(n_168),
.B2(n_178),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_15),
.A3(n_13),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.C(n_217),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_201),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_6),
.C2(n_7),
.Y(n_215)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_2),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_201),
.Y(n_217)
);

AOI31xp33_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_219),
.A3(n_7),
.B(n_8),
.Y(n_223)
);

NAND2xp67_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_2),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_208),
.B(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_10),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_205),
.C(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_8),
.C(n_10),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_224),
.C(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_229),
.Y(n_232)
);


endmodule