module fake_jpeg_8210_n_47 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_47);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_20),
.B1(n_8),
.B2(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_0),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_6),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

AOI31xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_43),
.A3(n_16),
.B(n_36),
.Y(n_47)
);


endmodule