module fake_jpeg_21731_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_21),
.Y(n_28)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_18),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_11),
.B1(n_10),
.B2(n_12),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_12),
.B(n_19),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_11),
.B1(n_10),
.B2(n_17),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_29),
.B1(n_21),
.B2(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_21),
.C(n_20),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_9),
.B(n_13),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_37),
.B1(n_31),
.B2(n_39),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_46),
.B1(n_48),
.B2(n_22),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_28),
.B1(n_10),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_10),
.B1(n_24),
.B2(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_48),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_56),
.B(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_22),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.C(n_58),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_24),
.C(n_18),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_14),
.B1(n_24),
.B2(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_13),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_66),
.B(n_70),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_45),
.C(n_46),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_15),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_15),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_27),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_0),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_79),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_55),
.B(n_56),
.C(n_15),
.D(n_14),
.Y(n_74)
);

OA21x2_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_81),
.B(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_78),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_80),
.Y(n_87)
);

AOI322xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_61),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_88),
.C(n_83),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_13),
.C(n_9),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_95),
.B1(n_88),
.B2(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_72),
.C(n_75),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_82),
.B(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI221xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_87),
.B(n_79),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_90),
.B(n_85),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_5),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_96),
.C(n_2),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

OAI221xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_104)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_8),
.B(n_0),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_109),
.B(n_106),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_1),
.Y(n_111)
);


endmodule