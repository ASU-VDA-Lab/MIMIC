module real_jpeg_28917_n_10 (n_8, n_57, n_0, n_54, n_2, n_55, n_58, n_52, n_9, n_6, n_60, n_59, n_7, n_53, n_3, n_5, n_4, n_1, n_56, n_10);

input n_8;
input n_57;
input n_0;
input n_54;
input n_2;
input n_55;
input n_58;
input n_52;
input n_9;
input n_6;
input n_60;
input n_59;
input n_7;
input n_53;
input n_3;
input n_5;
input n_4;
input n_1;
input n_56;

output n_10;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_49;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_20),
.C(n_37),
.Y(n_19)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_18),
.C(n_43),
.Y(n_17)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_12),
.Y(n_11)
);

FAx1_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_22),
.CI(n_25),
.CON(n_21),
.SN(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_16),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_46),
.C(n_47),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.C(n_40),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.C(n_34),
.Y(n_20)
);

BUFx24_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.C(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_52),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_53),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_54),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_55),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_56),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_57),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_58),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_59),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_60),
.Y(n_49)
);


endmodule