module fake_jpeg_11530_n_429 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_50),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_67),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_16),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_83),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_12),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_40),
.B(n_15),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_27),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_27),
.Y(n_93)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_93),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_27),
.B1(n_36),
.B2(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_97),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_39),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_27),
.B1(n_20),
.B2(n_38),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_20),
.B1(n_38),
.B2(n_43),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_38),
.B1(n_20),
.B2(n_39),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_48),
.B(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_48),
.B(n_39),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_35),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_138),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_35),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_140),
.C(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_34),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_26),
.B1(n_75),
.B2(n_41),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_151),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_33),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_21),
.B1(n_52),
.B2(n_44),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_172),
.B1(n_109),
.B2(n_89),
.Y(n_186)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_164),
.Y(n_189)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_111),
.A2(n_94),
.B1(n_112),
.B2(n_78),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_54),
.B1(n_62),
.B2(n_50),
.Y(n_200)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_169),
.A2(n_132),
.B1(n_98),
.B2(n_125),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_89),
.A2(n_21),
.B1(n_47),
.B2(n_55),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_93),
.B(n_132),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_141),
.B(n_154),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_165),
.B1(n_155),
.B2(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_186),
.B1(n_193),
.B2(n_125),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_139),
.A2(n_64),
.B1(n_58),
.B2(n_63),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_98),
.B1(n_95),
.B2(n_21),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_149),
.Y(n_212)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_135),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_212),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_147),
.B(n_150),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_208),
.B(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_156),
.B1(n_142),
.B2(n_164),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_175),
.B(n_146),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_179),
.C(n_198),
.Y(n_229)
);

NAND2xp33_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_26),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_223),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_194),
.B(n_184),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_177),
.B(n_195),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_200),
.B1(n_183),
.B2(n_194),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_157),
.B1(n_174),
.B2(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_183),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_109),
.B1(n_114),
.B2(n_92),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_151),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_137),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_92),
.B1(n_144),
.B2(n_162),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_179),
.B1(n_173),
.B2(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_177),
.B1(n_148),
.B2(n_169),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_229),
.B(n_207),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_202),
.B1(n_219),
.B2(n_228),
.Y(n_263)
);

BUFx4f_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_195),
.B1(n_192),
.B2(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_104),
.B1(n_49),
.B2(n_56),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_195),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_237),
.B(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_196),
.C(n_173),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_249),
.C(n_254),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_250),
.B1(n_252),
.B2(n_209),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_208),
.B(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_190),
.C(n_129),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_197),
.B1(n_192),
.B2(n_199),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_26),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_192),
.B1(n_199),
.B2(n_145),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_118),
.C(n_171),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_136),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_255),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_266),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_211),
.B1(n_221),
.B2(n_214),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_264),
.B1(n_267),
.B2(n_271),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_262),
.A2(n_284),
.B(n_238),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_214),
.B1(n_212),
.B2(n_203),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_204),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_273),
.C(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_230),
.A2(n_205),
.B1(n_224),
.B2(n_204),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_209),
.B1(n_204),
.B2(n_216),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_268),
.A2(n_280),
.B1(n_283),
.B2(n_232),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_234),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.Y(n_290)
);

AO22x1_ASAP7_75t_SL g270 ( 
.A1(n_230),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_117),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_277),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_41),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_276),
.B(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_239),
.B1(n_251),
.B2(n_253),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_231),
.A2(n_51),
.B1(n_87),
.B2(n_103),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_238),
.A2(n_98),
.B(n_33),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_281),
.A2(n_242),
.B(n_245),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_72),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_231),
.A2(n_95),
.B1(n_72),
.B2(n_82),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_41),
.B(n_34),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_251),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_233),
.B(n_12),
.Y(n_286)
);

XNOR2x2_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_289),
.A2(n_23),
.B(n_22),
.Y(n_335)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_291),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_262),
.A2(n_249),
.B1(n_229),
.B2(n_233),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_295),
.A2(n_23),
.B(n_22),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_302),
.B1(n_309),
.B2(n_279),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_253),
.B1(n_254),
.B2(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_300),
.B(n_306),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_246),
.C(n_235),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_308),
.C(n_284),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_269),
.A2(n_235),
.B1(n_34),
.B2(n_33),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_235),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_258),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_272),
.B(n_32),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_264),
.B(n_32),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_32),
.C(n_31),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_281),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_257),
.B(n_31),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_329),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_318),
.Y(n_343)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_256),
.B1(n_270),
.B2(n_267),
.Y(n_322)
);

NAND2x1p5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_332),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_285),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_330),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_327),
.C(n_331),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_261),
.C(n_274),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_312),
.A2(n_256),
.B1(n_260),
.B2(n_277),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_283),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_278),
.C(n_280),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_288),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_336),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_304),
.C(n_298),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_305),
.C(n_308),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_289),
.B(n_296),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_0),
.B(n_1),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_288),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_337),
.B(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_316),
.B(n_310),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_349),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_305),
.B1(n_297),
.B2(n_290),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_342),
.A2(n_344),
.B1(n_348),
.B2(n_357),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_328),
.A2(n_290),
.B1(n_305),
.B2(n_292),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_347),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_311),
.B1(n_310),
.B2(n_302),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_311),
.C(n_309),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_314),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_350),
.A2(n_335),
.B1(n_336),
.B2(n_315),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_0),
.C(n_1),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_317),
.C(n_326),
.Y(n_367)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_321),
.B(n_1),
.Y(n_356)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_323),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_357)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_318),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_363),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_343),
.B(n_315),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_354),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_373),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_367),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_338),
.A2(n_323),
.B1(n_331),
.B2(n_334),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_368),
.A2(n_346),
.B1(n_349),
.B2(n_355),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_344),
.A2(n_329),
.B1(n_322),
.B2(n_330),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_372),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_343),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_322),
.C(n_332),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_322),
.C(n_3),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_2),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_380),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_354),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_386),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_375),
.B(n_348),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_382),
.B(n_385),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_362),
.B(n_357),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_352),
.B(n_351),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_359),
.A2(n_339),
.B(n_351),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_373),
.B(n_351),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_SL g401 ( 
.A(n_388),
.B(n_4),
.C(n_5),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_363),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_372),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_390),
.B(n_393),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_371),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_395),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_376),
.A2(n_388),
.B1(n_378),
.B2(n_374),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_386),
.B1(n_5),
.B2(n_6),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_370),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_389),
.B(n_367),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_396),
.B(n_6),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_353),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_398),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_2),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_4),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_381),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_404),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_11),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_405),
.B(n_410),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_411),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_400),
.A2(n_5),
.B(n_6),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_408),
.A2(n_400),
.B(n_401),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_6),
.Y(n_411)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_414),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_7),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_415),
.B(n_416),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_7),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_403),
.A2(n_7),
.B(n_9),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_417),
.A2(n_9),
.B(n_10),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_412),
.B(n_405),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_420),
.B(n_422),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_414),
.A2(n_404),
.B(n_10),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_418),
.C(n_413),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_424),
.A2(n_421),
.B(n_419),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_425),
.C(n_10),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_427),
.B(n_11),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_11),
.Y(n_429)
);


endmodule