module real_aes_6822_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_1), .A2(n_135), .B(n_139), .C(n_220), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_2), .A2(n_169), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g513 ( .A(n_3), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_4), .B(n_236), .Y(n_255) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_169), .B(n_479), .Y(n_478) );
AND2x6_ASAP7_75t_L g135 ( .A(n_6), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g210 ( .A(n_7), .Y(n_210) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_8), .B(n_41), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_9), .A2(n_168), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_10), .B(n_147), .Y(n_222) );
INVx1_ASAP7_75t_L g483 ( .A(n_11), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_12), .B(n_250), .Y(n_538) );
INVx1_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
INVx1_ASAP7_75t_L g550 ( .A(n_14), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_15), .A2(n_145), .B(n_232), .C(n_234), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_16), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_17), .B(n_501), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_18), .B(n_169), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_19), .B(n_181), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_20), .A2(n_250), .B(n_265), .C(n_267), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_21), .B(n_236), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_22), .B(n_147), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_23), .A2(n_177), .B(n_234), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_24), .B(n_147), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_25), .Y(n_186) );
INVx1_ASAP7_75t_L g143 ( .A(n_26), .Y(n_143) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_27), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_28), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_29), .B(n_147), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_30), .A2(n_31), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_30), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_31), .Y(n_748) );
INVx1_ASAP7_75t_L g175 ( .A(n_32), .Y(n_175) );
INVx1_ASAP7_75t_L g492 ( .A(n_33), .Y(n_492) );
INVx2_ASAP7_75t_L g133 ( .A(n_34), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_35), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_36), .A2(n_250), .B(n_251), .C(n_253), .Y(n_249) );
INVxp67_ASAP7_75t_L g176 ( .A(n_37), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_38), .A2(n_139), .B(n_142), .C(n_150), .Y(n_138) );
CKINVDCx14_ASAP7_75t_R g248 ( .A(n_39), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_40), .A2(n_135), .B(n_139), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g491 ( .A(n_42), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_43), .A2(n_194), .B(n_208), .C(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_44), .B(n_147), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_45), .A2(n_746), .B1(n_747), .B2(n_750), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_45), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_46), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_47), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_48), .A2(n_104), .B1(n_113), .B2(n_759), .Y(n_103) );
INVx1_ASAP7_75t_L g263 ( .A(n_49), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_50), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_51), .B(n_169), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_52), .B(n_458), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_53), .A2(n_139), .B1(n_267), .B2(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_54), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_55), .Y(n_510) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_56), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_57), .A2(n_208), .B(n_253), .C(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_58), .Y(n_566) );
INVx1_ASAP7_75t_L g480 ( .A(n_59), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_60), .A2(n_89), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_60), .Y(n_450) );
INVx1_ASAP7_75t_L g136 ( .A(n_61), .Y(n_136) );
INVx1_ASAP7_75t_L g154 ( .A(n_62), .Y(n_154) );
INVx1_ASAP7_75t_SL g252 ( .A(n_63), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_65), .B(n_236), .Y(n_269) );
INVx1_ASAP7_75t_L g189 ( .A(n_66), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_67), .A2(n_253), .B(n_501), .C(n_502), .Y(n_500) );
INVxp67_ASAP7_75t_L g503 ( .A(n_68), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_69), .A2(n_120), .B1(n_121), .B2(n_122), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_69), .Y(n_120) );
INVx1_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_71), .A2(n_169), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_72), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_73), .A2(n_169), .B(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_74), .Y(n_495) );
INVx1_ASAP7_75t_L g560 ( .A(n_75), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_76), .A2(n_168), .B(n_170), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g137 ( .A(n_77), .Y(n_137) );
INVx1_ASAP7_75t_L g230 ( .A(n_78), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_79), .A2(n_135), .B(n_139), .C(n_562), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_80), .A2(n_169), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g233 ( .A(n_81), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_82), .B(n_144), .Y(n_526) );
INVx2_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g221 ( .A(n_84), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_85), .B(n_501), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_86), .A2(n_135), .B(n_139), .C(n_512), .Y(n_511) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_87), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g453 ( .A(n_87), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g465 ( .A(n_87), .B(n_455), .Y(n_465) );
INVx2_ASAP7_75t_L g469 ( .A(n_87), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_88), .A2(n_139), .B(n_188), .C(n_196), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_89), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_90), .B(n_151), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_91), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_92), .A2(n_135), .B(n_139), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_93), .Y(n_542) );
INVx1_ASAP7_75t_L g499 ( .A(n_94), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_95), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_96), .B(n_144), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_97), .B(n_159), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_98), .B(n_159), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g266 ( .A(n_100), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_101), .A2(n_169), .B(n_498), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_102), .A2(n_462), .B1(n_744), .B2(n_745), .C1(n_751), .C2(n_754), .Y(n_461) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g455 ( .A(n_109), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_460), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g758 ( .A(n_116), .Y(n_758) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_451), .B(n_457), .Y(n_118) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_448), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_123), .A2(n_463), .B1(n_466), .B2(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g752 ( .A(n_123), .Y(n_752) );
OR4x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_338), .C(n_385), .D(n_425), .Y(n_123) );
NAND3xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_284), .C(n_313), .Y(n_124) );
AOI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_199), .B(n_237), .C(n_277), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_126), .A2(n_297), .B(n_314), .C(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_161), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_128), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_SL g280 ( .A(n_128), .Y(n_280) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_128), .Y(n_292) );
AND2x4_ASAP7_75t_L g296 ( .A(n_128), .B(n_244), .Y(n_296) );
AND2x2_ASAP7_75t_L g307 ( .A(n_128), .B(n_184), .Y(n_307) );
OR2x2_ASAP7_75t_L g331 ( .A(n_128), .B(n_240), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_128), .B(n_245), .Y(n_344) );
AND2x2_ASAP7_75t_L g384 ( .A(n_128), .B(n_370), .Y(n_384) );
AND2x2_ASAP7_75t_L g391 ( .A(n_128), .B(n_354), .Y(n_391) );
AND2x2_ASAP7_75t_L g421 ( .A(n_128), .B(n_162), .Y(n_421) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_156), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_138), .C(n_151), .Y(n_129) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_130), .A2(n_186), .B(n_187), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_130), .A2(n_218), .B(n_219), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_130), .A2(n_179), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_130), .A2(n_510), .B(n_511), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_130), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
AND2x4_ASAP7_75t_L g169 ( .A(n_131), .B(n_135), .Y(n_169) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g149 ( .A(n_132), .Y(n_149) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g140 ( .A(n_133), .Y(n_140) );
INVx1_ASAP7_75t_L g268 ( .A(n_133), .Y(n_268) );
INVx1_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx3_ASAP7_75t_L g145 ( .A(n_134), .Y(n_145) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx1_ASAP7_75t_L g501 ( .A(n_134), .Y(n_501) );
BUFx3_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
INVx4_ASAP7_75t_SL g179 ( .A(n_135), .Y(n_179) );
INVx5_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g195 ( .A(n_140), .Y(n_195) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_140), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_146), .C(n_148), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_144), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_144), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_145), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_145), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_145), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
INVx4_ASAP7_75t_L g250 ( .A(n_147), .Y(n_250) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_149), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_151), .A2(n_204), .B(n_211), .Y(n_203) );
INVx1_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_151), .A2(n_545), .B(n_551), .Y(n_544) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_L g160 ( .A(n_152), .B(n_153), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_158), .A2(n_185), .B(n_197), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_158), .B(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
NOR2xp33_ASAP7_75t_SL g528 ( .A(n_158), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_159), .Y(n_227) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_159), .A2(n_497), .B(n_504), .Y(n_496) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_161), .B(n_348), .Y(n_360) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_183), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_162), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g298 ( .A(n_162), .B(n_183), .Y(n_298) );
BUFx3_ASAP7_75t_L g306 ( .A(n_162), .Y(n_306) );
OR2x2_ASAP7_75t_L g327 ( .A(n_162), .B(n_202), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_162), .B(n_348), .Y(n_438) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_180), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_164), .A2(n_241), .B(n_242), .Y(n_240) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_164), .A2(n_559), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_165), .A2(n_523), .B(n_524), .Y(n_522) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_166), .A2(n_488), .B(n_494), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_166), .B(n_495), .Y(n_494) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_166), .A2(n_509), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g241 ( .A(n_167), .Y(n_241) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_179), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g205 ( .A1(n_172), .A2(n_179), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g229 ( .A1(n_172), .A2(n_179), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_172), .A2(n_179), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_172), .A2(n_179), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_172), .A2(n_179), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_172), .A2(n_179), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_172), .A2(n_179), .B(n_547), .C(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_177), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_177), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_177), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g490 ( .A1(n_178), .A2(n_191), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g196 ( .A(n_179), .Y(n_196) );
INVx1_ASAP7_75t_L g242 ( .A(n_180), .Y(n_242) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_182), .B(n_198), .Y(n_197) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_182), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_L g243 ( .A(n_183), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g291 ( .A(n_183), .Y(n_291) );
AND2x2_ASAP7_75t_L g354 ( .A(n_183), .B(n_245), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_183), .A2(n_357), .B1(n_359), .B2(n_361), .C(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g370 ( .A(n_183), .B(n_240), .Y(n_370) );
AND2x2_ASAP7_75t_L g396 ( .A(n_183), .B(n_280), .Y(n_396) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g276 ( .A(n_184), .B(n_245), .Y(n_276) );
BUFx2_ASAP7_75t_L g410 ( .A(n_184), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_192), .C(n_193), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_190), .A2(n_193), .B(n_221), .C(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_193), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_193), .A2(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI32xp33_ASAP7_75t_L g376 ( .A1(n_200), .A2(n_337), .A3(n_351), .B1(n_377), .B2(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AND2x2_ASAP7_75t_L g317 ( .A(n_201), .B(n_259), .Y(n_317) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g299 ( .A(n_202), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_202), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g371 ( .A(n_202), .B(n_259), .Y(n_371) );
AND2x2_ASAP7_75t_L g382 ( .A(n_202), .B(n_274), .Y(n_382) );
BUFx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g283 ( .A(n_203), .B(n_260), .Y(n_283) );
AND2x2_ASAP7_75t_L g287 ( .A(n_203), .B(n_260), .Y(n_287) );
AND2x2_ASAP7_75t_L g322 ( .A(n_203), .B(n_273), .Y(n_322) );
AND2x2_ASAP7_75t_L g329 ( .A(n_203), .B(n_225), .Y(n_329) );
OAI211xp5_ASAP7_75t_L g334 ( .A1(n_203), .A2(n_280), .B(n_291), .C(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g388 ( .A(n_203), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_203), .B(n_214), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_212), .B(n_271), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_212), .B(n_287), .Y(n_377) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g282 ( .A(n_213), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_226), .Y(n_274) );
OR2x2_ASAP7_75t_L g289 ( .A(n_214), .B(n_226), .Y(n_289) );
AND2x2_ASAP7_75t_L g312 ( .A(n_214), .B(n_273), .Y(n_312) );
INVx1_ASAP7_75t_L g316 ( .A(n_214), .Y(n_316) );
AND2x2_ASAP7_75t_L g335 ( .A(n_214), .B(n_272), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_214), .A2(n_300), .B1(n_346), .B2(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_214), .B(n_388), .Y(n_412) );
AND2x2_ASAP7_75t_L g427 ( .A(n_214), .B(n_287), .Y(n_427) );
INVx4_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx3_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
AND2x2_ASAP7_75t_L g301 ( .A(n_215), .B(n_226), .Y(n_301) );
AND2x2_ASAP7_75t_L g303 ( .A(n_215), .B(n_259), .Y(n_303) );
AND3x2_ASAP7_75t_L g365 ( .A(n_215), .B(n_329), .C(n_366), .Y(n_365) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_216), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_216), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_216), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g400 ( .A(n_225), .B(n_272), .Y(n_400) );
INVx1_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g259 ( .A(n_226), .B(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_226), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_226), .B(n_271), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_226), .B(n_312), .C(n_388), .Y(n_440) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_235), .Y(n_226) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_227), .A2(n_246), .B(n_255), .Y(n_245) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_227), .A2(n_261), .B(n_269), .Y(n_260) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_236), .A2(n_478), .B(n_484), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_256), .B1(n_270), .B2(n_275), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_243), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_240), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g352 ( .A(n_240), .Y(n_352) );
OAI31xp33_ASAP7_75t_L g368 ( .A1(n_243), .A2(n_369), .A3(n_370), .B(n_371), .Y(n_368) );
AND2x2_ASAP7_75t_L g393 ( .A(n_243), .B(n_280), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_243), .B(n_306), .Y(n_439) );
AND2x2_ASAP7_75t_L g348 ( .A(n_244), .B(n_280), .Y(n_348) );
AND2x2_ASAP7_75t_L g409 ( .A(n_244), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g279 ( .A(n_245), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g337 ( .A(n_245), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_250), .B(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_254), .Y(n_539) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_257), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_258), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AOI221x1_ASAP7_75t_SL g325 ( .A1(n_259), .A2(n_326), .B1(n_328), .B2(n_330), .C(n_332), .Y(n_325) );
INVx2_ASAP7_75t_L g273 ( .A(n_260), .Y(n_273) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_260), .Y(n_367) );
INVx2_ASAP7_75t_L g515 ( .A(n_267), .Y(n_515) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g355 ( .A(n_270), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_271), .B(n_288), .Y(n_380) );
INVx1_ASAP7_75t_SL g443 ( .A(n_271), .Y(n_443) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g361 ( .A(n_274), .B(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g429 ( .A(n_275), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_275), .B(n_358), .Y(n_442) );
INVx2_ASAP7_75t_SL g281 ( .A(n_276), .Y(n_281) );
AND2x2_ASAP7_75t_L g324 ( .A(n_276), .B(n_280), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_276), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_276), .B(n_351), .Y(n_378) );
AOI21xp33_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_281), .B(n_282), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_279), .B(n_351), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_279), .B(n_306), .Y(n_447) );
OR2x2_ASAP7_75t_L g319 ( .A(n_280), .B(n_298), .Y(n_319) );
AND2x2_ASAP7_75t_L g418 ( .A(n_280), .B(n_409), .Y(n_418) );
OAI22xp5_ASAP7_75t_SL g293 ( .A1(n_281), .A2(n_294), .B1(n_299), .B2(n_302), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_281), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g341 ( .A(n_283), .B(n_289), .Y(n_341) );
INVx1_ASAP7_75t_L g405 ( .A(n_283), .Y(n_405) );
AOI311xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .A3(n_292), .B(n_293), .C(n_304), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_288), .A2(n_420), .B1(n_432), .B2(n_435), .C(n_437), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_288), .B(n_443), .Y(n_445) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g342 ( .A(n_290), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g332 ( .A1(n_291), .A2(n_333), .B(n_334), .C(n_336), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_SL g401 ( .A1(n_295), .A2(n_297), .B(n_402), .C(n_403), .Y(n_401) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_296), .B(n_370), .Y(n_436) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_299), .A2(n_319), .B1(n_320), .B2(n_323), .C(n_325), .Y(n_318) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g321 ( .A(n_301), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g404 ( .A(n_301), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_305), .A2(n_363), .B(n_364), .C(n_368), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_306), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_306), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g328 ( .A(n_312), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_316), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g430 ( .A(n_319), .Y(n_430) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_322), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g434 ( .A(n_322), .Y(n_434) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g375 ( .A(n_324), .B(n_351), .Y(n_375) );
INVx1_ASAP7_75t_SL g369 ( .A(n_331), .Y(n_369) );
INVx1_ASAP7_75t_L g346 ( .A(n_337), .Y(n_346) );
NAND3xp33_ASAP7_75t_SL g338 ( .A(n_339), .B(n_356), .C(n_372), .Y(n_338) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .A3(n_343), .B1(n_345), .B2(n_349), .C1(n_353), .C2(n_355), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_340), .A2(n_393), .B(n_394), .C(n_401), .Y(n_392) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_343), .A2(n_364), .B1(n_395), .B2(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_351), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g390 ( .A(n_351), .B(n_391), .Y(n_390) );
AOI32xp33_ASAP7_75t_L g441 ( .A1(n_351), .A2(n_442), .A3(n_443), .B1(n_444), .B2(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g363 ( .A(n_354), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_354), .A2(n_407), .B1(n_411), .B2(n_413), .C(n_416), .Y(n_406) );
AND2x2_ASAP7_75t_L g420 ( .A(n_354), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g423 ( .A(n_358), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g433 ( .A(n_358), .B(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g424 ( .A(n_367), .B(n_388), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_376), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_389), .B(n_392), .C(n_406), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_400), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g415 ( .A(n_412), .Y(n_415) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B(n_422), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_428), .B(n_431), .C(n_441), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_454), .B(n_469), .Y(n_756) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g468 ( .A(n_455), .B(n_469), .Y(n_468) );
AOI21xp33_ASAP7_75t_L g460 ( .A1(n_457), .A2(n_461), .B(n_757), .Y(n_460) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_463), .A2(n_466), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g753 ( .A(n_471), .Y(n_753) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_666), .C(n_711), .Y(n_472) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_589), .C(n_630), .D(n_647), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_505), .B(n_519), .C(n_552), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_476), .B(n_506), .Y(n_505) );
NOR4xp25_ASAP7_75t_L g613 ( .A(n_476), .B(n_607), .C(n_614), .D(n_620), .Y(n_613) );
AND2x2_ASAP7_75t_L g686 ( .A(n_476), .B(n_575), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_476), .B(n_651), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_476), .B(n_700), .Y(n_714) );
AND2x2_ASAP7_75t_L g727 ( .A(n_476), .B(n_518), .Y(n_727) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g572 ( .A(n_477), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_477), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g629 ( .A(n_477), .B(n_486), .Y(n_629) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_477), .B(n_575), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_477), .B(n_486), .Y(n_644) );
AND2x2_ASAP7_75t_L g653 ( .A(n_477), .B(n_578), .Y(n_653) );
BUFx2_ASAP7_75t_L g676 ( .A(n_477), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_477), .B(n_496), .Y(n_680) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_496), .Y(n_485) );
AND2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_496), .Y(n_518) );
BUFx2_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_486), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_614) );
OR2x2_ASAP7_75t_L g636 ( .A(n_486), .B(n_508), .Y(n_636) );
AND2x2_ASAP7_75t_L g700 ( .A(n_486), .B(n_578), .Y(n_700) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g568 ( .A(n_487), .B(n_508), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_487), .B(n_496), .Y(n_575) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_487), .Y(n_617) );
OR2x2_ASAP7_75t_L g652 ( .A(n_487), .B(n_507), .Y(n_652) );
INVx1_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
INVx3_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
BUFx2_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
AND2x2_ASAP7_75t_L g637 ( .A(n_496), .B(n_572), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_505), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_580), .Y(n_584) );
INVx1_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
INVx1_ASAP7_75t_L g590 ( .A(n_518), .Y(n_590) );
NAND2x1_ASAP7_75t_SL g519 ( .A(n_520), .B(n_530), .Y(n_519) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_543), .Y(n_588) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_520), .Y(n_662) );
AND2x2_ASAP7_75t_L g689 ( .A(n_520), .B(n_609), .Y(n_689) );
AND2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_659), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_520), .B(n_555), .Y(n_724) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g556 ( .A(n_521), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g573 ( .A(n_521), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g594 ( .A(n_521), .Y(n_594) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_521), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g633 ( .A(n_521), .B(n_558), .Y(n_633) );
OR2x2_ASAP7_75t_L g671 ( .A(n_521), .B(n_626), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g683 ( .A1(n_521), .A2(n_684), .A3(n_687), .B1(n_688), .B2(n_689), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_521), .B(n_659), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_521), .B(n_619), .Y(n_734) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g645 ( .A(n_531), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_543), .Y(n_531) );
INVx1_ASAP7_75t_L g607 ( .A(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_532), .B(n_557), .Y(n_626) );
AND2x2_ASAP7_75t_L g659 ( .A(n_532), .B(n_635), .Y(n_659) );
AND2x2_ASAP7_75t_L g696 ( .A(n_532), .B(n_558), .Y(n_696) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g555 ( .A(n_533), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_533), .B(n_557), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g634 ( .A(n_533), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_L g610 ( .A(n_543), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_543), .B(n_557), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_543), .B(n_601), .Y(n_682) );
INVx1_ASAP7_75t_L g704 ( .A(n_543), .Y(n_704) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_557), .Y(n_574) );
AND2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g635 ( .A(n_544), .Y(n_635) );
AOI221x1_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_567), .B1(n_573), .B2(n_575), .C(n_576), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_553), .A2(n_640), .B1(n_707), .B2(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
AND2x2_ASAP7_75t_L g598 ( .A(n_554), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g693 ( .A(n_554), .B(n_573), .Y(n_693) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g649 ( .A(n_555), .B(n_574), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
AND2x2_ASAP7_75t_L g672 ( .A(n_556), .B(n_659), .Y(n_672) );
AND2x2_ASAP7_75t_L g739 ( .A(n_556), .B(n_634), .Y(n_739) );
INVx2_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_568), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g691 ( .A(n_568), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_569), .B(n_652), .Y(n_655) );
INVx3_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_570), .A2(n_691), .B(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2xp33_ASAP7_75t_SL g713 ( .A(n_573), .B(n_599), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_574), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g665 ( .A(n_574), .B(n_593), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_574), .B(n_600), .Y(n_742) );
AND2x2_ASAP7_75t_L g611 ( .A(n_575), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g678 ( .A(n_575), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B(n_585), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g639 ( .A(n_578), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_578), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g663 ( .A(n_579), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_579), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_582), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_582), .A2(n_621), .B(n_651), .C(n_653), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_582), .A2(n_669), .B1(n_672), .B2(n_673), .C(n_677), .Y(n_668) );
AND2x2_ASAP7_75t_L g664 ( .A(n_583), .B(n_617), .Y(n_664) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g624 ( .A(n_588), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_597), .C(n_622), .Y(n_589) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_590), .B(n_709), .C(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
OR2x2_ASAP7_75t_L g681 ( .A(n_592), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_602), .B1(n_605), .B2(n_611), .C(n_613), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_599), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g621 ( .A(n_604), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
OR2x2_ASAP7_75t_L g741 ( .A(n_604), .B(n_652), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVxp67_ASAP7_75t_L g715 ( .A(n_607), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_609), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g616 ( .A(n_610), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_612), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_612), .B(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_612), .B(n_679), .Y(n_718) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g732 ( .A(n_621), .B(n_652), .Y(n_732) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g710 ( .A(n_627), .Y(n_710) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI322xp33_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_636), .A3(n_637), .B1(n_638), .B2(n_641), .C1(n_643), .C2(n_645), .Y(n_630) );
OAI322xp33_ASAP7_75t_L g712 ( .A1(n_631), .A2(n_713), .A3(n_714), .B1(n_715), .B2(n_716), .C1(n_717), .C2(n_719), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx4_ASAP7_75t_L g646 ( .A(n_633), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_633), .B(n_659), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_633), .B(n_721), .Y(n_720) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_636), .Y(n_731) );
INVx1_ASAP7_75t_L g709 ( .A(n_637), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OR2x2_ASAP7_75t_L g643 ( .A(n_639), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g726 ( .A(n_639), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_639), .B(n_680), .Y(n_737) );
OR2x2_ASAP7_75t_L g670 ( .A(n_642), .B(n_671), .Y(n_670) );
INVxp33_ASAP7_75t_L g687 ( .A(n_642), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_654), .C(n_656), .Y(n_647) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_646), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g730 ( .A(n_646), .Y(n_730) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_678), .A3(n_695), .B1(n_697), .B2(n_698), .C1(n_701), .C2(n_705), .Y(n_694) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_690), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_683), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_671), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
NAND2xp33_ASAP7_75t_SL g688 ( .A(n_674), .B(n_685), .Y(n_688) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
OAI322xp33_ASAP7_75t_L g728 ( .A1(n_676), .A2(n_729), .A3(n_731), .B1(n_732), .B2(n_733), .C1(n_735), .C2(n_738), .Y(n_728) );
AOI21xp33_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_686), .B(n_734), .Y(n_743) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_694), .C(n_706), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_722), .C(n_728), .D(n_740), .Y(n_711) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_742), .B(n_743), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule