module real_aes_6202_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g287 ( .A(n_0), .Y(n_287) );
AOI22xp33_ASAP7_75t_SL g126 ( .A1(n_1), .A2(n_33), .B1(n_127), .B2(n_131), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_2), .A2(n_31), .B1(n_200), .B2(n_212), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_3), .B(n_243), .Y(n_276) );
INVx1_ASAP7_75t_L g184 ( .A(n_4), .Y(n_184) );
AND2x6_ASAP7_75t_L g215 ( .A(n_4), .B(n_182), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_4), .B(n_507), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_5), .A2(n_80), .B1(n_81), .B2(n_162), .Y(n_79) );
INVx1_ASAP7_75t_L g162 ( .A(n_5), .Y(n_162) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_6), .A2(n_26), .B1(n_89), .B2(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g281 ( .A(n_7), .Y(n_281) );
INVx1_ASAP7_75t_L g196 ( .A(n_8), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_9), .B(n_204), .Y(n_203) );
AOI222xp33_ASAP7_75t_L g148 ( .A1(n_10), .A2(n_32), .B1(n_34), .B2(n_149), .C1(n_152), .C2(n_157), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_11), .B(n_241), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_12), .A2(n_66), .B1(n_136), .B2(n_140), .Y(n_135) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_13), .A2(n_236), .A3(n_240), .B1(n_242), .B2(n_243), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_14), .B(n_200), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_15), .A2(n_45), .B1(n_85), .B2(n_100), .Y(n_84) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_16), .A2(n_28), .B1(n_89), .B2(n_90), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_17), .B(n_241), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_18), .A2(n_42), .B1(n_200), .B2(n_212), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g252 ( .A1(n_19), .A2(n_61), .B1(n_200), .B2(n_204), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_20), .B(n_200), .Y(n_229) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_21), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_22), .B(n_192), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_23), .A2(n_46), .B1(n_143), .B2(n_146), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_24), .B(n_192), .Y(n_233) );
INVx2_ASAP7_75t_L g202 ( .A(n_25), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_27), .B(n_200), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g175 ( .A1(n_28), .A2(n_49), .B1(n_59), .B2(n_176), .C(n_177), .Y(n_175) );
INVxp67_ASAP7_75t_L g178 ( .A(n_28), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_29), .B(n_192), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_30), .A2(n_166), .B1(n_167), .B2(n_170), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_30), .Y(n_166) );
XOR2xp5_ASAP7_75t_L g514 ( .A(n_35), .B(n_80), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_36), .B(n_200), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_37), .A2(n_69), .B1(n_212), .B2(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_38), .B(n_200), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_39), .B(n_200), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_40), .A2(n_73), .B1(n_168), .B2(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_40), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_41), .B(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_SL g263 ( .A1(n_43), .A2(n_50), .B1(n_200), .B2(n_204), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_44), .A2(n_72), .B1(n_105), .B2(n_109), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_47), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_48), .B(n_200), .Y(n_300) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_49), .A2(n_64), .B1(n_89), .B2(n_90), .Y(n_88) );
INVxp67_ASAP7_75t_L g179 ( .A(n_49), .Y(n_179) );
INVx1_ASAP7_75t_L g513 ( .A(n_50), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_51), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g182 ( .A(n_52), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_53), .B(n_200), .Y(n_288) );
INVx1_ASAP7_75t_L g195 ( .A(n_54), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_55), .Y(n_176) );
AO32x2_ASAP7_75t_L g248 ( .A1(n_56), .A2(n_242), .A3(n_243), .B1(n_249), .B2(n_253), .Y(n_248) );
INVx1_ASAP7_75t_L g299 ( .A(n_57), .Y(n_299) );
INVx1_ASAP7_75t_L g224 ( .A(n_58), .Y(n_224) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_59), .A2(n_71), .B1(n_89), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_60), .B(n_204), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_62), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_63), .B(n_204), .Y(n_230) );
INVx2_ASAP7_75t_L g193 ( .A(n_65), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_67), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g163 ( .A1(n_68), .A2(n_164), .B1(n_165), .B2(n_171), .Y(n_163) );
INVx1_ASAP7_75t_L g171 ( .A(n_68), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_68), .B(n_204), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_70), .A2(n_76), .B1(n_204), .B2(n_205), .Y(n_262) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_70), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g168 ( .A(n_73), .Y(n_168) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_75), .B(n_204), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_172), .B1(n_185), .B2(n_496), .C(n_500), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_163), .Y(n_78) );
AOI22xp5_ASAP7_75t_SL g501 ( .A1(n_80), .A2(n_81), .B1(n_502), .B2(n_503), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND4xp75_ASAP7_75t_L g82 ( .A(n_83), .B(n_113), .C(n_134), .D(n_148), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_104), .Y(n_83) );
BUFx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
AND2x2_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_92), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_88), .B(n_93), .Y(n_103) );
INVx2_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
AND2x2_ASAP7_75t_L g130 ( .A(n_88), .B(n_97), .Y(n_130) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
INVx1_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
AND2x2_ASAP7_75t_L g118 ( .A(n_93), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
INVx1_ASAP7_75t_L g156 ( .A(n_93), .Y(n_156) );
AND2x4_ASAP7_75t_L g101 ( .A(n_95), .B(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g137 ( .A(n_95), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g141 ( .A(n_95), .B(n_118), .Y(n_141) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g108 ( .A(n_96), .B(n_99), .Y(n_108) );
OR2x2_ASAP7_75t_L g125 ( .A(n_96), .B(n_99), .Y(n_125) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g133 ( .A(n_97), .B(n_99), .Y(n_133) );
AND2x2_ASAP7_75t_L g155 ( .A(n_98), .B(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g112 ( .A(n_99), .Y(n_112) );
BUFx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OR2x6_ASAP7_75t_L g111 ( .A(n_103), .B(n_112), .Y(n_111) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx8_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2x1p5_ASAP7_75t_L g117 ( .A(n_108), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g147 ( .A(n_108), .B(n_138), .Y(n_147) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g129 ( .A(n_112), .Y(n_129) );
OA211x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_115), .B(n_120), .C(n_126), .Y(n_113) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g123 ( .A(n_118), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g138 ( .A(n_119), .B(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x6_ASAP7_75t_L g145 ( .A(n_124), .B(n_138), .Y(n_145) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x4_ASAP7_75t_L g154 ( .A(n_130), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g160 ( .A(n_130), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x6_ASAP7_75t_L g151 ( .A(n_133), .B(n_138), .Y(n_151) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_142), .Y(n_134) );
BUFx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx11_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx12f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_167), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
AND3x1_ASAP7_75t_SL g174 ( .A(n_175), .B(n_180), .C(n_183), .Y(n_174) );
INVxp67_ASAP7_75t_L g507 ( .A(n_175), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_180), .A2(n_499), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_180), .Y(n_518) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_181), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_181), .B(n_184), .Y(n_512) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_SL g517 ( .A(n_183), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_418), .Y(n_185) );
NAND5xp2_ASAP7_75t_L g186 ( .A(n_187), .B(n_337), .C(n_352), .D(n_378), .E(n_400), .Y(n_186) );
NOR2xp33_ASAP7_75t_SL g187 ( .A(n_188), .B(n_317), .Y(n_187) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_254), .B1(n_290), .B2(n_306), .C(n_307), .Y(n_188) );
NOR2xp33_ASAP7_75t_SL g189 ( .A(n_190), .B(n_244), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_190), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g494 ( .A(n_190), .Y(n_494) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_217), .Y(n_190) );
INVx1_ASAP7_75t_L g334 ( .A(n_191), .Y(n_334) );
AND2x2_ASAP7_75t_L g336 ( .A(n_191), .B(n_235), .Y(n_336) );
AND2x2_ASAP7_75t_L g346 ( .A(n_191), .B(n_234), .Y(n_346) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_191), .Y(n_364) );
INVx1_ASAP7_75t_L g374 ( .A(n_191), .Y(n_374) );
OR2x2_ASAP7_75t_L g412 ( .A(n_191), .B(n_311), .Y(n_412) );
INVx2_ASAP7_75t_L g462 ( .A(n_191), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_191), .B(n_310), .Y(n_479) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_197), .B(n_216), .Y(n_191) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_192), .A2(n_221), .B(n_233), .Y(n_220) );
INVx2_ASAP7_75t_L g253 ( .A(n_192), .Y(n_253) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AND2x2_ASAP7_75t_L g241 ( .A(n_193), .B(n_194), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_209), .B(n_215), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_203), .B(n_206), .Y(n_198) );
INVx3_ASAP7_75t_L g223 ( .A(n_200), .Y(n_223) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g212 ( .A(n_201), .Y(n_212) );
BUFx3_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g205 ( .A(n_202), .Y(n_205) );
INVx1_ASAP7_75t_L g275 ( .A(n_202), .Y(n_275) );
INVx2_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_208), .Y(n_214) );
INVx3_ASAP7_75t_L g227 ( .A(n_208), .Y(n_227) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_208), .Y(n_232) );
AND2x2_ASAP7_75t_L g499 ( .A(n_208), .B(n_275), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g298 ( .A1(n_213), .A2(n_286), .B(n_299), .C(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_214), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
OAI22xp5_ASAP7_75t_SL g249 ( .A1(n_214), .A2(n_227), .B1(n_250), .B2(n_252), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_214), .A2(n_238), .B1(n_262), .B2(n_263), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_215), .A2(n_222), .B(n_228), .Y(n_221) );
BUFx3_ASAP7_75t_L g242 ( .A(n_215), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_215), .A2(n_268), .B(n_271), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_215), .A2(n_280), .B(n_285), .Y(n_279) );
AND2x4_ASAP7_75t_L g498 ( .A(n_215), .B(n_499), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g217 ( .A(n_218), .B(n_234), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_219), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_219), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_219), .B(n_334), .Y(n_394) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_220), .Y(n_246) );
INVx2_ASAP7_75t_L g311 ( .A(n_220), .Y(n_311) );
OR2x2_ASAP7_75t_L g373 ( .A(n_220), .B(n_374), .Y(n_373) );
O2A1O1Ixp5_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B(n_225), .C(n_226), .Y(n_222) );
INVx2_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_226), .A2(n_269), .B(n_270), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_226), .A2(n_296), .B(n_297), .Y(n_295) );
INVx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
INVx4_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g312 ( .A(n_234), .B(n_248), .Y(n_312) );
AND2x2_ASAP7_75t_L g329 ( .A(n_234), .B(n_309), .Y(n_329) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g247 ( .A(n_235), .B(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g332 ( .A(n_235), .Y(n_332) );
AND2x2_ASAP7_75t_L g461 ( .A(n_235), .B(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_238), .A2(n_272), .B(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_238), .A2(n_286), .B(n_287), .C(n_288), .Y(n_285) );
INVx2_ASAP7_75t_L g278 ( .A(n_240), .Y(n_278) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_241), .Y(n_243) );
NAND3xp33_ASAP7_75t_L g260 ( .A(n_242), .B(n_261), .C(n_264), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_242), .A2(n_295), .B(n_298), .Y(n_294) );
INVx4_ASAP7_75t_L g264 ( .A(n_243), .Y(n_264) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_267), .B(n_276), .Y(n_266) );
INVx1_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
AND2x2_ASAP7_75t_L g424 ( .A(n_245), .B(n_312), .Y(n_424) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g425 ( .A(n_246), .B(n_336), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_247), .A2(n_393), .B(n_395), .C(n_397), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_247), .B(n_393), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_247), .A2(n_323), .B1(n_466), .B2(n_467), .C(n_469), .Y(n_465) );
INVx1_ASAP7_75t_L g309 ( .A(n_248), .Y(n_309) );
INVx1_ASAP7_75t_L g345 ( .A(n_248), .Y(n_345) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_265), .Y(n_255) );
AND2x2_ASAP7_75t_L g371 ( .A(n_256), .B(n_316), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_256), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_257), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g463 ( .A(n_257), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g495 ( .A(n_257), .Y(n_495) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g325 ( .A(n_258), .Y(n_325) );
AND2x2_ASAP7_75t_L g351 ( .A(n_258), .B(n_305), .Y(n_351) );
NOR2x1_ASAP7_75t_L g360 ( .A(n_258), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_258), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
AO21x1_ASAP7_75t_L g302 ( .A1(n_261), .A2(n_264), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_265), .B(n_407), .Y(n_442) );
INVx1_ASAP7_75t_SL g446 ( .A(n_265), .Y(n_446) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_277), .Y(n_265) );
INVx3_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
AND2x2_ASAP7_75t_L g316 ( .A(n_266), .B(n_293), .Y(n_316) );
AND2x2_ASAP7_75t_L g338 ( .A(n_266), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g383 ( .A(n_266), .B(n_377), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_266), .B(n_315), .Y(n_464) );
INVx2_ASAP7_75t_L g286 ( .A(n_274), .Y(n_286) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_277), .B(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_277), .B(n_377), .Y(n_376) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_289), .Y(n_277) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_278), .A2(n_294), .B(n_301), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_283), .C(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_304), .Y(n_291) );
INVx1_ASAP7_75t_L g356 ( .A(n_292), .Y(n_356) );
AND2x2_ASAP7_75t_L g398 ( .A(n_292), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_292), .B(n_319), .Y(n_404) );
AOI21xp5_ASAP7_75t_SL g478 ( .A1(n_292), .A2(n_310), .B(n_333), .Y(n_478) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_302), .Y(n_292) );
OR2x2_ASAP7_75t_L g321 ( .A(n_293), .B(n_302), .Y(n_321) );
AND2x2_ASAP7_75t_L g368 ( .A(n_293), .B(n_305), .Y(n_368) );
INVx2_ASAP7_75t_L g377 ( .A(n_293), .Y(n_377) );
INVx1_ASAP7_75t_L g483 ( .A(n_293), .Y(n_483) );
AND2x2_ASAP7_75t_L g407 ( .A(n_302), .B(n_377), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_302), .Y(n_432) );
AND2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_325), .Y(n_341) );
AND2x2_ASAP7_75t_L g353 ( .A(n_304), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_SL g471 ( .A(n_304), .Y(n_471) );
INVx2_ASAP7_75t_L g361 ( .A(n_305), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_305), .B(n_315), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_305), .B(n_483), .Y(n_482) );
OAI21xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_313), .Y(n_307) );
AND2x2_ASAP7_75t_L g414 ( .A(n_308), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g468 ( .A(n_308), .Y(n_468) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g388 ( .A(n_309), .Y(n_388) );
BUFx2_ASAP7_75t_L g487 ( .A(n_309), .Y(n_487) );
BUFx2_ASAP7_75t_L g358 ( .A(n_310), .Y(n_358) );
AND2x2_ASAP7_75t_L g460 ( .A(n_310), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g443 ( .A(n_311), .Y(n_443) );
AND2x4_ASAP7_75t_L g370 ( .A(n_312), .B(n_333), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_312), .B(n_394), .Y(n_406) );
AOI32xp33_ASAP7_75t_L g330 ( .A1(n_313), .A2(n_331), .A3(n_333), .B1(n_335), .B2(n_336), .Y(n_330) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx3_ASAP7_75t_L g319 ( .A(n_314), .Y(n_319) );
OR2x2_ASAP7_75t_L g455 ( .A(n_314), .B(n_411), .Y(n_455) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g324 ( .A(n_315), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g431 ( .A(n_315), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g323 ( .A(n_316), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g335 ( .A(n_316), .B(n_325), .Y(n_335) );
INVx1_ASAP7_75t_L g456 ( .A(n_316), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_316), .B(n_431), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B(n_326), .C(n_330), .Y(n_317) );
OAI322xp33_ASAP7_75t_L g426 ( .A1(n_318), .A2(n_363), .A3(n_427), .B1(n_429), .B2(n_433), .C1(n_434), .C2(n_438), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVxp67_ASAP7_75t_L g391 ( .A(n_319), .Y(n_391) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g445 ( .A(n_321), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_321), .B(n_361), .Y(n_492) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
OR2x2_ASAP7_75t_L g470 ( .A(n_325), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_328), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_358), .Y(n_379) );
AND2x2_ASAP7_75t_L g450 ( .A(n_329), .B(n_363), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_329), .B(n_437), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_331), .A2(n_338), .B1(n_341), .B2(n_342), .C(n_347), .Y(n_337) );
OR2x2_ASAP7_75t_L g348 ( .A(n_331), .B(n_344), .Y(n_348) );
AND2x2_ASAP7_75t_L g436 ( .A(n_331), .B(n_437), .Y(n_436) );
AOI32xp33_ASAP7_75t_L g475 ( .A1(n_331), .A2(n_361), .A3(n_476), .B1(n_477), .B2(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_332), .B(n_368), .C(n_391), .Y(n_409) );
AND2x2_ASAP7_75t_L g435 ( .A(n_332), .B(n_428), .Y(n_435) );
INVxp67_ASAP7_75t_L g415 ( .A(n_333), .Y(n_415) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_336), .B(n_388), .Y(n_444) );
INVx2_ASAP7_75t_L g454 ( .A(n_336), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_336), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g423 ( .A(n_339), .Y(n_423) );
OR2x2_ASAP7_75t_L g349 ( .A(n_340), .B(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_342), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_345), .Y(n_428) );
AND2x2_ASAP7_75t_L g387 ( .A(n_346), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g433 ( .A(n_346), .Y(n_433) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_346), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AOI21xp33_ASAP7_75t_SL g372 ( .A1(n_348), .A2(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g466 ( .A(n_351), .B(n_376), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B(n_365), .C(n_372), .Y(n_352) );
AND2x2_ASAP7_75t_L g396 ( .A(n_354), .B(n_364), .Y(n_396) );
INVx2_ASAP7_75t_L g411 ( .A(n_354), .Y(n_411) );
OR2x2_ASAP7_75t_L g449 ( .A(n_354), .B(n_412), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_354), .B(n_492), .Y(n_491) );
AOI211xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_357), .B(n_359), .C(n_362), .Y(n_355) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_358), .B(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_359), .A2(n_454), .B(n_478), .C(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g417 ( .A(n_361), .B(n_407), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_366), .B(n_369), .Y(n_365) );
INVxp33_ASAP7_75t_L g473 ( .A(n_367), .Y(n_473) );
AND2x2_ASAP7_75t_L g452 ( .A(n_368), .B(n_431), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_373), .A2(n_435), .B(n_436), .Y(n_434) );
OAI322xp33_ASAP7_75t_L g453 ( .A1(n_375), .A2(n_454), .A3(n_455), .B1(n_456), .B2(n_457), .C1(n_459), .C2(n_463), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_385), .B2(n_389), .C(n_392), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g430 ( .A(n_383), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g474 ( .A(n_387), .Y(n_474) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_390), .B(n_410), .Y(n_476) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g439 ( .A(n_399), .B(n_407), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_403), .A2(n_420), .B1(n_424), .B2(n_425), .C(n_426), .Y(n_419) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_407), .B(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_413), .B2(n_416), .Y(n_408) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx2_ASAP7_75t_SL g437 ( .A(n_412), .Y(n_437) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND5xp2_ASAP7_75t_L g418 ( .A(n_419), .B(n_440), .C(n_465), .D(n_475), .E(n_485), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_421), .B(n_423), .Y(n_420) );
NOR4xp25_ASAP7_75t_L g493 ( .A(n_422), .B(n_428), .C(n_494), .D(n_495), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_425), .A2(n_486), .B1(n_488), .B2(n_490), .C(n_493), .Y(n_485) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
OAI322xp33_ASAP7_75t_L g441 ( .A1(n_435), .A2(n_442), .A3(n_443), .B1(n_444), .B2(n_445), .C1(n_447), .C2(n_451), .Y(n_441) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_453), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g486 ( .A(n_461), .B(n_487), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI322xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_504), .A3(n_508), .B1(n_509), .B2(n_513), .C1(n_514), .C2(n_515), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_502), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
endmodule