module fake_jpeg_31675_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_55),
.Y(n_129)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_60),
.B(n_77),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_61),
.Y(n_115)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_62),
.Y(n_156)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_19),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_71),
.A2(n_73),
.B(n_24),
.Y(n_152)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_21),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_100),
.Y(n_124)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_104),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_19),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_35),
.B1(n_33),
.B2(n_43),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_130),
.B1(n_74),
.B2(n_54),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_43),
.C(n_33),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_152),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_26),
.B1(n_37),
.B2(n_44),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_62),
.B(n_34),
.CON(n_131),
.SN(n_131)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_23),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_135),
.B(n_144),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_26),
.B1(n_37),
.B2(n_44),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_142),
.B1(n_83),
.B2(n_67),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_73),
.A2(n_26),
.B1(n_103),
.B2(n_44),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_23),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_64),
.B(n_48),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_161),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_78),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_158),
.B(n_162),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_90),
.A2(n_38),
.B1(n_48),
.B2(n_27),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_55),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_55),
.B(n_38),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_168),
.Y(n_222)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_166),
.B(n_204),
.Y(n_269)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_37),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_169),
.B(n_192),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_177),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_44),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_184),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_174),
.A2(n_216),
.B(n_121),
.C(n_24),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_176),
.A2(n_188),
.B1(n_203),
.B2(n_143),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_25),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_25),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_179),
.B(n_181),
.Y(n_260)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_180),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_45),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_44),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_185),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_187),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_59),
.B1(n_57),
.B2(n_66),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_114),
.Y(n_192)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_194),
.B(n_201),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_126),
.Y(n_199)
);

BUFx4f_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_105),
.B(n_40),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_110),
.A2(n_86),
.B1(n_95),
.B2(n_94),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_205),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_40),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_213),
.B1(n_214),
.B2(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_34),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_208),
.B(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_215),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_126),
.A2(n_89),
.B1(n_88),
.B2(n_96),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_24),
.B1(n_121),
.B2(n_3),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_152),
.A2(n_49),
.B(n_45),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_130),
.B(n_49),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_149),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_106),
.B(n_28),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_146),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_220),
.A2(n_221),
.B1(n_213),
.B2(n_204),
.Y(n_250)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_154),
.B1(n_139),
.B2(n_146),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_194),
.A2(n_133),
.B1(n_139),
.B2(n_154),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_233),
.B1(n_244),
.B2(n_220),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_121),
.B(n_106),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_229),
.A2(n_246),
.B(n_250),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_28),
.B(n_24),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_195),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_138),
.C(n_143),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_237),
.C(n_259),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_138),
.C(n_111),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_179),
.B(n_202),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_173),
.A2(n_111),
.B1(n_24),
.B2(n_106),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_248),
.A2(n_255),
.B1(n_258),
.B2(n_2),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_190),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_189),
.A2(n_9),
.B1(n_17),
.B2(n_15),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_171),
.B(n_18),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_181),
.B(n_1),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_177),
.B(n_1),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_216),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_272),
.B(n_279),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_220),
.B1(n_221),
.B2(n_214),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_276),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_200),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_282),
.Y(n_317)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_278),
.A2(n_225),
.B1(n_248),
.B2(n_231),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_228),
.B(n_175),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_280),
.B(n_281),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_238),
.B(n_165),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_164),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_260),
.A2(n_167),
.B1(n_218),
.B2(n_199),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_287),
.B1(n_288),
.B2(n_304),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_166),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_284),
.B(n_293),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_182),
.B1(n_191),
.B2(n_183),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_251),
.A2(n_186),
.B1(n_196),
.B2(n_207),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_232),
.B(n_178),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_193),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_295),
.Y(n_350)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_227),
.B(n_170),
.Y(n_293)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

BUFx24_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_204),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_230),
.B(n_12),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_296),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_223),
.Y(n_300)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_257),
.A2(n_12),
.B(n_18),
.C(n_14),
.Y(n_302)
);

XNOR2x2_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_241),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_303),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_251),
.A2(n_213),
.B1(n_18),
.B2(n_14),
.Y(n_304)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_305),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_13),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_309),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_3),
.Y(n_309)
);

BUFx8_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_310),
.Y(n_352)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_312),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_237),
.C(n_235),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_331),
.C(n_277),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_302),
.C(n_309),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_233),
.B1(n_254),
.B2(n_246),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_329),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_341),
.B1(n_286),
.B2(n_285),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_297),
.A2(n_244),
.B1(n_259),
.B2(n_262),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_298),
.C(n_289),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_266),
.B1(n_261),
.B2(n_234),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_342),
.Y(n_356)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_274),
.A2(n_252),
.A3(n_239),
.B1(n_268),
.B2(n_247),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_272),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_278),
.A2(n_234),
.B1(n_256),
.B2(n_249),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_283),
.B1(n_287),
.B2(n_291),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_280),
.A2(n_239),
.B1(n_264),
.B2(n_236),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_345),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_277),
.B(n_236),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_282),
.A2(n_264),
.B1(n_247),
.B2(n_245),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_310),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_333),
.Y(n_354)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_357),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_338),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_365),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_290),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_336),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_360),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_361),
.A2(n_363),
.B(n_364),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_304),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_362),
.B(n_382),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_313),
.B(n_273),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_338),
.A2(n_313),
.B(n_271),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_345),
.Y(n_365)
);

INVx3_ASAP7_75t_SL g366 ( 
.A(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_367),
.A2(n_373),
.B1(n_386),
.B2(n_348),
.Y(n_404)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_368),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_270),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_369),
.Y(n_419)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_343),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_311),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_374),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_337),
.A2(n_252),
.B1(n_307),
.B2(n_300),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_334),
.B(n_276),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_378),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_317),
.B(n_305),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_347),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_383),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_310),
.Y(n_380)
);

AO21x1_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_387),
.B(n_324),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_303),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_385),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_292),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_320),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_314),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_384),
.B(n_314),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_337),
.Y(n_385)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_294),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_388),
.B(n_352),
.Y(n_389)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

FAx1_ASAP7_75t_SL g391 ( 
.A(n_371),
.B(n_331),
.CI(n_322),
.CON(n_391),
.SN(n_391)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_395),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_360),
.B(n_316),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_380),
.A2(n_348),
.B1(n_328),
.B2(n_341),
.Y(n_396)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

OA22x2_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_411),
.B1(n_418),
.B2(n_381),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_364),
.A2(n_358),
.B(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_417),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_367),
.B1(n_366),
.B2(n_355),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_363),
.A2(n_326),
.B1(n_342),
.B2(n_321),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_369),
.B(n_321),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_359),
.C(n_379),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_410),
.Y(n_428)
);

AO22x1_ASAP7_75t_L g411 ( 
.A1(n_386),
.A2(n_325),
.B1(n_332),
.B2(n_329),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_372),
.A2(n_326),
.B1(n_325),
.B2(n_319),
.Y(n_412)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_412),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_3),
.C(n_4),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_356),
.A2(n_330),
.B(n_319),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_387),
.A2(n_355),
.B1(n_365),
.B2(n_374),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_420),
.A2(n_430),
.B1(n_434),
.B2(n_436),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_356),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_443),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_395),
.B(n_354),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_437),
.Y(n_449)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_376),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_427),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_376),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_378),
.B1(n_384),
.B2(n_375),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_413),
.A2(n_366),
.B1(n_370),
.B2(n_388),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_431),
.A2(n_414),
.B1(n_390),
.B2(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_445),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_275),
.Y(n_433)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_399),
.A2(n_383),
.B1(n_320),
.B2(n_301),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_411),
.A2(n_330),
.B1(n_357),
.B2(n_368),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_389),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_397),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_439),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_411),
.A2(n_330),
.B1(n_357),
.B2(n_368),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_440),
.A2(n_396),
.B1(n_414),
.B2(n_390),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_394),
.B(n_253),
.Y(n_441)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_253),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_405),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_408),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_412),
.C(n_418),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_456),
.C(n_460),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_416),
.C(n_417),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_426),
.A2(n_402),
.B(n_392),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_400),
.B(n_420),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_SL g458 ( 
.A(n_438),
.B(n_401),
.C(n_416),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_SL g483 ( 
.A(n_458),
.B(n_419),
.C(n_432),
.Y(n_483)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_403),
.C(n_393),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_403),
.C(n_393),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_461),
.B(n_465),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_466),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_446),
.A2(n_423),
.B1(n_442),
.B2(n_426),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_467),
.A2(n_483),
.B1(n_432),
.B2(n_448),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_449),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_474),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_476),
.B(n_436),
.Y(n_488)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_450),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_457),
.A2(n_400),
.B(n_440),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_442),
.B1(n_423),
.B2(n_428),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_477),
.A2(n_463),
.B1(n_451),
.B2(n_452),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_419),
.Y(n_479)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_443),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_447),
.Y(n_490)
);

AOI21xp33_ASAP7_75t_L g481 ( 
.A1(n_458),
.A2(n_432),
.B(n_398),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_481),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_450),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_474),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_486),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_475),
.B(n_453),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_455),
.C(n_460),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_487),
.B(n_493),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_490),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_496),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_462),
.C(n_456),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_494),
.A2(n_498),
.B1(n_468),
.B2(n_451),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_462),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_471),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_472),
.B(n_465),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_444),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_488),
.B(n_490),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_498),
.A2(n_468),
.B1(n_482),
.B2(n_483),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_506),
.B(n_507),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_473),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_509),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_478),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_407),
.Y(n_517)
);

AOI31xp33_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_492),
.A3(n_478),
.B(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_512),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_506),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_516),
.A2(n_517),
.B1(n_502),
.B2(n_409),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_407),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_518),
.B(n_409),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_501),
.C(n_502),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_519),
.A2(n_520),
.B(n_522),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_523),
.A2(n_511),
.B1(n_514),
.B2(n_500),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_524),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_516),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_522),
.B(n_5),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_527),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_529),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_525),
.Y(n_531)
);

AOI221xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_528),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_4),
.B(n_5),
.Y(n_533)
);


endmodule