module fake_jpeg_30080_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_22),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_20),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_26),
.B(n_19),
.C(n_18),
.Y(n_48)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_25),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_50),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_67),
.Y(n_80)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_16),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_72),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_20),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_82),
.B(n_43),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_57),
.B1(n_62),
.B2(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_24),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_65),
.C(n_58),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_23),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_65),
.B1(n_55),
.B2(n_56),
.Y(n_99)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_6),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_6),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_58),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_98),
.C(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_72),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_25),
.A3(n_3),
.B1(n_0),
.B2(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_94),
.C(n_86),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_110),
.C(n_100),
.Y(n_115)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_109),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_100),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_120),
.C(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_87),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_122),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_115),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_102),
.B1(n_91),
.B2(n_113),
.Y(n_127)
);

AOI31xp67_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_102),
.A3(n_101),
.B(n_120),
.Y(n_131)
);

BUFx4f_ASAP7_75t_SL g128 ( 
.A(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_104),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_122),
.Y(n_135)
);

AOI31xp67_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_125),
.A3(n_118),
.B(n_128),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_100),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_126),
.C(n_96),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_133),
.A3(n_102),
.B1(n_87),
.B2(n_81),
.C1(n_71),
.C2(n_45),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_64),
.C(n_76),
.Y(n_140)
);

OA21x2_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_138),
.B(n_76),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_45),
.Y(n_142)
);


endmodule