module fake_jpeg_20357_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_46),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_48),
.B1(n_53),
.B2(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_51),
.B1(n_40),
.B2(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_48),
.B1(n_53),
.B2(n_52),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_79),
.B1(n_83),
.B2(n_66),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_46),
.B1(n_50),
.B2(n_23),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_99),
.Y(n_104)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_5),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_95),
.C(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_76),
.C(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_105),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_103),
.B(n_101),
.Y(n_110)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_111),
.A3(n_109),
.B1(n_96),
.B2(n_97),
.C(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_104),
.C(n_99),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_7),
.C(n_9),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_10),
.B(n_14),
.Y(n_114)
);

OAI21x1_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_17),
.B(n_18),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_27),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_29),
.B(n_30),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_32),
.C(n_35),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_36),
.Y(n_119)
);


endmodule