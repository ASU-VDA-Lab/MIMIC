module fake_ariane_2730_n_2328 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2328);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2328;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_221;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_60),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_29),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_105),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_40),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_41),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_58),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_73),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_84),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_189),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_108),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_89),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_117),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_81),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_129),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_135),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_62),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_36),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_75),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_113),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_127),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_84),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_38),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_85),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_152),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_46),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_33),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_65),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_126),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_24),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_10),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_6),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_99),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_171),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_67),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_58),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_50),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_55),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_31),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_128),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_81),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_70),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_19),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_103),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_190),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_161),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_28),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_119),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_142),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_185),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_151),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_107),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_9),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_131),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_45),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_153),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_11),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_88),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_209),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_57),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_217),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_14),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_40),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_20),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_194),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_144),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_150),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_214),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_157),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_204),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_78),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_20),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_19),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_11),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_122),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_23),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_71),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_191),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_116),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_201),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_140),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_93),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_73),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_62),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_139),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_79),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_25),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_13),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_56),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_77),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_121),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_14),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_21),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_137),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_32),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_199),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_75),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_47),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_47),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_133),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_115),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_43),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_23),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_49),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_213),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_167),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_61),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_87),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_59),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_59),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_18),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_18),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_37),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_25),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_154),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_68),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_76),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_35),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_179),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_147),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_195),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_205),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_67),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_78),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_17),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_54),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_210),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_158),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_36),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_168),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_41),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_55),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_28),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_91),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_69),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_54),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_177),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_186),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_42),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_74),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_79),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_3),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_114),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_57),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_130),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_118),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_97),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_89),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_202),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_80),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_51),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_101),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_169),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_207),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_106),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_94),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_98),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_132),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_99),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_39),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_95),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_86),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_148),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_44),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_165),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_7),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_183),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_92),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_72),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_421),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_279),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_273),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_280),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_220),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_349),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_219),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_219),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_229),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_291),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_229),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_233),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_233),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_295),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_301),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_311),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_366),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_399),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_247),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_247),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_225),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_248),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_416),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_258),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_227),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_258),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_349),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_239),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_232),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_252),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_256),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_287),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_259),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_261),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_349),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_385),
.B(n_0),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_267),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_268),
.Y(n_477)
);

INVxp33_ASAP7_75t_SL g478 ( 
.A(n_270),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_267),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_241),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_271),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_274),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_272),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_303),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_272),
.B(n_0),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_328),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_278),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_275),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_275),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_304),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_304),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_353),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_224),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_363),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_317),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_317),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_287),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_375),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_375),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_321),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_236),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_321),
.B(n_1),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_324),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_281),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_284),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_286),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_287),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_315),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_288),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_324),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_333),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_333),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_289),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_360),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_290),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_360),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_236),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_341),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_224),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_375),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_292),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_296),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_341),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_381),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_306),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_237),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_383),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_230),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_308),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_383),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_388),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_392),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_309),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_R g536 ( 
.A(n_221),
.B(n_100),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_310),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_287),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_360),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_287),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_237),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_392),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_230),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_405),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_314),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_540),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_467),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_442),
.A2(n_234),
.B1(n_426),
.B2(n_222),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_540),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_237),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_502),
.B(n_485),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_471),
.A2(n_405),
.B(n_307),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_432),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_471),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_508),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_434),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_466),
.B(n_253),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_439),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_497),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_497),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_454),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_507),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_507),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_441),
.B(n_285),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_441),
.B(n_285),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_444),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_446),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_485),
.B(n_287),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_448),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_448),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_527),
.B(n_253),
.Y(n_592)
);

NOR2xp67_ASAP7_75t_L g593 ( 
.A(n_449),
.B(n_415),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_449),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_450),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_440),
.B(n_414),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_456),
.B(n_253),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_462),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_456),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_457),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_457),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_447),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_469),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_459),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_451),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_452),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_459),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_460),
.B(n_415),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_514),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_453),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_455),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_470),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_461),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_480),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_465),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_473),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_477),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_481),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_465),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_476),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_487),
.Y(n_624)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_476),
.A2(n_307),
.B(n_298),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_479),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_504),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_474),
.B(n_298),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_479),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_483),
.Y(n_630)
);

OA21x2_ASAP7_75t_L g631 ( 
.A1(n_483),
.A2(n_307),
.B(n_298),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_488),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_488),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_489),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_541),
.B(n_305),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_609),
.B(n_260),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_549),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_609),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_609),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_609),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_549),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_592),
.B(n_498),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_611),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_592),
.B(n_499),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_501),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_609),
.B(n_589),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_592),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_609),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_549),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_611),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_609),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_586),
.B(n_501),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_468),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_609),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_586),
.B(n_517),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_517),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_597),
.A2(n_443),
.B1(n_437),
.B2(n_472),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_260),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_546),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_546),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_597),
.B(n_520),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_629),
.B(n_478),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_546),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_552),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_619),
.B(n_505),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_618),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_552),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_590),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_635),
.B(n_520),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_590),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_560),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_629),
.B(n_506),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_591),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_591),
.Y(n_682)
);

NAND3x1_ASAP7_75t_L g683 ( 
.A(n_628),
.B(n_238),
.C(n_235),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_548),
.A2(n_475),
.B1(n_529),
.B2(n_519),
.Y(n_684)
);

OR2x2_ASAP7_75t_SL g685 ( 
.A(n_551),
.B(n_458),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_628),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_629),
.B(n_509),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_547),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_635),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_604),
.A2(n_475),
.B1(n_374),
.B2(n_342),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_552),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_559),
.Y(n_692)
);

INVxp33_ASAP7_75t_L g693 ( 
.A(n_551),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_550),
.B(n_489),
.Y(n_694)
);

INVx5_ASAP7_75t_L g695 ( 
.A(n_565),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_550),
.B(n_569),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_629),
.B(n_490),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_550),
.B(n_493),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_591),
.B(n_594),
.Y(n_699)
);

BUFx4f_ASAP7_75t_L g700 ( 
.A(n_625),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_625),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_559),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_559),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_559),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_601),
.B(n_513),
.Y(n_705)
);

AND3x4_ASAP7_75t_L g706 ( 
.A(n_593),
.B(n_346),
.C(n_305),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_604),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_594),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_569),
.B(n_490),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_491),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_548),
.A2(n_588),
.B1(n_631),
.B2(n_625),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_547),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_617),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_601),
.B(n_515),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_596),
.B(n_491),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_596),
.B(n_260),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_559),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_562),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_604),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_562),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_602),
.B(n_521),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_562),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_596),
.B(n_495),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_630),
.B(n_260),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_598),
.B(n_320),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_630),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_630),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_625),
.B(n_631),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_598),
.B(n_543),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_525),
.C(n_522),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_615),
.B(n_464),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_618),
.B(n_495),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_598),
.B(n_496),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_571),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_562),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_632),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_560),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_585),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_575),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_530),
.Y(n_741)
);

INVx4_ASAP7_75t_SL g742 ( 
.A(n_565),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_632),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_605),
.B(n_535),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_615),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_565),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_632),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_605),
.B(n_537),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_615),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_585),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_620),
.A2(n_234),
.B1(n_426),
.B2(n_222),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_634),
.Y(n_752)
);

INVxp67_ASAP7_75t_SL g753 ( 
.A(n_593),
.Y(n_753)
);

INVx4_ASAP7_75t_SL g754 ( 
.A(n_565),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_634),
.B(n_496),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_565),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_620),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_565),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_545),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_575),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_608),
.B(n_516),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_634),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_556),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_585),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_556),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_613),
.B(n_500),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_613),
.B(n_500),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_562),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_539),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_598),
.B(n_385),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_598),
.B(n_503),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_557),
.Y(n_772)
);

BUFx4f_ASAP7_75t_L g773 ( 
.A(n_625),
.Y(n_773)
);

NAND3x1_ASAP7_75t_L g774 ( 
.A(n_580),
.B(n_238),
.C(n_235),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_598),
.B(n_503),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_621),
.B(n_438),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_622),
.B(n_435),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_623),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_557),
.Y(n_779)
);

AO22x2_ASAP7_75t_L g780 ( 
.A1(n_588),
.A2(n_511),
.B1(n_512),
.B2(n_510),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_565),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_617),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_558),
.Y(n_783)
);

OAI221xp5_ASAP7_75t_L g784 ( 
.A1(n_580),
.A2(n_246),
.B1(n_249),
.B2(n_262),
.C(n_264),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_621),
.A2(n_318),
.B1(n_326),
.B2(n_325),
.Y(n_785)
);

BUFx8_ASAP7_75t_SL g786 ( 
.A(n_603),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_585),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_558),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_564),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_623),
.B(n_510),
.Y(n_790)
);

AND2x6_ASAP7_75t_SL g791 ( 
.A(n_786),
.B(n_246),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_672),
.B(n_626),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_745),
.B(n_624),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_707),
.Y(n_795)
);

NAND2x1_ASAP7_75t_L g796 ( 
.A(n_679),
.B(n_626),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_770),
.B(n_583),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_733),
.B(n_583),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_743),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_643),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_700),
.B(n_624),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_761),
.B(n_627),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_743),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_769),
.B(n_627),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_706),
.A2(n_554),
.B1(n_631),
.B2(n_625),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_700),
.B(n_773),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_745),
.B(n_599),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_777),
.B(n_249),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_733),
.B(n_610),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_700),
.B(n_553),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_660),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_686),
.B(n_610),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_654),
.B(n_587),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_706),
.A2(n_554),
.B1(n_631),
.B2(n_512),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_668),
.B(n_587),
.Y(n_816)
);

AND2x6_ASAP7_75t_SL g817 ( 
.A(n_705),
.B(n_262),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_739),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_770),
.B(n_587),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_697),
.A2(n_699),
.B(n_656),
.C(n_674),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_773),
.B(n_553),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_726),
.A2(n_554),
.B1(n_631),
.B2(n_518),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_667),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_726),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_715),
.B(n_587),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_773),
.B(n_553),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_679),
.B(n_599),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_696),
.B(n_564),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_726),
.A2(n_554),
.B1(n_631),
.B2(n_518),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_667),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_722),
.A2(n_536),
.B1(n_600),
.B2(n_595),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_720),
.B(n_603),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_606),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_741),
.B(n_595),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_726),
.A2(n_554),
.B1(n_523),
.B2(n_524),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_674),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_726),
.A2(n_554),
.B1(n_523),
.B2(n_524),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_660),
.Y(n_838)
);

AND2x6_ASAP7_75t_SL g839 ( 
.A(n_744),
.B(n_264),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_749),
.B(n_607),
.C(n_606),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_677),
.A2(n_567),
.B(n_566),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_748),
.B(n_595),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_677),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_739),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_778),
.A2(n_567),
.B1(n_568),
.B2(n_566),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_759),
.A2(n_600),
.B1(n_633),
.B2(n_595),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_679),
.B(n_600),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_681),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_681),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_750),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_749),
.B(n_600),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_648),
.B(n_633),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_646),
.B(n_653),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_651),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_682),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_701),
.B(n_633),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_701),
.B(n_660),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_735),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_657),
.B(n_658),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_750),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_SL g861 ( 
.A(n_659),
.B(n_484),
.C(n_482),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_701),
.B(n_633),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_648),
.B(n_568),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_750),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_642),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_732),
.B(n_607),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_734),
.B(n_511),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_689),
.B(n_526),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_689),
.B(n_526),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_680),
.B(n_528),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_682),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_708),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_732),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_687),
.B(n_528),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_660),
.B(n_531),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_671),
.B(n_612),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_764),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_642),
.B(n_531),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_660),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_688),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_642),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_708),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_645),
.B(n_532),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_711),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_707),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_645),
.B(n_532),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_676),
.B(n_533),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_645),
.B(n_533),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_778),
.A2(n_346),
.B1(n_347),
.B2(n_305),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_666),
.B(n_534),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_764),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_714),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_694),
.B(n_534),
.Y(n_893)
);

NOR2x2_ASAP7_75t_L g894 ( 
.A(n_770),
.B(n_346),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_694),
.B(n_542),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_638),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_764),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_709),
.B(n_542),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_726),
.A2(n_354),
.B1(n_544),
.B2(n_263),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_709),
.B(n_544),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_729),
.A2(n_561),
.B(n_555),
.Y(n_901)
);

BUFx5_ASAP7_75t_L g902 ( 
.A(n_639),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_676),
.B(n_320),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_696),
.A2(n_226),
.B1(n_228),
.B2(n_223),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_698),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_698),
.B(n_612),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_757),
.B(n_614),
.Y(n_907)
);

BUFx5_ASAP7_75t_L g908 ( 
.A(n_639),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_757),
.B(n_731),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_770),
.B(n_347),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_696),
.B(n_614),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_676),
.B(n_320),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_787),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_710),
.B(n_347),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_710),
.B(n_350),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_711),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_727),
.A2(n_370),
.B(n_395),
.C(n_350),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_735),
.B(n_616),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_787),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_734),
.B(n_350),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_734),
.A2(n_240),
.B1(n_242),
.B2(n_231),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_727),
.Y(n_922)
);

AO221x1_ASAP7_75t_L g923 ( 
.A1(n_751),
.A2(n_785),
.B1(n_690),
.B2(n_780),
.C(n_678),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_771),
.B(n_775),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_370),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_684),
.A2(n_265),
.B1(n_332),
.B2(n_236),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_370),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_782),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_397),
.B1(n_395),
.B2(n_338),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_780),
.A2(n_265),
.B1(n_332),
.B2(n_236),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_775),
.B(n_395),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_775),
.B(n_397),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_688),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_698),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_676),
.Y(n_935)
);

AND2x6_ASAP7_75t_SL g936 ( 
.A(n_740),
.B(n_266),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_737),
.A2(n_561),
.B(n_555),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_675),
.B(n_616),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_787),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_676),
.B(n_738),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_780),
.A2(n_265),
.B1(n_403),
.B2(n_332),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_730),
.B(n_397),
.Y(n_942)
);

O2A1O1Ixp5_ASAP7_75t_L g943 ( 
.A1(n_678),
.A2(n_561),
.B(n_563),
.C(n_555),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_730),
.B(n_572),
.Y(n_944)
);

BUFx12f_ASAP7_75t_SL g945 ( 
.A(n_730),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_753),
.B(n_486),
.Y(n_946)
);

INVx5_ASAP7_75t_L g947 ( 
.A(n_638),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_738),
.B(n_340),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_644),
.B(n_492),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_738),
.B(n_340),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_664),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_737),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_738),
.B(n_340),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_738),
.B(n_417),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_747),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_638),
.B(n_376),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_763),
.B(n_572),
.Y(n_957)
);

AND2x6_ASAP7_75t_SL g958 ( 
.A(n_740),
.B(n_266),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_664),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_638),
.B(n_376),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_678),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_765),
.B(n_572),
.Y(n_962)
);

INVx8_ASAP7_75t_L g963 ( 
.A(n_638),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_865),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_951),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_SL g966 ( 
.A(n_802),
.B(n_760),
.C(n_776),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_865),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_873),
.B(n_866),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_885),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_853),
.B(n_859),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_951),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_963),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_880),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_959),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_798),
.B(n_766),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_810),
.B(n_767),
.Y(n_977)
);

AO22x1_ASAP7_75t_L g978 ( 
.A1(n_804),
.A2(n_760),
.B1(n_858),
.B2(n_949),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_881),
.B(n_683),
.Y(n_979)
);

AO22x1_ASAP7_75t_L g980 ( 
.A1(n_858),
.A2(n_713),
.B1(n_494),
.B2(n_685),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_SL g981 ( 
.A(n_918),
.B(n_713),
.C(n_339),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_881),
.Y(n_982)
);

AND2x6_ASAP7_75t_SL g983 ( 
.A(n_907),
.B(n_876),
.Y(n_983)
);

AND3x2_ASAP7_75t_SL g984 ( 
.A(n_923),
.B(n_683),
.C(n_408),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_813),
.B(n_790),
.Y(n_985)
);

BUFx4f_ASAP7_75t_L g986 ( 
.A(n_794),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_824),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_870),
.B(n_765),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_824),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_938),
.A2(n_779),
.B1(n_783),
.B2(n_772),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_808),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_963),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_824),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_945),
.B(n_685),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_793),
.Y(n_995)
);

NAND3xp33_ASAP7_75t_SL g996 ( 
.A(n_840),
.B(n_344),
.C(n_329),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_806),
.B(n_747),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_823),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_880),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_874),
.B(n_772),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_819),
.B(n_779),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_890),
.B(n_878),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_800),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_963),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_883),
.B(n_783),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_886),
.B(n_888),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_793),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_819),
.B(n_788),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_854),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_928),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_836),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_843),
.A2(n_752),
.B(n_762),
.C(n_784),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_963),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_893),
.B(n_788),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_R g1016 ( 
.A(n_945),
.B(n_647),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_895),
.B(n_789),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_909),
.A2(n_789),
.B1(n_762),
.B2(n_752),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_848),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_832),
.B(n_911),
.C(n_827),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_905),
.B(n_780),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_827),
.B(n_365),
.C(n_361),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_833),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_818),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_818),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_898),
.B(n_716),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_896),
.B(n_728),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_844),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_849),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_838),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_844),
.Y(n_1031)
);

AND3x2_ASAP7_75t_SL g1032 ( 
.A(n_817),
.B(n_408),
.C(n_376),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_819),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_900),
.B(n_724),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_906),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_855),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_871),
.Y(n_1037)
);

INVx8_ASAP7_75t_L g1038 ( 
.A(n_819),
.Y(n_1038)
);

INVx6_ASAP7_75t_L g1039 ( 
.A(n_828),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_896),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_872),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_828),
.B(n_637),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_825),
.A2(n_755),
.B1(n_641),
.B2(n_650),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_828),
.B(n_712),
.Y(n_1044)
);

BUFx10_ASAP7_75t_L g1045 ( 
.A(n_946),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_807),
.B(n_265),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_809),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_934),
.B(n_637),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_795),
.B(n_641),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_910),
.B(n_774),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_838),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_882),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_884),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_868),
.B(n_665),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_850),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_924),
.B(n_650),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_916),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_838),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_869),
.B(n_665),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_806),
.B(n_662),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_850),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_933),
.B(n_662),
.Y(n_1062)
);

CKINVDCx8_ASAP7_75t_R g1063 ( 
.A(n_791),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_834),
.B(n_669),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_838),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_961),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_892),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_842),
.B(n_669),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_812),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_860),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_922),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_867),
.B(n_332),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_812),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_894),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_894),
.Y(n_1075)
);

AOI22x1_ASAP7_75t_L g1076 ( 
.A1(n_841),
.A2(n_663),
.B1(n_673),
.B2(n_670),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_867),
.B(n_670),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_792),
.B(n_851),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_851),
.B(n_673),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_896),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_879),
.Y(n_1081)
);

BUFx8_ASAP7_75t_L g1082 ( 
.A(n_799),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_801),
.B(n_663),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_914),
.B(n_691),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_910),
.B(n_774),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_860),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_864),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_856),
.A2(n_647),
.B(n_640),
.Y(n_1088)
);

CKINVDCx11_ASAP7_75t_R g1089 ( 
.A(n_936),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_952),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_861),
.B(n_661),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_879),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_915),
.B(n_691),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_801),
.B(n_640),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_955),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_SL g1096 ( 
.A(n_929),
.B(n_368),
.C(n_367),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_910),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_961),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_864),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_942),
.B(n_692),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_930),
.A2(n_661),
.B1(n_725),
.B2(n_717),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_839),
.B(n_717),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_904),
.B(n_372),
.C(n_371),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_902),
.B(n_640),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_814),
.B(n_692),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_816),
.B(n_702),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_877),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_917),
.B(n_384),
.C(n_378),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_863),
.B(n_702),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_910),
.Y(n_1110)
);

NOR2x1p5_ASAP7_75t_L g1111 ( 
.A(n_920),
.B(n_276),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_R g1112 ( 
.A(n_935),
.B(n_725),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_831),
.B(n_703),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_803),
.B(n_797),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_852),
.Y(n_1115)
);

OR2x6_ASAP7_75t_SL g1116 ( 
.A(n_889),
.B(n_386),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_957),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_797),
.A2(n_649),
.B1(n_655),
.B2(n_652),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_797),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_797),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_962),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_796),
.B(n_649),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_896),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_896),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_925),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_921),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_958),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_944),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_927),
.B(n_703),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_877),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_SL g1131 ( 
.A(n_845),
.B(n_403),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_931),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_891),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_932),
.B(n_704),
.Y(n_1134)
);

BUFx4f_ASAP7_75t_L g1135 ( 
.A(n_954),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_891),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_897),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_815),
.B(n_704),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_899),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_897),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_941),
.A2(n_649),
.B1(n_655),
.B2(n_652),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_947),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_913),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_913),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_926),
.B(n_718),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_856),
.B(n_652),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_919),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_917),
.B(n_390),
.C(n_387),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_947),
.B(n_742),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_919),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_846),
.B(n_718),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_857),
.B(n_954),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_902),
.B(n_655),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_947),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_947),
.B(n_935),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_939),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_R g1157 ( 
.A(n_935),
.B(n_636),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1076),
.A2(n_901),
.B(n_821),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_970),
.A2(n_821),
.B(n_811),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_988),
.A2(n_826),
.B1(n_811),
.B2(n_939),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_1001),
.A2(n_820),
.B(n_943),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_985),
.B(n_835),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1064),
.A2(n_826),
.B(n_862),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1083),
.A2(n_1094),
.B(n_1060),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1083),
.A2(n_729),
.B(n_937),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_1113),
.A2(n_721),
.A3(n_723),
.B(n_719),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_L g1167 ( 
.A(n_1023),
.B(n_947),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1138),
.A2(n_721),
.A3(n_723),
.B(n_719),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1094),
.A2(n_729),
.B(n_857),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1060),
.A2(n_960),
.B(n_956),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_972),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1068),
.A2(n_862),
.B(n_847),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1067),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1015),
.A2(n_847),
.B(n_940),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_976),
.B(n_977),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1003),
.B(n_837),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_989),
.Y(n_1177)
);

BUFx2_ASAP7_75t_R g1178 ( 
.A(n_1063),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1146),
.A2(n_768),
.A3(n_736),
.B(n_573),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1035),
.B(n_403),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1142),
.B(n_1002),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_968),
.B(n_875),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1017),
.A2(n_940),
.B(n_887),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_991),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1002),
.B(n_875),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1126),
.A2(n_887),
.B1(n_908),
.B2(n_902),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1056),
.A2(n_829),
.B(n_822),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1128),
.B(n_805),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1007),
.B(n_902),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1117),
.B(n_902),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_997),
.A2(n_956),
.B(n_960),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_986),
.B(n_403),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_997),
.A2(n_912),
.B(n_903),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_998),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1121),
.B(n_902),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_999),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1012),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1088),
.A2(n_912),
.B(n_903),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_SL g1199 ( 
.A1(n_989),
.A2(n_1149),
.B(n_1009),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_1142),
.B(n_948),
.Y(n_1200)
);

CKINVDCx16_ASAP7_75t_R g1201 ( 
.A(n_981),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1039),
.B(n_902),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1046),
.B(n_978),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1043),
.A2(n_950),
.B(n_948),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_972),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1151),
.A2(n_953),
.B(n_950),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_SL g1207 ( 
.A1(n_989),
.A2(n_953),
.B(n_408),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1104),
.A2(n_768),
.B(n_736),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1104),
.A2(n_561),
.B(n_555),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1105),
.A2(n_636),
.B(n_746),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_990),
.A2(n_1018),
.B(n_1020),
.C(n_1026),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1019),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_974),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1013),
.A2(n_574),
.B(n_573),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1056),
.A2(n_758),
.B(n_695),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1106),
.A2(n_1034),
.B(n_1006),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1153),
.A2(n_570),
.B(n_563),
.Y(n_1217)
);

NOR2x1_ASAP7_75t_L g1218 ( 
.A(n_1010),
.B(n_417),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1089),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1010),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1013),
.A2(n_377),
.B(n_356),
.C(n_276),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1029),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_980),
.A2(n_393),
.B1(n_396),
.B2(n_398),
.C(n_401),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1000),
.B(n_277),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1125),
.B(n_908),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1153),
.A2(n_570),
.B(n_563),
.Y(n_1226)
);

AOI211x1_ASAP7_75t_L g1227 ( 
.A1(n_1036),
.A2(n_277),
.B(n_282),
.C(n_283),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1146),
.A2(n_573),
.A3(n_584),
.B(n_579),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1054),
.A2(n_756),
.B(n_746),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1059),
.A2(n_756),
.B(n_746),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1132),
.B(n_908),
.Y(n_1231)
);

NOR2x1_ASAP7_75t_SL g1232 ( 
.A(n_1142),
.B(n_1040),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1038),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1115),
.B(n_908),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1072),
.B(n_908),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1044),
.A2(n_570),
.B(n_563),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1037),
.B(n_908),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1041),
.B(n_908),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1078),
.A2(n_756),
.B(n_746),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_965),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_965),
.A2(n_584),
.A3(n_574),
.B(n_576),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_971),
.A2(n_584),
.A3(n_574),
.B(n_576),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_SL g1243 ( 
.A1(n_1109),
.A2(n_754),
.B(n_742),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_1040),
.A2(n_283),
.B(n_282),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1079),
.A2(n_577),
.B(n_570),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1052),
.Y(n_1246)
);

NOR2x1_ASAP7_75t_SL g1247 ( 
.A(n_1142),
.B(n_746),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1084),
.A2(n_758),
.B(n_695),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1093),
.A2(n_781),
.B(n_756),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1129),
.A2(n_577),
.B(n_578),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1053),
.B(n_402),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1002),
.B(n_756),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1038),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1038),
.B(n_1050),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1009),
.A2(n_379),
.B1(n_302),
.B2(n_312),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1011),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1077),
.A2(n_758),
.B(n_695),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_972),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1131),
.B(n_1096),
.C(n_1108),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1040),
.A2(n_312),
.B(n_302),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_972),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1134),
.A2(n_579),
.B(n_576),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1009),
.A2(n_362),
.B1(n_316),
.B2(n_327),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_966),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1100),
.A2(n_581),
.B(n_579),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_971),
.A2(n_577),
.B(n_578),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1071),
.B(n_404),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1090),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_SL g1270 ( 
.A1(n_1080),
.A2(n_1033),
.B(n_1123),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1139),
.B(n_316),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1095),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1062),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1141),
.A2(n_758),
.B(n_695),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_973),
.A2(n_577),
.B(n_578),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_986),
.B(n_409),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_973),
.A2(n_975),
.B(n_1027),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1149),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_975),
.A2(n_582),
.B(n_578),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1039),
.A2(n_357),
.B1(n_327),
.B2(n_331),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1049),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1130),
.A2(n_581),
.B(n_582),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1027),
.A2(n_1008),
.B(n_995),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_995),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1042),
.B(n_410),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1133),
.A2(n_758),
.B(n_695),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1042),
.B(n_412),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_987),
.B(n_781),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1122),
.A2(n_781),
.B(n_244),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1122),
.A2(n_781),
.B(n_245),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_969),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_979),
.B(n_422),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1140),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_983),
.B(n_428),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_994),
.B(n_430),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1101),
.A2(n_356),
.B(n_379),
.C(n_373),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_979),
.B(n_431),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1008),
.A2(n_582),
.B(n_581),
.Y(n_1299)
);

OAI22x1_ASAP7_75t_L g1300 ( 
.A1(n_1047),
.A2(n_424),
.B1(n_345),
.B2(n_419),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1144),
.A2(n_582),
.B(n_337),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_994),
.B(n_781),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1024),
.A2(n_337),
.B(n_331),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1024),
.A2(n_355),
.B(n_345),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_987),
.A2(n_250),
.B(n_243),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1149),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1089),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_979),
.B(n_355),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1025),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1025),
.A2(n_362),
.B(n_357),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1101),
.A2(n_424),
.B1(n_419),
.B2(n_418),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_964),
.B(n_369),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1152),
.A2(n_373),
.B(n_369),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_969),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1033),
.B(n_417),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_967),
.B(n_377),
.Y(n_1316)
);

NAND3x1_ASAP7_75t_L g1317 ( 
.A(n_1032),
.B(n_413),
.C(n_394),
.Y(n_1317)
);

AOI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1145),
.A2(n_413),
.B(n_394),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_992),
.B(n_1045),
.Y(n_1319)
);

O2A1O1Ixp5_ASAP7_75t_L g1320 ( 
.A1(n_1058),
.A2(n_418),
.B(n_754),
.C(n_742),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1075),
.B(n_1),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1028),
.A2(n_754),
.B(n_742),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1004),
.B(n_251),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1028),
.A2(n_754),
.A3(n_260),
.B(n_565),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1082),
.Y(n_1325)
);

BUFx10_ASAP7_75t_L g1326 ( 
.A(n_1325),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1245),
.A2(n_1236),
.B(n_1250),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1175),
.A2(n_1126),
.B1(n_1116),
.B2(n_1022),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1220),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1236),
.A2(n_1245),
.B(n_1163),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1240),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1211),
.A2(n_1123),
.B(n_1103),
.C(n_1154),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1173),
.B(n_1074),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_L g1334 ( 
.A(n_1279),
.B(n_1058),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1158),
.A2(n_1055),
.B(n_1031),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1311),
.A2(n_1085),
.B1(n_1050),
.B2(n_1047),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1271),
.A2(n_1223),
.B1(n_1102),
.B2(n_1091),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1240),
.Y(n_1338)
);

OAI221xp5_ASAP7_75t_L g1339 ( 
.A1(n_1295),
.A2(n_996),
.B1(n_1148),
.B2(n_1127),
.C(n_1085),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1285),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

AOI22x1_ASAP7_75t_L g1342 ( 
.A1(n_1159),
.A2(n_1066),
.B1(n_1098),
.B2(n_1124),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1309),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1177),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1250),
.A2(n_1055),
.B(n_1031),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1279),
.B(n_1080),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1279),
.B(n_1080),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1309),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1166),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1256),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1273),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1241),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1158),
.A2(n_1070),
.B(n_1061),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1203),
.B(n_1045),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1241),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1220),
.Y(n_1356)
);

AND2x4_ASAP7_75t_SL g1357 ( 
.A(n_1254),
.B(n_1045),
.Y(n_1357)
);

OAI222xp33_ASAP7_75t_L g1358 ( 
.A1(n_1162),
.A2(n_1021),
.B1(n_1085),
.B2(n_1050),
.C1(n_1063),
.C2(n_1032),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1296),
.A2(n_1102),
.B1(n_1091),
.B2(n_1021),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1177),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1241),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1202),
.B(n_1069),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1178),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1166),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1185),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1248),
.A2(n_1112),
.B(n_1118),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1254),
.B(n_1021),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1164),
.A2(n_1070),
.B(n_1061),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1296),
.A2(n_1111),
.B1(n_1082),
.B2(n_982),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1216),
.A2(n_993),
.B(n_987),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1198),
.A2(n_1087),
.B(n_1086),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1166),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1317),
.A2(n_1114),
.B1(n_1120),
.B2(n_1097),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1198),
.A2(n_1217),
.B(n_1209),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1211),
.B(n_1114),
.C(n_1082),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1209),
.A2(n_1087),
.B(n_1086),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1217),
.A2(n_1107),
.B(n_1099),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1166),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1226),
.A2(n_1107),
.B(n_1099),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1226),
.A2(n_1204),
.B(n_1267),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1204),
.A2(n_1137),
.B(n_1136),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1180),
.A2(n_1110),
.B1(n_1119),
.B2(n_1048),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1160),
.A2(n_1137),
.A3(n_1156),
.B(n_1136),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1297),
.A2(n_993),
.B(n_1048),
.C(n_1135),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1267),
.A2(n_1147),
.B(n_1143),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1185),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1319),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1185),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1275),
.A2(n_1147),
.B(n_1143),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1275),
.A2(n_1156),
.B(n_1150),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1282),
.B(n_1048),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1241),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1189),
.A2(n_1182),
.B1(n_1195),
.B2(n_1190),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1242),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1187),
.A2(n_1112),
.B(n_1157),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1306),
.B(n_1155),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1164),
.A2(n_1150),
.B(n_984),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1213),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1224),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_SL g1400 ( 
.A1(n_1297),
.A2(n_1066),
.B(n_1098),
.C(n_1005),
.Y(n_1400)
);

AO21x2_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_1221),
.B(n_1215),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1295),
.A2(n_1016),
.B1(n_984),
.B2(n_1157),
.C(n_1092),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1242),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1221),
.A2(n_1135),
.B(n_993),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1303),
.A2(n_1016),
.B(n_1155),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1306),
.B(n_1058),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1325),
.Y(n_1407)
);

OAI222xp33_ASAP7_75t_L g1408 ( 
.A1(n_1255),
.A2(n_1152),
.B1(n_1092),
.B2(n_1066),
.C1(n_1098),
.C2(n_1155),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1306),
.B(n_1065),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1292),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1165),
.A2(n_1065),
.B(n_1124),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1259),
.A2(n_1065),
.B(n_1124),
.C(n_1005),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1182),
.B(n_1069),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1165),
.A2(n_1014),
.B(n_1005),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1234),
.A2(n_1051),
.B(n_1030),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1242),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1314),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1254),
.B(n_1069),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1314),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1249),
.A2(n_1051),
.B(n_1030),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1201),
.A2(n_1152),
.B1(n_1081),
.B2(n_1073),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1242),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1278),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1188),
.B(n_1069),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1184),
.B(n_1073),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1276),
.A2(n_1014),
.B(n_4),
.C(n_5),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1287),
.A2(n_1172),
.B(n_1229),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1179),
.Y(n_1428)
);

OAI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1186),
.A2(n_1014),
.B1(n_254),
.B2(n_348),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1177),
.B(n_1030),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1252),
.B(n_1073),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1174),
.A2(n_352),
.B(n_257),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1289),
.A2(n_1051),
.B(n_1030),
.C(n_1081),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1235),
.A2(n_1051),
.B1(n_992),
.B2(n_1081),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1206),
.A2(n_336),
.B(n_269),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1179),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1181),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1168),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_SL g1439 ( 
.A1(n_1270),
.A2(n_1081),
.B(n_1073),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1194),
.B(n_992),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1179),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1179),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1183),
.A2(n_351),
.B(n_429),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1206),
.A2(n_1169),
.B(n_1322),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1169),
.A2(n_992),
.B(n_260),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1302),
.B(n_2),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1319),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1230),
.A2(n_315),
.B(n_323),
.Y(n_1448)
);

NOR2x1_ASAP7_75t_SL g1449 ( 
.A(n_1289),
.B(n_315),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1307),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1302),
.B(n_2),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1322),
.A2(n_260),
.B(n_389),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1192),
.B(n_1196),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1237),
.A2(n_315),
.B(n_323),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1170),
.A2(n_260),
.B(n_389),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1199),
.B(n_315),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1214),
.A2(n_260),
.B(n_315),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1257),
.A2(n_323),
.B(n_389),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1170),
.A2(n_389),
.B(n_323),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1265),
.B(n_425),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1197),
.B(n_4),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1253),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_R g1463 ( 
.A(n_1307),
.B(n_255),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1280),
.A2(n_389),
.B(n_323),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1280),
.A2(n_1193),
.B(n_1239),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1253),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1214),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1168),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_L g1469 ( 
.A(n_1262),
.B(n_102),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1212),
.B(n_5),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1193),
.A2(n_389),
.B(n_323),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1208),
.A2(n_212),
.B(n_211),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1222),
.B(n_6),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1208),
.A2(n_206),
.B(n_203),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1214),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1293),
.A2(n_7),
.B(n_12),
.C(n_15),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1238),
.A2(n_420),
.B1(n_411),
.B2(n_407),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1243),
.A2(n_197),
.B(n_193),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1231),
.A2(n_1176),
.B(n_1320),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1277),
.A2(n_188),
.B(n_184),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1228),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1210),
.A2(n_400),
.B(n_391),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1181),
.Y(n_1483)
);

CKINVDCx16_ASAP7_75t_R g1484 ( 
.A(n_1219),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1277),
.A2(n_176),
.B(n_175),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1318),
.A2(n_382),
.B(n_380),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1246),
.B(n_12),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1168),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1228),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1299),
.A2(n_364),
.B(n_359),
.Y(n_1490)
);

CKINVDCx14_ASAP7_75t_R g1491 ( 
.A(n_1219),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1260),
.B(n_15),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1317),
.A2(n_358),
.B1(n_343),
.B2(n_335),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1284),
.A2(n_173),
.B(n_166),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1228),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1225),
.A2(n_334),
.B(n_330),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1269),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1284),
.A2(n_164),
.B(n_162),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1299),
.A2(n_159),
.B(n_146),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1168),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1274),
.A2(n_322),
.B(n_319),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1272),
.B(n_16),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1171),
.Y(n_1503)
);

AOI21xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1300),
.A2(n_16),
.B(n_17),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1456),
.B(n_1315),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1370),
.A2(n_1202),
.B(n_1247),
.Y(n_1506)
);

AO31x2_ASAP7_75t_L g1507 ( 
.A1(n_1349),
.A2(n_1294),
.A3(n_1291),
.B(n_1290),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1357),
.B(n_1233),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1321),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1493),
.A2(n_1308),
.B(n_1304),
.C(n_1310),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1328),
.A2(n_1298),
.B1(n_1286),
.B2(n_1288),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1456),
.B(n_1315),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1359),
.A2(n_1227),
.B1(n_1264),
.B2(n_1312),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1497),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1337),
.A2(n_1336),
.B1(n_1493),
.B2(n_1375),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1331),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1350),
.B(n_1323),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1407),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1486),
.A2(n_1281),
.B1(n_1218),
.B2(n_1251),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1268),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1338),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1413),
.B(n_1252),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1484),
.B(n_1316),
.C(n_1305),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1365),
.B(n_1228),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1331),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1340),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1340),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1327),
.A2(n_1161),
.B(n_1263),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1336),
.A2(n_1233),
.B1(n_1313),
.B2(n_1167),
.Y(n_1529)
);

CKINVDCx6p67_ASAP7_75t_R g1530 ( 
.A(n_1407),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1329),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1363),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1329),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1504),
.A2(n_1301),
.B1(n_1207),
.B2(n_1262),
.C(n_1200),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1446),
.A2(n_1451),
.B1(n_1470),
.B2(n_1461),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1341),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1363),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1356),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1343),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1341),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1431),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1348),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1357),
.B(n_1171),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1348),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1327),
.A2(n_1266),
.B(n_1263),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1471),
.A2(n_1266),
.B(n_1263),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1356),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1396),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1395),
.A2(n_1486),
.B1(n_1502),
.B2(n_1492),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1437),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1487),
.A2(n_1200),
.B1(n_1266),
.B2(n_1191),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1486),
.A2(n_1261),
.B1(n_1244),
.B2(n_1283),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1437),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1504),
.A2(n_1258),
.B1(n_1171),
.B2(n_1205),
.Y(n_1555)
);

INVxp33_ASAP7_75t_L g1556 ( 
.A(n_1333),
.Y(n_1556)
);

NOR2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1450),
.B(n_1171),
.Y(n_1557)
);

AND2x6_ASAP7_75t_L g1558 ( 
.A(n_1437),
.B(n_1205),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1386),
.B(n_1205),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1450),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1456),
.A2(n_1369),
.B1(n_1398),
.B2(n_1339),
.Y(n_1561)
);

OAI222xp33_ASAP7_75t_L g1562 ( 
.A1(n_1373),
.A2(n_313),
.B1(n_300),
.B2(n_299),
.C1(n_297),
.C2(n_294),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1460),
.A2(n_1283),
.B1(n_1191),
.B2(n_1258),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1425),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1386),
.B(n_1205),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1453),
.A2(n_293),
.B1(n_1324),
.B2(n_24),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1481),
.A2(n_1232),
.B(n_1324),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1391),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1326),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1492),
.B(n_21),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1326),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1399),
.A2(n_1191),
.B1(n_1258),
.B2(n_1324),
.Y(n_1572)
);

AO21x2_ASAP7_75t_L g1573 ( 
.A1(n_1481),
.A2(n_1258),
.B(n_143),
.Y(n_1573)
);

CKINVDCx6p67_ASAP7_75t_R g1574 ( 
.A(n_1484),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1388),
.B(n_22),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1351),
.Y(n_1576)
);

CKINVDCx16_ASAP7_75t_R g1577 ( 
.A(n_1491),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1502),
.B(n_22),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1456),
.B(n_138),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1326),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1410),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1388),
.B(n_26),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1440),
.B(n_26),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1419),
.B(n_30),
.Y(n_1584)
);

CKINVDCx16_ASAP7_75t_R g1585 ( 
.A(n_1462),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1417),
.B(n_31),
.Y(n_1586)
);

INVx4_ASAP7_75t_SL g1587 ( 
.A(n_1437),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1423),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1462),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1396),
.B(n_1409),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1395),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1466),
.Y(n_1592)
);

BUFx4f_ASAP7_75t_SL g1593 ( 
.A(n_1466),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1354),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1393),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1384),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1467),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1424),
.B(n_48),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1476),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.C(n_53),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1427),
.A2(n_60),
.B(n_63),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1396),
.Y(n_1601)
);

NOR3xp33_ASAP7_75t_SL g1602 ( 
.A(n_1426),
.B(n_1358),
.C(n_1402),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1395),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1603)
);

INVx6_ASAP7_75t_L g1604 ( 
.A(n_1437),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1387),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1424),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1368),
.Y(n_1607)
);

NOR2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1418),
.B(n_64),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1396),
.B(n_66),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1382),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1373),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1429),
.A2(n_76),
.B1(n_77),
.B2(n_82),
.Y(n_1612)
);

NOR3xp33_ASAP7_75t_SL g1613 ( 
.A(n_1496),
.B(n_1477),
.C(n_1412),
.Y(n_1613)
);

OAI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1429),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1352),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1387),
.B(n_83),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1447),
.B(n_86),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1332),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.C(n_92),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1352),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_L g1620 ( 
.A(n_1443),
.B(n_90),
.C(n_93),
.D(n_94),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1409),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1409),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1409),
.B(n_95),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1355),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1367),
.B(n_96),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1355),
.Y(n_1626)
);

OR2x6_ASAP7_75t_SL g1627 ( 
.A(n_1418),
.B(n_96),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1367),
.B(n_97),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1404),
.A2(n_98),
.B1(n_104),
.B2(n_109),
.Y(n_1629)
);

INVx6_ASAP7_75t_L g1630 ( 
.A(n_1431),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_L g1631 ( 
.A(n_1439),
.B(n_110),
.Y(n_1631)
);

OR2x6_ASAP7_75t_L g1632 ( 
.A(n_1483),
.B(n_1447),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1483),
.B(n_111),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1432),
.A2(n_112),
.B1(n_123),
.B2(n_124),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1501),
.A2(n_125),
.B1(n_136),
.B2(n_1421),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1430),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1503),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1334),
.B(n_1503),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1362),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1334),
.B(n_1344),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1467),
.A2(n_1475),
.B1(n_1479),
.B2(n_1489),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1475),
.B(n_1344),
.Y(n_1642)
);

CKINVDCx16_ASAP7_75t_R g1643 ( 
.A(n_1463),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1361),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1482),
.A2(n_1400),
.B1(n_1489),
.B2(n_1495),
.C(n_1406),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1430),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1361),
.B(n_1392),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1392),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1430),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1394),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1394),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1406),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1406),
.B(n_1346),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1346),
.A2(n_1347),
.B1(n_1469),
.B2(n_1434),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1346),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1501),
.A2(n_1495),
.B1(n_1397),
.B2(n_1441),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1368),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1368),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1501),
.A2(n_1397),
.B1(n_1441),
.B2(n_1436),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1427),
.A2(n_1342),
.B(n_1420),
.Y(n_1660)
);

CKINVDCx14_ASAP7_75t_R g1661 ( 
.A(n_1463),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1347),
.A2(n_1469),
.B1(n_1416),
.B2(n_1422),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1433),
.A2(n_1454),
.B(n_1436),
.C(n_1442),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1428),
.A2(n_1442),
.B(n_1403),
.C(n_1422),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1408),
.A2(n_1401),
.B1(n_1416),
.B2(n_1403),
.C(n_1428),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1457),
.A2(n_1378),
.B(n_1349),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1342),
.A2(n_1347),
.B1(n_1490),
.B2(n_1435),
.C(n_1415),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1401),
.A2(n_1449),
.B1(n_1366),
.B2(n_1490),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1397),
.B(n_1344),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1360),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1360),
.B(n_1405),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1427),
.A2(n_1366),
.B(n_1458),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1368),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1381),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1494),
.A2(n_1498),
.B(n_1480),
.C(n_1485),
.Y(n_1675)
);

OAI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1490),
.A2(n_1435),
.B1(n_1448),
.B2(n_1360),
.C(n_1397),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1405),
.Y(n_1677)
);

CKINVDCx6p67_ASAP7_75t_R g1678 ( 
.A(n_1439),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1366),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1405),
.A2(n_1401),
.B1(n_1490),
.B2(n_1435),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1383),
.B(n_1500),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1335),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1411),
.B(n_1445),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1383),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1381),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1435),
.A2(n_1378),
.B1(n_1372),
.B2(n_1364),
.Y(n_1686)
);

CKINVDCx11_ASAP7_75t_R g1687 ( 
.A(n_1364),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1383),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1620),
.A2(n_1372),
.B1(n_1438),
.B2(n_1468),
.C(n_1488),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1515),
.A2(n_1458),
.B1(n_1468),
.B2(n_1488),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1611),
.A2(n_1438),
.B1(n_1335),
.B2(n_1457),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1509),
.B(n_1445),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1535),
.B(n_1480),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1535),
.A2(n_1458),
.B1(n_1330),
.B2(n_1383),
.C(n_1335),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1599),
.B(n_1335),
.C(n_1449),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1568),
.B(n_1371),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1599),
.A2(n_1498),
.B1(n_1494),
.B2(n_1485),
.C(n_1474),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1581),
.B(n_1411),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1594),
.A2(n_1371),
.B1(n_1345),
.B2(n_1390),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_R g1700 ( 
.A1(n_1627),
.A2(n_1499),
.B1(n_1474),
.B2(n_1472),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1596),
.A2(n_1330),
.B(n_1499),
.C(n_1472),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_SL g1702 ( 
.A(n_1618),
.B(n_1478),
.C(n_1471),
.D(n_1459),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1513),
.A2(n_1345),
.B1(n_1389),
.B2(n_1390),
.Y(n_1703)
);

INVxp33_ASAP7_75t_L g1704 ( 
.A(n_1517),
.Y(n_1704)
);

OAI332xp33_ASAP7_75t_L g1705 ( 
.A1(n_1595),
.A2(n_1455),
.A3(n_1459),
.B1(n_1353),
.B2(n_1330),
.B3(n_1465),
.C1(n_1379),
.C2(n_1377),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1510),
.A2(n_1414),
.B1(n_1478),
.B2(n_1380),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1514),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1561),
.A2(n_1389),
.B1(n_1385),
.B2(n_1376),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1602),
.A2(n_1414),
.B1(n_1380),
.B2(n_1353),
.Y(n_1709)
);

OAI222xp33_ASAP7_75t_L g1710 ( 
.A1(n_1549),
.A2(n_1455),
.B1(n_1385),
.B2(n_1377),
.C1(n_1379),
.C2(n_1376),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1513),
.A2(n_1444),
.B1(n_1465),
.B2(n_1464),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1588),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1618),
.A2(n_1444),
.B1(n_1464),
.B2(n_1452),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1614),
.A2(n_1610),
.B1(n_1595),
.B2(n_1600),
.C(n_1612),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1600),
.A2(n_1374),
.B(n_1452),
.C(n_1591),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1596),
.A2(n_1374),
.B1(n_1610),
.B2(n_1579),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1532),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1576),
.B(n_1520),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1602),
.A2(n_1603),
.B1(n_1613),
.B2(n_1523),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_SL g1720 ( 
.A(n_1632),
.B(n_1579),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1577),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1561),
.A2(n_1608),
.B1(n_1511),
.B2(n_1634),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1613),
.A2(n_1634),
.B(n_1562),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1523),
.A2(n_1609),
.B1(n_1623),
.B2(n_1629),
.Y(n_1724)
);

OAI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1579),
.A2(n_1582),
.B1(n_1556),
.B2(n_1585),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_SL g1726 ( 
.A1(n_1566),
.A2(n_1578),
.B1(n_1570),
.B2(n_1679),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1531),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1609),
.A2(n_1639),
.B1(n_1643),
.B2(n_1529),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1547),
.B(n_1590),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1549),
.B(n_1519),
.C(n_1680),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1562),
.A2(n_1641),
.B1(n_1676),
.B2(n_1564),
.C(n_1555),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1635),
.A2(n_1661),
.B1(n_1524),
.B2(n_1628),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1623),
.A2(n_1593),
.B1(n_1574),
.B2(n_1575),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1625),
.A2(n_1584),
.B1(n_1583),
.B2(n_1668),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1516),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1575),
.A2(n_1592),
.B1(n_1589),
.B2(n_1580),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1605),
.A2(n_1598),
.B1(n_1534),
.B2(n_1557),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1668),
.B(n_1563),
.C(n_1676),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1606),
.A2(n_1665),
.B1(n_1537),
.B2(n_1586),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_SL g1740 ( 
.A1(n_1573),
.A2(n_1633),
.B1(n_1667),
.B2(n_1551),
.Y(n_1740)
);

INVxp33_ASAP7_75t_L g1741 ( 
.A(n_1531),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1590),
.B(n_1533),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1597),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1548),
.B(n_1601),
.Y(n_1744)
);

BUFx4f_ASAP7_75t_SL g1745 ( 
.A(n_1530),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1641),
.A2(n_1665),
.B1(n_1551),
.B2(n_1667),
.C(n_1645),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1534),
.A2(n_1622),
.B1(n_1637),
.B2(n_1571),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1525),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1538),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1506),
.A2(n_1660),
.B(n_1675),
.Y(n_1750)
);

AOI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1541),
.A2(n_1527),
.B1(n_1542),
.B2(n_1536),
.C1(n_1544),
.C2(n_1526),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1645),
.A2(n_1522),
.B1(n_1672),
.B2(n_1656),
.C(n_1626),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1573),
.A2(n_1633),
.B1(n_1684),
.B2(n_1505),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1505),
.B(n_1512),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1522),
.A2(n_1505),
.B1(n_1512),
.B2(n_1518),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1541),
.B(n_1552),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1548),
.B(n_1601),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1537),
.A2(n_1687),
.B1(n_1659),
.B2(n_1512),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1537),
.A2(n_1630),
.B1(n_1617),
.B2(n_1616),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1672),
.A2(n_1650),
.B1(n_1648),
.B2(n_1619),
.C(n_1644),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1622),
.A2(n_1571),
.B1(n_1553),
.B2(n_1621),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1569),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1540),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1615),
.A2(n_1624),
.B1(n_1651),
.B2(n_1664),
.C(n_1688),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1663),
.A2(n_1572),
.B1(n_1518),
.B2(n_1631),
.C(n_1565),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1538),
.Y(n_1766)
);

OAI211xp5_ASAP7_75t_L g1767 ( 
.A1(n_1660),
.A2(n_1642),
.B(n_1597),
.C(n_1559),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1647),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1630),
.A2(n_1662),
.B1(n_1508),
.B2(n_1538),
.Y(n_1769)
);

INVx5_ASAP7_75t_SL g1770 ( 
.A(n_1632),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1642),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1559),
.B(n_1565),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1521),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1653),
.B(n_1587),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1539),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1669),
.B(n_1671),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1652),
.A2(n_1655),
.B1(n_1649),
.B2(n_1654),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1587),
.B(n_1543),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1640),
.B(n_1638),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1640),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1673),
.A2(n_1682),
.B1(n_1686),
.B2(n_1681),
.C(n_1677),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1550),
.B(n_1604),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1655),
.A2(n_1649),
.B1(n_1560),
.B2(n_1678),
.Y(n_1783)
);

AOI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1682),
.A2(n_1681),
.B1(n_1607),
.B2(n_1658),
.C(n_1657),
.Y(n_1784)
);

AOI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1674),
.A2(n_1685),
.B1(n_1646),
.B2(n_1636),
.C(n_1683),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1550),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1554),
.A2(n_1604),
.B1(n_1558),
.B2(n_1567),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1636),
.A2(n_1646),
.B1(n_1506),
.B2(n_1554),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1558),
.A2(n_1567),
.B1(n_1666),
.B2(n_1587),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1670),
.A2(n_1528),
.B(n_1545),
.C(n_1507),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1670),
.B(n_1558),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1683),
.A2(n_1558),
.B1(n_1507),
.B2(n_1546),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1666),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1507),
.A2(n_970),
.B(n_1506),
.Y(n_1794)
);

BUFx8_ASAP7_75t_SL g1795 ( 
.A(n_1532),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1581),
.B(n_858),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1660),
.A2(n_1327),
.B(n_1545),
.Y(n_1797)
);

NOR2x1_ASAP7_75t_SL g1798 ( 
.A(n_1632),
.B(n_1579),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1589),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1535),
.A2(n_751),
.B1(n_804),
.B2(n_802),
.C(n_1504),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1802)
);

OAI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1515),
.A2(n_1620),
.B1(n_1611),
.B2(n_1336),
.Y(n_1803)
);

AOI21xp33_ASAP7_75t_L g1804 ( 
.A1(n_1535),
.A2(n_804),
.B(n_802),
.Y(n_1804)
);

AOI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1535),
.A2(n_804),
.B(n_802),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1589),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1515),
.A2(n_970),
.B1(n_804),
.B2(n_802),
.Y(n_1808)
);

OAI222xp33_ASAP7_75t_L g1809 ( 
.A1(n_1515),
.A2(n_1611),
.B1(n_1336),
.B2(n_1549),
.C1(n_1493),
.C2(n_1596),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1514),
.B(n_1606),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_713),
.B2(n_688),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1600),
.A2(n_1535),
.B(n_1457),
.Y(n_1812)
);

AO221x1_ASAP7_75t_L g1813 ( 
.A1(n_1629),
.A2(n_1596),
.B1(n_1595),
.B2(n_1594),
.C(n_1614),
.Y(n_1813)
);

OAI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1620),
.A2(n_802),
.B1(n_804),
.B2(n_1295),
.C(n_1337),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1620),
.A2(n_802),
.B(n_804),
.C(n_1599),
.Y(n_1815)
);

INVx5_ASAP7_75t_SL g1816 ( 
.A(n_1530),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1576),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1599),
.B(n_804),
.C(n_802),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1660),
.A2(n_1672),
.B(n_1675),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1620),
.A2(n_802),
.B1(n_804),
.B2(n_1295),
.C(n_1337),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1514),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1594),
.A2(n_980),
.B1(n_1358),
.B2(n_548),
.C1(n_1328),
.C2(n_1599),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1514),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1514),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1597),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1561),
.A2(n_451),
.B1(n_452),
.B2(n_447),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1509),
.B(n_1547),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1514),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_L g1834 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1561),
.A2(n_451),
.B1(n_452),
.B2(n_447),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1514),
.Y(n_1838)
);

BUFx12f_ASAP7_75t_L g1839 ( 
.A(n_1532),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1620),
.A2(n_923),
.B1(n_1594),
.B2(n_804),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1509),
.B(n_1547),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1568),
.B(n_1497),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_SL g1843 ( 
.A1(n_1561),
.A2(n_451),
.B1(n_452),
.B2(n_447),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1506),
.A2(n_970),
.B(n_1456),
.Y(n_1844)
);

OA21x2_ASAP7_75t_L g1845 ( 
.A1(n_1660),
.A2(n_1672),
.B(n_1675),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1509),
.B(n_1547),
.Y(n_1846)
);

OAI222xp33_ASAP7_75t_L g1847 ( 
.A1(n_1515),
.A2(n_1611),
.B1(n_1336),
.B2(n_1549),
.C1(n_1493),
.C2(n_1596),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1547),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1509),
.B(n_1547),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1743),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1776),
.B(n_1720),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1743),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1793),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1771),
.B(n_1826),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1798),
.B(n_1791),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1692),
.B(n_1830),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1773),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1744),
.B(n_1757),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1826),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1848),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1754),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1819),
.B(n_1829),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1841),
.B(n_1846),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1754),
.B(n_1738),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1756),
.B(n_1772),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1735),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1849),
.B(n_1748),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1808),
.A2(n_1823),
.B1(n_1803),
.B2(n_1818),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1707),
.B(n_1822),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1833),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1763),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1768),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1775),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1795),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_SL g1875 ( 
.A(n_1723),
.B(n_1809),
.Y(n_1875)
);

AOI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1813),
.A2(n_1835),
.B1(n_1843),
.B2(n_1828),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1810),
.B(n_1824),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1825),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1780),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1831),
.B(n_1838),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1696),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1712),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1837),
.B(n_1842),
.Y(n_1883)
);

OAI321xp33_ASAP7_75t_L g1884 ( 
.A1(n_1719),
.A2(n_1815),
.A3(n_1803),
.B1(n_1722),
.B2(n_1800),
.C(n_1814),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1751),
.B(n_1698),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1714),
.A2(n_1801),
.B1(n_1840),
.B2(n_1802),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1774),
.B(n_1787),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1729),
.B(n_1746),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1693),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1801),
.A2(n_1802),
.B1(n_1840),
.B2(n_1827),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1796),
.B(n_1799),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1778),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1760),
.B(n_1794),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1806),
.A2(n_1827),
.B1(n_1836),
.B2(n_1832),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1820),
.B(n_1845),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1785),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1820),
.B(n_1845),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1820),
.B(n_1845),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1718),
.B(n_1742),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1817),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1792),
.Y(n_1901)
);

AOI322xp5_ASAP7_75t_L g1902 ( 
.A1(n_1806),
.A2(n_1832),
.A3(n_1836),
.B1(n_1834),
.B2(n_1811),
.C1(n_1805),
.C2(n_1804),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1797),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1767),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1752),
.B(n_1784),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1749),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1812),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1689),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1774),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1779),
.B(n_1730),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1703),
.B(n_1694),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1764),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1739),
.B(n_1770),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1703),
.B(n_1740),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1787),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1708),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1781),
.B(n_1750),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1731),
.B(n_1844),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1690),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1709),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1711),
.B(n_1699),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1711),
.B(n_1699),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1706),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1789),
.B(n_1782),
.Y(n_1924)
);

CKINVDCx6p67_ASAP7_75t_R g1925 ( 
.A(n_1762),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1788),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1788),
.B(n_1716),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1727),
.B(n_1734),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1716),
.B(n_1725),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1790),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1792),
.Y(n_1931)
);

INVxp67_ASAP7_75t_SL g1932 ( 
.A(n_1701),
.Y(n_1932)
);

NAND2x1_ASAP7_75t_L g1933 ( 
.A(n_1761),
.B(n_1747),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1734),
.B(n_1759),
.Y(n_1934)
);

AO21x2_ASAP7_75t_L g1935 ( 
.A1(n_1691),
.A2(n_1710),
.B(n_1695),
.Y(n_1935)
);

INVx4_ASAP7_75t_L g1936 ( 
.A(n_1786),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1766),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1759),
.B(n_1736),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1758),
.B(n_1713),
.Y(n_1940)
);

BUFx2_ASAP7_75t_L g1941 ( 
.A(n_1783),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1755),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_SL g1943 ( 
.A(n_1875),
.B(n_1721),
.Y(n_1943)
);

AOI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1884),
.A2(n_1821),
.B(n_1847),
.C(n_1724),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1868),
.B(n_1834),
.C(n_1726),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1924),
.B(n_1737),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1850),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1875),
.A2(n_1732),
.B1(n_1753),
.B2(n_1700),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1859),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1853),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1852),
.Y(n_1951)
);

OAI31xp33_ASAP7_75t_L g1952 ( 
.A1(n_1894),
.A2(n_1715),
.A3(n_1732),
.B(n_1777),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1874),
.Y(n_1953)
);

CKINVDCx8_ASAP7_75t_R g1954 ( 
.A(n_1941),
.Y(n_1954)
);

OAI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1868),
.A2(n_1939),
.B1(n_1894),
.B2(n_1929),
.Y(n_1955)
);

AOI31xp33_ASAP7_75t_L g1956 ( 
.A1(n_1939),
.A2(n_1733),
.A3(n_1783),
.B(n_1728),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1925),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1856),
.B(n_1758),
.Y(n_1958)
);

AOI33xp33_ASAP7_75t_L g1959 ( 
.A1(n_1886),
.A2(n_1713),
.A3(n_1691),
.B1(n_1777),
.B2(n_1769),
.B3(n_1704),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1870),
.B(n_1741),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1855),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1852),
.Y(n_1962)
);

AO21x2_ASAP7_75t_L g1963 ( 
.A1(n_1907),
.A2(n_1697),
.B(n_1765),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1855),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1853),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1866),
.Y(n_1966)
);

OAI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1890),
.A2(n_1769),
.B1(n_1807),
.B2(n_1717),
.C(n_1702),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1856),
.B(n_1816),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1884),
.A2(n_1745),
.B(n_1816),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1866),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1865),
.B(n_1816),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1879),
.Y(n_1972)
);

AOI211xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1932),
.A2(n_1745),
.B(n_1839),
.C(n_1929),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1904),
.B(n_1902),
.C(n_1917),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1858),
.B(n_1901),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1862),
.B(n_1883),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1854),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_L g1978 ( 
.A(n_1904),
.B(n_1902),
.C(n_1917),
.Y(n_1978)
);

NOR3xp33_ASAP7_75t_SL g1979 ( 
.A(n_1930),
.B(n_1932),
.C(n_1891),
.Y(n_1979)
);

OAI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1885),
.A2(n_1918),
.B1(n_1896),
.B2(n_1905),
.Y(n_1980)
);

INVxp67_ASAP7_75t_L g1981 ( 
.A(n_1937),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1858),
.B(n_1901),
.Y(n_1982)
);

OAI222xp33_ASAP7_75t_L g1983 ( 
.A1(n_1885),
.A2(n_1905),
.B1(n_1914),
.B2(n_1934),
.C1(n_1896),
.C2(n_1876),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1909),
.B(n_1887),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1858),
.B(n_1867),
.Y(n_1985)
);

NAND4xp25_ASAP7_75t_L g1986 ( 
.A(n_1930),
.B(n_1922),
.C(n_1921),
.D(n_1920),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1914),
.A2(n_1908),
.B1(n_1934),
.B2(n_1919),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1862),
.B(n_1883),
.Y(n_1988)
);

OAI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1907),
.A2(n_1903),
.B(n_1920),
.Y(n_1989)
);

AOI221x1_ASAP7_75t_L g1990 ( 
.A1(n_1912),
.A2(n_1908),
.B1(n_1918),
.B2(n_1915),
.C(n_1919),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1865),
.B(n_1877),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1854),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1921),
.A2(n_1922),
.B1(n_1912),
.B2(n_1911),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1877),
.B(n_1860),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1878),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1858),
.B(n_1867),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1927),
.A2(n_1864),
.B1(n_1941),
.B2(n_1913),
.Y(n_1997)
);

AOI21xp33_ASAP7_75t_L g1998 ( 
.A1(n_1935),
.A2(n_1893),
.B(n_1911),
.Y(n_1998)
);

INVx5_ASAP7_75t_L g1999 ( 
.A(n_1864),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1940),
.A2(n_1910),
.B1(n_1935),
.B2(n_1915),
.Y(n_2000)
);

OAI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1927),
.A2(n_1893),
.B(n_1889),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1863),
.B(n_1931),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1935),
.A2(n_1933),
.B(n_1923),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1860),
.B(n_1872),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1863),
.B(n_1931),
.Y(n_2005)
);

AOI33xp33_ASAP7_75t_L g2006 ( 
.A1(n_1888),
.A2(n_1938),
.A3(n_1940),
.B1(n_1895),
.B2(n_1897),
.B3(n_1898),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1879),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_R g2008 ( 
.A(n_1925),
.B(n_1909),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_L g2009 ( 
.A(n_1920),
.B(n_1926),
.C(n_1923),
.Y(n_2009)
);

INVxp67_ASAP7_75t_SL g2010 ( 
.A(n_1895),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1888),
.A2(n_1935),
.B1(n_1864),
.B2(n_1938),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1860),
.B(n_1869),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1950),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1991),
.B(n_1916),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_2010),
.B(n_1897),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1947),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1975),
.B(n_1898),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1977),
.B(n_1881),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1962),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1975),
.B(n_1899),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1977),
.B(n_1881),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1953),
.B(n_1925),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1962),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1982),
.B(n_1899),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1953),
.B(n_1936),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1982),
.B(n_1923),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1947),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_2008),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1984),
.B(n_1892),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_1974),
.A2(n_1872),
.B1(n_1926),
.B2(n_1882),
.C(n_1878),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1985),
.B(n_1996),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1965),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1992),
.B(n_1882),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1992),
.B(n_2006),
.Y(n_2034)
);

NAND2x1p5_ASAP7_75t_L g2035 ( 
.A(n_1999),
.B(n_1933),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1994),
.B(n_1880),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2003),
.B(n_1906),
.Y(n_2037)
);

NAND2x1p5_ASAP7_75t_L g2038 ( 
.A(n_1999),
.B(n_1861),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1976),
.B(n_1871),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2002),
.B(n_1900),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1966),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1988),
.B(n_1871),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1951),
.B(n_1910),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2005),
.B(n_1909),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1971),
.B(n_1936),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1966),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1971),
.B(n_1936),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1970),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1970),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2012),
.B(n_1851),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1995),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1949),
.B(n_1857),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1998),
.B(n_1873),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1957),
.B(n_1936),
.Y(n_2054)
);

AND2x2_ASAP7_75t_SL g2055 ( 
.A(n_2011),
.B(n_1887),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_2004),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1989),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1958),
.B(n_1887),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1995),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1989),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_2004),
.B(n_1942),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_1961),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1957),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_2034),
.B(n_2009),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2057),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2017),
.B(n_1972),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2017),
.B(n_1972),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2057),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_2035),
.B(n_1954),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2057),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2034),
.B(n_2043),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2017),
.B(n_2007),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2041),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_2055),
.A2(n_2000),
.B1(n_1948),
.B2(n_1974),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2041),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2043),
.B(n_2001),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2015),
.B(n_2007),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2019),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2060),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2015),
.B(n_1958),
.Y(n_2080)
);

BUFx3_ASAP7_75t_L g2081 ( 
.A(n_2063),
.Y(n_2081)
);

OAI21xp33_ASAP7_75t_SL g2082 ( 
.A1(n_2055),
.A2(n_2030),
.B(n_2015),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2046),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2016),
.B(n_1978),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2060),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2046),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2016),
.B(n_1978),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2027),
.B(n_1955),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2048),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2060),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2035),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_2061),
.B(n_1986),
.Y(n_2093)
);

NOR2x1p5_ASAP7_75t_SL g2094 ( 
.A(n_2027),
.B(n_1903),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2049),
.Y(n_2095)
);

AOI21xp33_ASAP7_75t_SL g2096 ( 
.A1(n_2035),
.A2(n_1969),
.B(n_1980),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2049),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2031),
.B(n_1961),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2051),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2013),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2035),
.A2(n_1952),
.B(n_1944),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2018),
.B(n_2021),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2059),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2018),
.B(n_2011),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2021),
.B(n_1981),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2013),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2059),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_2037),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2030),
.B(n_2033),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2033),
.B(n_1979),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2061),
.B(n_1960),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2039),
.B(n_1993),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2031),
.B(n_1964),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2052),
.Y(n_2114)
);

OAI21xp33_ASAP7_75t_L g2115 ( 
.A1(n_2037),
.A2(n_1944),
.B(n_1945),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2109),
.B(n_2056),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2100),
.Y(n_2117)
);

NOR2x1_ASAP7_75t_R g2118 ( 
.A(n_2081),
.B(n_2028),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2100),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2064),
.B(n_2036),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2100),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_2115),
.A2(n_2055),
.B1(n_1945),
.B2(n_1943),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2073),
.Y(n_2123)
);

AND2x2_ASAP7_75t_SL g2124 ( 
.A(n_2064),
.B(n_2028),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_L g2125 ( 
.A(n_2115),
.B(n_2022),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2109),
.B(n_2056),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2080),
.B(n_2031),
.Y(n_2127)
);

NAND2xp33_ASAP7_75t_R g2128 ( 
.A(n_2101),
.B(n_2058),
.Y(n_2128)
);

INVxp67_ASAP7_75t_SL g2129 ( 
.A(n_2084),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2080),
.B(n_2020),
.Y(n_2130)
);

NOR4xp25_ASAP7_75t_SL g2131 ( 
.A(n_2096),
.B(n_1967),
.C(n_1973),
.D(n_1956),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2073),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2064),
.B(n_2036),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_L g2134 ( 
.A(n_2082),
.B(n_1990),
.C(n_1987),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2075),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2106),
.A2(n_2053),
.B(n_2032),
.Y(n_2136)
);

AOI211xp5_ASAP7_75t_L g2137 ( 
.A1(n_2082),
.A2(n_2101),
.B(n_2096),
.C(n_1983),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2080),
.B(n_2062),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2098),
.B(n_2020),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2075),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2141)
);

NAND2xp33_ASAP7_75t_R g2142 ( 
.A(n_2092),
.B(n_2058),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2083),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_2081),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_2092),
.B(n_2029),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2083),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2084),
.B(n_2052),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2113),
.B(n_2024),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2087),
.B(n_2039),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2086),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2087),
.B(n_2042),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2086),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2113),
.B(n_2024),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2113),
.B(n_2050),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2071),
.B(n_2042),
.Y(n_2156)
);

NAND2xp33_ASAP7_75t_L g2157 ( 
.A(n_2110),
.B(n_2069),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2066),
.B(n_2026),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2071),
.B(n_2026),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2066),
.B(n_2026),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2089),
.Y(n_2161)
);

INVx4_ASAP7_75t_L g2162 ( 
.A(n_2081),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2066),
.B(n_2044),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2067),
.B(n_2044),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2129),
.B(n_2088),
.Y(n_2165)
);

OAI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2137),
.A2(n_2088),
.B(n_2074),
.Y(n_2166)
);

OAI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_2134),
.A2(n_1954),
.B1(n_1990),
.B2(n_2093),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2123),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_2144),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2125),
.B(n_2076),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2129),
.B(n_2076),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_2137),
.B(n_2110),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_2118),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2123),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2124),
.B(n_2093),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2124),
.B(n_2108),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2120),
.B(n_2105),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2132),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_L g2179 ( 
.A1(n_2134),
.A2(n_2094),
.B(n_2104),
.C(n_2112),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2120),
.B(n_2105),
.Y(n_2180)
);

AOI321xp33_ASAP7_75t_L g2181 ( 
.A1(n_2122),
.A2(n_2116),
.A3(n_2126),
.B1(n_2104),
.B2(n_2128),
.C(n_2152),
.Y(n_2181)
);

AO21x1_ASAP7_75t_L g2182 ( 
.A1(n_2116),
.A2(n_2112),
.B(n_2102),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_2124),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_SL g2184 ( 
.A1(n_2126),
.A2(n_2108),
.B(n_2077),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2132),
.Y(n_2185)
);

OAI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_2157),
.A2(n_2078),
.B(n_2077),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2127),
.Y(n_2187)
);

CKINVDCx16_ASAP7_75t_R g2188 ( 
.A(n_2131),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2135),
.Y(n_2189)
);

AOI21xp33_ASAP7_75t_L g2190 ( 
.A1(n_2148),
.A2(n_2118),
.B(n_2150),
.Y(n_2190)
);

AOI31xp33_ASAP7_75t_L g2191 ( 
.A1(n_2144),
.A2(n_2025),
.A3(n_2078),
.B(n_2054),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2142),
.A2(n_1946),
.B1(n_1997),
.B2(n_2058),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2150),
.A2(n_1946),
.B1(n_1928),
.B2(n_1963),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2133),
.B(n_2156),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2135),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2131),
.A2(n_2102),
.B(n_2053),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2152),
.B(n_2114),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2156),
.B(n_2114),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2140),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2140),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2130),
.B(n_2040),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2127),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2133),
.B(n_2111),
.Y(n_2203)
);

OAI221xp5_ASAP7_75t_SL g2204 ( 
.A1(n_2181),
.A2(n_2148),
.B1(n_2159),
.B2(n_1959),
.C(n_2127),
.Y(n_2204)
);

AOI22x1_ASAP7_75t_L g2205 ( 
.A1(n_2188),
.A2(n_2162),
.B1(n_2138),
.B2(n_2145),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2168),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2174),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2170),
.B(n_2130),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2178),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2187),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2170),
.A2(n_2179),
.B1(n_2167),
.B2(n_2172),
.Y(n_2211)
);

NAND2x1_ASAP7_75t_L g2212 ( 
.A(n_2191),
.B(n_2162),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2172),
.B(n_2158),
.Y(n_2213)
);

O2A1O1Ixp5_ASAP7_75t_L g2214 ( 
.A1(n_2182),
.A2(n_2162),
.B(n_2153),
.C(n_2143),
.Y(n_2214)
);

OAI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2179),
.A2(n_2159),
.B1(n_2117),
.B2(n_2119),
.C(n_2121),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2165),
.B(n_2169),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2167),
.A2(n_2162),
.B(n_2147),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2186),
.A2(n_2158),
.B1(n_2160),
.B2(n_2145),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2169),
.B(n_2158),
.Y(n_2219)
);

NOR2x1_ASAP7_75t_L g2220 ( 
.A(n_2183),
.B(n_2063),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2171),
.B(n_2160),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2173),
.B(n_2138),
.Y(n_2222)
);

OAI31xp33_ASAP7_75t_L g2223 ( 
.A1(n_2184),
.A2(n_2138),
.A3(n_2119),
.B(n_2121),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2185),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2187),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2189),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2195),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2199),
.Y(n_2228)
);

AOI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2166),
.A2(n_2196),
.B1(n_2175),
.B2(n_2193),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2192),
.A2(n_2117),
.B1(n_2121),
.B2(n_2119),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2176),
.A2(n_2117),
.B1(n_1963),
.B2(n_1946),
.Y(n_2231)
);

A2O1A1Ixp33_ASAP7_75t_L g2232 ( 
.A1(n_2190),
.A2(n_2094),
.B(n_2136),
.C(n_2160),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2214),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2211),
.B(n_2194),
.Y(n_2234)
);

NAND4xp25_ASAP7_75t_L g2235 ( 
.A(n_2222),
.B(n_2202),
.C(n_2200),
.D(n_2177),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2208),
.B(n_2213),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2210),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2210),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2225),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2220),
.B(n_2202),
.Y(n_2240)
);

INVxp67_ASAP7_75t_SL g2241 ( 
.A(n_2212),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2219),
.B(n_2203),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2225),
.B(n_2216),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2215),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_2212),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2206),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_2222),
.B(n_2180),
.Y(n_2247)
);

AOI221x1_ASAP7_75t_L g2248 ( 
.A1(n_2217),
.A2(n_2197),
.B1(n_2198),
.B2(n_2143),
.C(n_2147),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2207),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_R g2250 ( 
.A(n_2209),
.B(n_2063),
.Y(n_2250)
);

NOR2xp67_ASAP7_75t_SL g2251 ( 
.A(n_2224),
.B(n_2226),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_2205),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2229),
.B(n_2201),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2227),
.Y(n_2254)
);

NOR4xp25_ASAP7_75t_SL g2255 ( 
.A(n_2204),
.B(n_2161),
.C(n_2153),
.D(n_2151),
.Y(n_2255)
);

O2A1O1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_2232),
.A2(n_2161),
.B(n_2151),
.C(n_2023),
.Y(n_2256)
);

INVxp67_ASAP7_75t_L g2257 ( 
.A(n_2251),
.Y(n_2257)
);

OAI221xp5_ASAP7_75t_L g2258 ( 
.A1(n_2233),
.A2(n_2229),
.B1(n_2232),
.B2(n_2223),
.C(n_2231),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2247),
.B(n_2221),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2251),
.B(n_2228),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2237),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2234),
.B(n_2139),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2252),
.B(n_2218),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2255),
.B(n_2139),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2233),
.B(n_2149),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2242),
.B(n_2253),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2236),
.B(n_2149),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2248),
.B(n_2154),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_2248),
.A2(n_2230),
.B(n_2145),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2235),
.B(n_2145),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2250),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2261),
.Y(n_2272)
);

O2A1O1Ixp33_ASAP7_75t_L g2273 ( 
.A1(n_2258),
.A2(n_2257),
.B(n_2266),
.C(n_2244),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_R g2274 ( 
.A(n_2271),
.B(n_2252),
.Y(n_2274)
);

OAI211xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2263),
.A2(n_2256),
.B(n_2243),
.C(n_2241),
.Y(n_2275)
);

A2O1A1Ixp33_ASAP7_75t_L g2276 ( 
.A1(n_2269),
.A2(n_2244),
.B(n_2237),
.C(n_2239),
.Y(n_2276)
);

AOI211xp5_ASAP7_75t_L g2277 ( 
.A1(n_2268),
.A2(n_2240),
.B(n_2245),
.C(n_2254),
.Y(n_2277)
);

NOR4xp75_ASAP7_75t_L g2278 ( 
.A(n_2265),
.B(n_2264),
.C(n_2259),
.D(n_2262),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2260),
.B(n_2245),
.Y(n_2279)
);

NAND5xp2_ASAP7_75t_L g2280 ( 
.A(n_2270),
.B(n_2240),
.C(n_2249),
.D(n_2246),
.E(n_2238),
.Y(n_2280)
);

OAI211xp5_ASAP7_75t_SL g2281 ( 
.A1(n_2270),
.A2(n_2245),
.B(n_2254),
.C(n_2246),
.Y(n_2281)
);

AOI221x1_ASAP7_75t_L g2282 ( 
.A1(n_2267),
.A2(n_2239),
.B1(n_2238),
.B2(n_2249),
.C(n_2070),
.Y(n_2282)
);

AOI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2258),
.A2(n_2090),
.B1(n_2065),
.B2(n_2068),
.C(n_2070),
.Y(n_2283)
);

AOI211xp5_ASAP7_75t_L g2284 ( 
.A1(n_2258),
.A2(n_2146),
.B(n_2141),
.C(n_2136),
.Y(n_2284)
);

AOI221xp5_ASAP7_75t_L g2285 ( 
.A1(n_2258),
.A2(n_2090),
.B1(n_2065),
.B2(n_2068),
.C(n_2070),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2277),
.B(n_2163),
.Y(n_2286)
);

XNOR2xp5_ASAP7_75t_L g2287 ( 
.A(n_2278),
.B(n_2038),
.Y(n_2287)
);

XNOR2xp5_ASAP7_75t_L g2288 ( 
.A(n_2284),
.B(n_2038),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2276),
.A2(n_2090),
.B1(n_2085),
.B2(n_2079),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_R g2290 ( 
.A(n_2272),
.B(n_2045),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2274),
.B(n_2275),
.Y(n_2291)
);

XOR2xp5_ASAP7_75t_L g2292 ( 
.A(n_2279),
.B(n_2111),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2273),
.B(n_2163),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_R g2294 ( 
.A(n_2280),
.B(n_2047),
.Y(n_2294)
);

A2O1A1Ixp33_ASAP7_75t_SL g2295 ( 
.A1(n_2286),
.A2(n_2281),
.B(n_2282),
.C(n_2283),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2291),
.B(n_2292),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_2293),
.B(n_2141),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2287),
.B(n_2285),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_2290),
.Y(n_2299)
);

OAI211xp5_ASAP7_75t_SL g2300 ( 
.A1(n_2294),
.A2(n_2097),
.B(n_2095),
.C(n_2091),
.Y(n_2300)
);

NOR2x1p5_ASAP7_75t_L g2301 ( 
.A(n_2288),
.B(n_2141),
.Y(n_2301)
);

NOR3xp33_ASAP7_75t_L g2302 ( 
.A(n_2289),
.B(n_2136),
.C(n_2085),
.Y(n_2302)
);

NAND5xp2_ASAP7_75t_L g2303 ( 
.A(n_2296),
.B(n_2298),
.C(n_2302),
.D(n_2295),
.E(n_2301),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2299),
.B(n_2163),
.Y(n_2304)
);

O2A1O1Ixp33_ASAP7_75t_L g2305 ( 
.A1(n_2300),
.A2(n_2079),
.B(n_2085),
.C(n_2065),
.Y(n_2305)
);

NOR2x1p5_ASAP7_75t_L g2306 ( 
.A(n_2297),
.B(n_2146),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2295),
.A2(n_2146),
.B(n_2164),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_SL g2308 ( 
.A(n_2296),
.B(n_2154),
.C(n_2164),
.Y(n_2308)
);

NAND4xp25_ASAP7_75t_SL g2309 ( 
.A(n_2298),
.B(n_2164),
.C(n_2077),
.D(n_2067),
.Y(n_2309)
);

XOR2xp5_ASAP7_75t_L g2310 ( 
.A(n_2298),
.B(n_2014),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2304),
.Y(n_2311)
);

NOR2x1_ASAP7_75t_L g2312 ( 
.A(n_2303),
.B(n_2308),
.Y(n_2312)
);

CKINVDCx12_ASAP7_75t_R g2313 ( 
.A(n_2309),
.Y(n_2313)
);

CKINVDCx16_ASAP7_75t_R g2314 ( 
.A(n_2310),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2314),
.A2(n_2307),
.B1(n_2306),
.B2(n_2079),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2312),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2315),
.A2(n_2311),
.B1(n_2313),
.B2(n_2305),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2316),
.A2(n_2103),
.B(n_2089),
.Y(n_2318)
);

BUFx2_ASAP7_75t_L g2319 ( 
.A(n_2317),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_2318),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_2317),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2320),
.A2(n_2068),
.B1(n_2106),
.B2(n_2107),
.Y(n_2322)
);

XNOR2xp5_ASAP7_75t_L g2323 ( 
.A(n_2321),
.B(n_1968),
.Y(n_2323)
);

AOI222xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2323),
.A2(n_2319),
.B1(n_2023),
.B2(n_2019),
.C1(n_2091),
.C2(n_2107),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2322),
.Y(n_2325)
);

NAND3xp33_ASAP7_75t_L g2326 ( 
.A(n_2325),
.B(n_2106),
.C(n_2095),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_R g2327 ( 
.A1(n_2326),
.A2(n_2324),
.B1(n_2067),
.B2(n_2072),
.C(n_2155),
.Y(n_2327)
);

AOI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2327),
.A2(n_2097),
.B(n_2103),
.C(n_2099),
.Y(n_2328)
);


endmodule