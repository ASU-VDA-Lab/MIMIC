module fake_jpeg_31644_n_519 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_59),
.Y(n_118)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_28),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_8),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_7),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_74),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_9),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_96),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_9),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_34),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_100),
.B(n_103),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_29),
.B1(n_23),
.B2(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_110),
.A2(n_124),
.B1(n_64),
.B2(n_57),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_114),
.B(n_136),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_52),
.A2(n_29),
.B1(n_31),
.B2(n_37),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_74),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_88),
.A2(n_37),
.B1(n_31),
.B2(n_42),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_53),
.A2(n_50),
.B1(n_40),
.B2(n_38),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_56),
.A2(n_50),
.B1(n_40),
.B2(n_38),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_92),
.A2(n_37),
.B1(n_31),
.B2(n_42),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_68),
.A2(n_29),
.B(n_45),
.C(n_31),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_47),
.B(n_103),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_54),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_161),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_60),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_69),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_164),
.A2(n_167),
.B1(n_202),
.B2(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_112),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_189),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_84),
.B1(n_76),
.B2(n_99),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_173),
.B(n_13),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_22),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_150),
.B(n_128),
.C(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_181),
.B(n_45),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_106),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_120),
.A2(n_89),
.B1(n_83),
.B2(n_97),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_124),
.B1(n_144),
.B2(n_148),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_81),
.B1(n_102),
.B2(n_55),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_194),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_62),
.C(n_95),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_120),
.Y(n_196)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_37),
.B1(n_49),
.B2(n_47),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_49),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_144),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_129),
.A2(n_77),
.B1(n_86),
.B2(n_85),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_117),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_126),
.A2(n_103),
.B1(n_35),
.B2(n_45),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_147),
.A2(n_93),
.B1(n_39),
.B2(n_45),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_208),
.A2(n_209),
.B1(n_216),
.B2(n_109),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_126),
.A2(n_135),
.B1(n_107),
.B2(n_111),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_212),
.Y(n_242)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.Y(n_244)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_215),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_108),
.A2(n_45),
.B1(n_39),
.B2(n_2),
.Y(n_216)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_252),
.B1(n_258),
.B2(n_164),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_250),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_226),
.A2(n_0),
.B(n_1),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_238),
.B(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_175),
.B(n_157),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_253),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_10),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_202),
.A2(n_151),
.B1(n_110),
.B2(n_155),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_201),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_163),
.B(n_109),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_163),
.C(n_203),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_181),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_154),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_280),
.B1(n_281),
.B2(n_285),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_261),
.A2(n_183),
.B1(n_195),
.B2(n_167),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_284),
.B1(n_287),
.B2(n_298),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_265),
.B(n_275),
.Y(n_309)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_244),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_192),
.C(n_172),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_286),
.C(n_288),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_235),
.A2(n_165),
.B(n_189),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_180),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_274),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_200),
.B1(n_214),
.B2(n_199),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_176),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_187),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_178),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_282),
.Y(n_338)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g279 ( 
.A1(n_226),
.A2(n_198),
.A3(n_211),
.B1(n_205),
.B2(n_215),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_219),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_252),
.A2(n_196),
.B1(n_177),
.B2(n_217),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_196),
.B1(n_213),
.B2(n_193),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_179),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_210),
.B1(n_171),
.B2(n_39),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_184),
.B1(n_11),
.B2(n_3),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_227),
.C(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_194),
.C(n_1),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_299),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_228),
.Y(n_326)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_295),
.Y(n_339)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_219),
.B(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_242),
.B(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_249),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_301),
.A2(n_285),
.B1(n_281),
.B2(n_280),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_302),
.A2(n_246),
.B1(n_255),
.B2(n_259),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_320),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_263),
.A2(n_221),
.B1(n_224),
.B2(n_223),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_305),
.A2(n_307),
.B1(n_312),
.B2(n_314),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_306),
.B(n_318),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_221),
.B1(n_224),
.B2(n_243),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_220),
.B(n_236),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_310),
.A2(n_323),
.B(n_330),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_233),
.B1(n_245),
.B2(n_254),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_268),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_229),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_319),
.B(n_333),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_264),
.A2(n_254),
.B1(n_228),
.B2(n_255),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_236),
.B(n_262),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_289),
.B(n_229),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_275),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_293),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_262),
.B(n_232),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_337),
.B1(n_282),
.B2(n_276),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_270),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_222),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_269),
.C(n_274),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_297),
.A2(n_237),
.B1(n_222),
.B2(n_241),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_341),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_342),
.A2(n_348),
.B1(n_350),
.B2(n_362),
.Y(n_382)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_302),
.B1(n_298),
.B2(n_279),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_345),
.A2(n_267),
.B(n_283),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_297),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_354),
.C(n_313),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_329),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_351),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_310),
.A2(n_271),
.B(n_301),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_349),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_303),
.A2(n_291),
.B1(n_295),
.B2(n_288),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_338),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_358),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_353),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_306),
.B(n_269),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_272),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_363),
.Y(n_378)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_271),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_361),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_337),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_364),
.A2(n_327),
.B1(n_311),
.B2(n_314),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_339),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_367),
.A2(n_368),
.B1(n_370),
.B2(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_300),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_316),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_313),
.B(n_292),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_326),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_357),
.A2(n_303),
.B1(n_315),
.B2(n_327),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_374),
.A2(n_386),
.B1(n_398),
.B2(n_342),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_364),
.A2(n_315),
.B(n_323),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_393),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_382),
.B(n_367),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_363),
.A2(n_320),
.B1(n_311),
.B2(n_312),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_383),
.A2(n_385),
.B1(n_366),
.B2(n_368),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_388),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_357),
.A2(n_332),
.B1(n_330),
.B2(n_339),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_326),
.C(n_328),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_391),
.C(n_396),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_328),
.C(n_317),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_343),
.A2(n_317),
.B(n_296),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_237),
.C(n_324),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_331),
.C(n_324),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_350),
.C(n_362),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_343),
.A2(n_331),
.B(n_316),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_401),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_267),
.B(n_247),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_351),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_259),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_366),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_405),
.A2(n_385),
.B1(n_375),
.B2(n_393),
.Y(n_439)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_390),
.A2(n_341),
.B1(n_345),
.B2(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_400),
.Y(n_410)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_412),
.Y(n_436)
);

XOR2x2_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_358),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_423),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_352),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_417),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_426),
.C(n_427),
.Y(n_431)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_355),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_418),
.B(n_422),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_360),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_419),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_425),
.B1(n_386),
.B2(n_374),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_370),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_421),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_361),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_424),
.B(n_395),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_383),
.A2(n_359),
.B1(n_356),
.B2(n_344),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_232),
.C(n_278),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_294),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_266),
.C(n_234),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_429),
.C(n_387),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_234),
.Y(n_429)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_395),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_448),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_449),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_439),
.A2(n_420),
.B1(n_394),
.B2(n_405),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_373),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

OAI31xp33_ASAP7_75t_L g447 ( 
.A1(n_406),
.A2(n_398),
.A3(n_394),
.B(n_402),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_447),
.A2(n_402),
.B(n_422),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_373),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_418),
.B(n_388),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_427),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_426),
.C(n_404),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_453),
.C(n_463),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_404),
.C(n_428),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_456),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_401),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_459),
.A2(n_437),
.B1(n_438),
.B2(n_445),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_415),
.C(n_413),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_464),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g468 ( 
.A1(n_462),
.A2(n_447),
.B(n_432),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_423),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_465),
.Y(n_483)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_12),
.Y(n_481)
);

OAI221xp5_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_379),
.B1(n_392),
.B2(n_389),
.C(n_380),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_467),
.A2(n_397),
.B(n_429),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_479),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_443),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_470),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_449),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_471),
.A2(n_473),
.B1(n_478),
.B2(n_480),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_SL g472 ( 
.A(n_460),
.B(n_409),
.C(n_446),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_475),
.B(n_482),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_459),
.A2(n_432),
.B1(n_442),
.B2(n_441),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_461),
.A2(n_441),
.B(n_439),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_446),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_458),
.A2(n_440),
.B1(n_414),
.B2(n_409),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_0),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_462),
.A2(n_440),
.B(n_4),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_473),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_486),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_474),
.A2(n_482),
.B1(n_454),
.B2(n_451),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_452),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_492),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_464),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_491),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_453),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_5),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_5),
.C(n_10),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_495),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_5),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_5),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_475),
.B(n_483),
.C(n_468),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_498),
.A2(n_502),
.B(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_471),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_505),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g502 ( 
.A1(n_495),
.A2(n_478),
.B(n_470),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_13),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_12),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_500),
.B(n_491),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_501),
.A2(n_485),
.B1(n_489),
.B2(n_490),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_508),
.A2(n_510),
.B1(n_497),
.B2(n_499),
.Y(n_513)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_509),
.Y(n_511)
);

NAND2x1_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_513),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_512),
.A2(n_504),
.B(n_13),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_13),
.C(n_17),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_516),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_517),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_518),
.B(n_514),
.Y(n_519)
);


endmodule