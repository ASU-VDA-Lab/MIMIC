module fake_jpeg_30540_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_18),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_23),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_2),
.C(n_3),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.B(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_28),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_11),
.B1(n_8),
.B2(n_13),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_31),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_12),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_25),
.C(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_32),
.C(n_35),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_8),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_35),
.C(n_34),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_45),
.B(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_8),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_45),
.B(n_47),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_23),
.B2(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_23),
.Y(n_52)
);


endmodule