module fake_jpeg_21922_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_1),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_23),
.B1(n_24),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_24),
.B1(n_19),
.B2(n_12),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_12),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_46),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_18),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_23),
.B1(n_18),
.B2(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_10),
.B1(n_36),
.B2(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_39),
.B(n_35),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_72),
.C(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_44),
.C(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_63),
.B1(n_59),
.B2(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_83),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_63),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_64),
.B(n_66),
.C(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_88),
.B1(n_81),
.B2(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

BUFx12f_ASAP7_75t_SL g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_88),
.C(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_89),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_97),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.Y(n_103)
);


endmodule