module fake_jpeg_19065_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_30),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_30),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_60),
.B1(n_68),
.B2(n_43),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_17),
.Y(n_78)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_37),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_69),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_35),
.B1(n_25),
.B2(n_23),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_26),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_19),
.CON(n_75),
.SN(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_30),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_56),
.B(n_74),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_76),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_97),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_43),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g134 ( 
.A(n_89),
.B(n_101),
.Y(n_134)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_106),
.B1(n_112),
.B2(n_67),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_110),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_48),
.B1(n_46),
.B2(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_48),
.B1(n_71),
.B2(n_17),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_16),
.B1(n_18),
.B2(n_26),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_67),
.B1(n_36),
.B2(n_18),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_28),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_28),
.C(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_121),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_125),
.B1(n_86),
.B2(n_96),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_33),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_49),
.B1(n_45),
.B2(n_18),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_149),
.B1(n_113),
.B2(n_77),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_145),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_16),
.B1(n_29),
.B2(n_36),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_106),
.B1(n_110),
.B2(n_101),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_19),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_58),
.C(n_82),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_90),
.A2(n_36),
.B1(n_29),
.B2(n_58),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_103),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_163),
.B1(n_167),
.B2(n_171),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_158),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_87),
.B1(n_98),
.B2(n_94),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_160),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_124),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_85),
.B1(n_81),
.B2(n_80),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_173),
.B1(n_183),
.B2(n_160),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_144),
.B1(n_121),
.B2(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_118),
.B1(n_129),
.B2(n_126),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_130),
.B1(n_136),
.B2(n_123),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_58),
.B1(n_57),
.B2(n_33),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_82),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_103),
.B1(n_82),
.B2(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_177),
.Y(n_201)
);

HAxp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_19),
.CON(n_178),
.SN(n_178)
);

AOI32xp33_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_21),
.A3(n_22),
.B1(n_8),
.B2(n_9),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_185),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_159),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_189),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_138),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_215),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_143),
.B1(n_145),
.B2(n_118),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_192),
.A2(n_202),
.B1(n_166),
.B2(n_156),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_199),
.B1(n_200),
.B2(n_174),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_21),
.B(n_132),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_177),
.B(n_170),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_126),
.B(n_21),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_208),
.B(n_212),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_34),
.C(n_129),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_204),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_181),
.B1(n_157),
.B2(n_168),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_34),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_166),
.B1(n_183),
.B2(n_164),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_6),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_226),
.B1(n_239),
.B2(n_244),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_240),
.B1(n_243),
.B2(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_159),
.C(n_157),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_237),
.C(n_241),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_228),
.B(n_229),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_232),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_194),
.B1(n_217),
.B2(n_201),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_13),
.C(n_6),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_6),
.B1(n_11),
.B2(n_9),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_186),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_12),
.C(n_7),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_7),
.B1(n_12),
.B2(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_188),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_221),
.B1(n_223),
.B2(n_225),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_189),
.B1(n_199),
.B2(n_206),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_253),
.A2(n_239),
.B1(n_244),
.B2(n_240),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_188),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_249),
.B(n_195),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_215),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_214),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_207),
.Y(n_261)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_196),
.Y(n_268)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_227),
.B(n_187),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_227),
.B(n_242),
.Y(n_274)
);

AOI31xp33_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_211),
.A3(n_236),
.B(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_234),
.B1(n_222),
.B2(n_223),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_277),
.B1(n_251),
.B2(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_282),
.B1(n_256),
.B2(n_246),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_273),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_276),
.B(n_278),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_196),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_241),
.C(n_202),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_7),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_260),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_259),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_284),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_289),
.B1(n_267),
.B2(n_274),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_257),
.B1(n_265),
.B2(n_263),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_265),
.B(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_293),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_247),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_272),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_12),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_277),
.B1(n_278),
.B2(n_273),
.Y(n_303)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_306),
.B1(n_289),
.B2(n_285),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_280),
.C(n_260),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_307),
.C(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_259),
.B1(n_255),
.B2(n_283),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_3),
.B(n_4),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_316),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_287),
.B1(n_294),
.B2(n_298),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_293),
.C(n_295),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_301),
.B(n_307),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_320),
.C(n_322),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_299),
.B1(n_300),
.B2(n_4),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_300),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_318),
.B(n_314),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_309),
.B(n_322),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_327),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_319),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_311),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_323),
.Y(n_333)
);


endmodule