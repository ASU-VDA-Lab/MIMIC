module fake_netlist_1_677_n_1240 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1240);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1240;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_283;
wire n_756;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_270;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1195;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
HB1xp67_ASAP7_75t_L g269 ( .A(n_215), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_112), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_119), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_102), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_226), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_4), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_158), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_4), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_135), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_233), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_100), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_133), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_28), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_71), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_113), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_149), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_52), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_208), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_140), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_202), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_29), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_205), .Y(n_290) );
CKINVDCx14_ASAP7_75t_R g291 ( .A(n_16), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_192), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_97), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_28), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_34), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_137), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_136), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_123), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_134), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_0), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_178), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_87), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_124), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_131), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_75), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_260), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_79), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_142), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_250), .B(n_198), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_6), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_241), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_224), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_12), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_82), .Y(n_315) );
INVxp33_ASAP7_75t_SL g316 ( .A(n_78), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_235), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_76), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_64), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_187), .Y(n_320) );
BUFx5_ASAP7_75t_L g321 ( .A(n_212), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_144), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_50), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_48), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_69), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_25), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_176), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_164), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_152), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_27), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_228), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_243), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_213), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_214), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_37), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_180), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_191), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_90), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_193), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_240), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_105), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_96), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_128), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_109), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_181), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_265), .B(n_261), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_170), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_238), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_216), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_160), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_34), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_68), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_44), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_46), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_266), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_52), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_70), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_17), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_229), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_211), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_48), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_83), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_162), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_199), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_84), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_117), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_166), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_157), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_174), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_104), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_118), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_23), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_16), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_29), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_245), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_120), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_36), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_194), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_165), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_249), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_255), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_251), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_239), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_148), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_167), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_13), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_47), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_179), .Y(n_388) );
INVxp33_ASAP7_75t_SL g389 ( .A(n_30), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_59), .B(n_88), .Y(n_390) );
BUFx5_ASAP7_75t_L g391 ( .A(n_65), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_43), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_143), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_31), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_60), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_132), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_155), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_72), .B(n_227), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_111), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_59), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_125), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_263), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_321), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_318), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_363), .B(n_0), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_321), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_321), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_321), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_386), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_289), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_289), .Y(n_411) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_386), .B(n_1), .Y(n_412) );
BUFx8_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_300), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_300), .B(n_1), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_291), .Y(n_416) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_346), .B(n_66), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_319), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_319), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_277), .A2(n_307), .B(n_288), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_298), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_321), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_373), .B(n_2), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_271), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_278), .Y(n_426) );
OA21x2_ASAP7_75t_L g427 ( .A1(n_277), .A2(n_73), .B(n_67), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_280), .Y(n_428) );
AND2x6_ASAP7_75t_L g429 ( .A(n_298), .B(n_74), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_283), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_291), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_431) );
INVx5_ASAP7_75t_L g432 ( .A(n_305), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_284), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_321), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_389), .A2(n_3), .B1(n_5), .B2(n_7), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_415), .A2(n_274), .B1(n_285), .B2(n_281), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_404), .B(n_362), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_429), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_415), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_404), .B(n_326), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_403), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_425), .B(n_269), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_416), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_415), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_415), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_424), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_425), .B(n_282), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_417), .A2(n_389), .B1(n_303), .B2(n_312), .Y(n_450) );
OR2x6_ASAP7_75t_L g451 ( .A(n_431), .B(n_330), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
AND2x6_ASAP7_75t_L g453 ( .A(n_424), .B(n_390), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_426), .B(n_394), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_426), .B(n_328), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_405), .B(n_394), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_422), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_428), .B(n_297), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_406), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_422), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_420), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
BUFx10_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_408), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_408), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_417), .A2(n_303), .B1(n_312), .B2(n_270), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_428), .B(n_297), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_430), .B(n_347), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_347), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_408), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
INVx4_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
NAND2xp33_ASAP7_75t_SL g479 ( .A(n_405), .B(n_270), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_424), .B(n_294), .Y(n_480) );
OR2x6_ASAP7_75t_L g481 ( .A(n_431), .B(n_295), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_413), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_445), .A2(n_420), .B(n_427), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_475), .B(n_417), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_450), .A2(n_413), .B1(n_424), .B2(n_339), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_475), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_463), .A2(n_413), .B1(n_324), .B2(n_392), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_458), .B(n_433), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_482), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_439), .Y(n_491) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_451), .A2(n_435), .B1(n_324), .B2(n_392), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_458), .B(n_455), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_440), .B(n_433), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_438), .B(n_350), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_440), .B(n_354), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_445), .A2(n_420), .B(n_427), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_409), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_479), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_480), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_473), .B(n_420), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_438), .B(n_350), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_439), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_474), .B(n_409), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_480), .B(n_453), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_480), .B(n_409), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_409), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_444), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_453), .A2(n_339), .B1(n_344), .B2(n_343), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_469), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_444), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_451), .B(n_435), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_453), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_453), .A2(n_343), .B1(n_375), .B2(n_344), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_437), .B(n_412), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_436), .B(n_377), .C(n_356), .Y(n_520) );
INVx3_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_442), .B(n_316), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_453), .A2(n_412), .B1(n_316), .B2(n_429), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_451), .B(n_358), .Y(n_524) );
NOR2x1p5_ASAP7_75t_L g525 ( .A(n_449), .B(n_396), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_446), .B(n_304), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_453), .A2(n_429), .B1(n_434), .B2(n_423), .Y(n_527) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_453), .B(n_429), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_456), .B(n_446), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_446), .B(n_423), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_447), .B(n_399), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_472), .A2(n_380), .B1(n_384), .B2(n_375), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_447), .B(n_366), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_451), .A2(n_276), .B1(n_384), .B2(n_380), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_447), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_447), .Y(n_536) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_467), .B(n_429), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_451), .B(n_410), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_481), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_441), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_460), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_472), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_481), .Y(n_543) );
NOR2x2_ASAP7_75t_L g544 ( .A(n_481), .B(n_276), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_481), .B(n_410), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_441), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_448), .B(n_434), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_443), .B(n_411), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_448), .Y(n_550) );
AND2x6_ASAP7_75t_L g551 ( .A(n_454), .B(n_315), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_469), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_454), .B(n_429), .Y(n_553) );
INVx5_ASAP7_75t_L g554 ( .A(n_438), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_459), .B(n_399), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_443), .B(n_411), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_459), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_457), .A2(n_314), .B1(n_323), .B2(n_310), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_457), .A2(n_335), .B1(n_353), .B2(n_351), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_462), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_465), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_462), .B(n_402), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_465), .A2(n_427), .B(n_309), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_464), .A2(n_372), .B1(n_374), .B2(n_361), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_464), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_466), .B(n_471), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_478), .B(n_414), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_414), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_471), .A2(n_387), .B1(n_400), .B2(n_395), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_550), .Y(n_570) );
INVx3_ASAP7_75t_SL g571 ( .A(n_544), .Y(n_571) );
CKINVDCx14_ASAP7_75t_R g572 ( .A(n_524), .Y(n_572) );
INVx4_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_502), .A2(n_478), .B(n_477), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_554), .B(n_478), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_493), .B(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_489), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_554), .B(n_469), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_566), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_493), .A2(n_468), .B(n_470), .C(n_452), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_484), .A2(n_468), .B(n_470), .C(n_452), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_568), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_488), .B(n_452), .Y(n_584) );
BUFx10_ASAP7_75t_L g585 ( .A(n_488), .Y(n_585) );
CKINVDCx16_ASAP7_75t_R g586 ( .A(n_524), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_484), .A2(n_470), .B(n_476), .C(n_468), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_501), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_554), .B(n_273), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_494), .B(n_476), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_490), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_554), .B(n_275), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_512), .A2(n_419), .B1(n_421), .B2(n_418), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_487), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_489), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_521), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_517), .B(n_279), .Y(n_597) );
OAI21x1_ASAP7_75t_SL g598 ( .A1(n_539), .A2(n_427), .B(n_388), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_543), .A2(n_476), .B1(n_286), .B2(n_364), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_486), .A2(n_418), .B(n_421), .C(n_419), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_496), .B(n_272), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_522), .B(n_342), .Y(n_602) );
OAI22x1_ASAP7_75t_L g603 ( .A1(n_532), .A2(n_360), .B1(n_308), .B2(n_311), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_534), .B(n_7), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_519), .B(n_292), .Y(n_605) );
O2A1O1Ixp5_ASAP7_75t_L g606 ( .A1(n_528), .A2(n_288), .B(n_337), .C(n_307), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_519), .B(n_357), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_502), .A2(n_497), .B(n_483), .Y(n_608) );
OR2x6_ASAP7_75t_L g609 ( .A(n_516), .B(n_352), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_545), .A2(n_290), .B(n_293), .C(n_287), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_513), .B(n_359), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_521), .Y(n_612) );
BUFx3_ASAP7_75t_L g613 ( .A(n_549), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_537), .A2(n_299), .B(n_296), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_563), .A2(n_302), .B(n_301), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_560), .B(n_365), .Y(n_616) );
NOR2xp67_ASAP7_75t_SL g617 ( .A(n_506), .B(n_379), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_562), .B(n_306), .Y(n_618) );
CKINVDCx8_ASAP7_75t_R g619 ( .A(n_500), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_538), .A2(n_317), .B(n_320), .C(n_313), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_518), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_556), .B(n_322), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_491), .A2(n_498), .B(n_507), .C(n_504), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_530), .A2(n_327), .B(n_325), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_485), .Y(n_625) );
BUFx12f_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_492), .A2(n_329), .B(n_332), .C(n_331), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_530), .A2(n_336), .B(n_333), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_508), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_514), .A2(n_340), .B(n_338), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_506), .B(n_341), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_553), .A2(n_348), .B(n_345), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_515), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_529), .A2(n_505), .B(n_499), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_542), .B(n_8), .Y(n_636) );
CKINVDCx8_ASAP7_75t_R g637 ( .A(n_551), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
NOR3xp33_ASAP7_75t_SL g639 ( .A(n_520), .B(n_355), .C(n_349), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_562), .B(n_367), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_535), .Y(n_641) );
INVx8_ASAP7_75t_L g642 ( .A(n_551), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_508), .Y(n_643) );
NOR2xp33_ASAP7_75t_SL g644 ( .A(n_513), .B(n_398), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_509), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_536), .A2(n_376), .B(n_401), .C(n_397), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_531), .B(n_368), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_505), .A2(n_370), .B(n_369), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g649 ( .A1(n_509), .A2(n_382), .B(n_383), .C(n_371), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_559), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_551), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_495), .A2(n_393), .B(n_381), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_547), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_551), .Y(n_655) );
CKINVDCx10_ASAP7_75t_R g656 ( .A(n_564), .Y(n_656) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_510), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_523), .B(n_555), .Y(n_658) );
BUFx10_ASAP7_75t_L g659 ( .A(n_526), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_558), .B(n_315), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_541), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_513), .B(n_385), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_546), .B(n_385), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_546), .B(n_321), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_533), .B(n_8), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_503), .B(n_9), .C(n_10), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_548), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_569), .B(n_391), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_567), .A2(n_334), .B(n_305), .C(n_432), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_546), .B(n_305), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_548), .Y(n_671) );
INVx4_ASAP7_75t_L g672 ( .A(n_552), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_552), .B(n_391), .Y(n_673) );
BUFx4f_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g675 ( .A1(n_561), .A2(n_9), .B(n_10), .C(n_11), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_552), .B(n_391), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_527), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_502), .A2(n_432), .B(n_334), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_554), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_488), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_496), .B(n_11), .Y(n_681) );
CKINVDCx6p67_ASAP7_75t_R g682 ( .A(n_524), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_566), .Y(n_683) );
BUFx2_ASAP7_75t_L g684 ( .A(n_524), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_493), .A2(n_12), .B(n_13), .C(n_14), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_550), .Y(n_686) );
INVx1_ASAP7_75t_SL g687 ( .A(n_550), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_566), .Y(n_688) );
OR2x6_ASAP7_75t_L g689 ( .A(n_524), .B(n_334), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_493), .A2(n_14), .B(n_15), .C(n_17), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_502), .A2(n_432), .B(n_391), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_566), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_493), .B(n_391), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_484), .A2(n_391), .B1(n_432), .B2(n_19), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_502), .A2(n_432), .B(n_391), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_493), .A2(n_15), .B(n_18), .C(n_19), .Y(n_696) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_554), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_493), .B(n_18), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_577), .B(n_20), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_580), .Y(n_700) );
OAI221xp5_ASAP7_75t_SL g701 ( .A1(n_627), .A2(n_20), .B1(n_21), .B2(n_22), .C(n_23), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g702 ( .A1(n_658), .A2(n_147), .B(n_268), .C(n_267), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_608), .A2(n_432), .B(n_77), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_683), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_688), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_586), .B(n_21), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_692), .A2(n_22), .B(n_24), .C(n_25), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_635), .A2(n_24), .B(n_26), .C(n_27), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_687), .Y(n_709) );
AO31x2_ASAP7_75t_L g710 ( .A1(n_615), .A2(n_26), .A3(n_30), .B(n_31), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_667), .Y(n_711) );
AO21x1_ASAP7_75t_L g712 ( .A1(n_678), .A2(n_81), .B(n_80), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_671), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_621), .A2(n_32), .B1(n_33), .B2(n_35), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_583), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_585), .B(n_32), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_576), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_651), .A2(n_33), .B1(n_35), .B2(n_36), .C(n_37), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_654), .B(n_38), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_585), .B(n_38), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_SL g721 ( .A1(n_623), .A2(n_163), .B(n_262), .C(n_259), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_646), .A2(n_39), .B(n_40), .C(n_41), .Y(n_722) );
AO31x2_ASAP7_75t_L g723 ( .A1(n_691), .A2(n_39), .A3(n_40), .B(n_41), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_SL g724 ( .A1(n_669), .A2(n_168), .B(n_258), .C(n_257), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_665), .A2(n_42), .B(n_43), .C(n_44), .Y(n_725) );
INVxp33_ASAP7_75t_L g726 ( .A(n_636), .Y(n_726) );
INVx8_ASAP7_75t_L g727 ( .A(n_689), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_574), .A2(n_161), .B(n_256), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g729 ( .A1(n_581), .A2(n_159), .B(n_253), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_682), .A2(n_42), .B1(n_45), .B2(n_46), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_689), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_679), .Y(n_732) );
AND2x6_ASAP7_75t_SL g733 ( .A(n_604), .B(n_45), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_695), .A2(n_47), .A3(n_49), .B(n_50), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g735 ( .A1(n_582), .A2(n_172), .B(n_252), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_572), .A2(n_51), .B1(n_53), .B2(n_54), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_650), .Y(n_737) );
NOR2xp67_ASAP7_75t_L g738 ( .A(n_591), .B(n_51), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_638), .Y(n_739) );
BUFx2_ASAP7_75t_L g740 ( .A(n_689), .Y(n_740) );
INVx3_ASAP7_75t_SL g741 ( .A(n_571), .Y(n_741) );
AO32x1_ASAP7_75t_L g742 ( .A1(n_599), .A2(n_53), .A3(n_54), .B1(n_55), .B2(n_56), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_625), .B(n_55), .Y(n_743) );
AO32x2_ASAP7_75t_L g744 ( .A1(n_573), .A2(n_56), .A3(n_57), .B1(n_58), .B2(n_60), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_680), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_613), .B(n_57), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_594), .A2(n_58), .B1(n_61), .B2(n_62), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_L g748 ( .A1(n_698), .A2(n_61), .B(n_62), .C(n_63), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_684), .B(n_63), .Y(n_749) );
OAI21x1_ASAP7_75t_L g750 ( .A1(n_670), .A2(n_85), .B(n_86), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_573), .A2(n_89), .B1(n_91), .B2(n_92), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_614), .A2(n_93), .B(n_94), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_647), .A2(n_95), .B(n_98), .C(n_99), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_590), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_681), .B(n_101), .Y(n_755) );
OR2x6_ASAP7_75t_L g756 ( .A(n_642), .B(n_103), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_610), .A2(n_106), .B(n_107), .C(n_108), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_649), .A2(n_110), .B(n_114), .C(n_115), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_638), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_694), .A2(n_116), .B1(n_121), .B2(n_122), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_584), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_587), .A2(n_126), .B(n_127), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_640), .A2(n_129), .B(n_130), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_622), .A2(n_601), .B1(n_593), .B2(n_603), .C(n_600), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_629), .B(n_138), .Y(n_765) );
OAI21x1_ASAP7_75t_SL g766 ( .A1(n_694), .A2(n_139), .B(n_141), .Y(n_766) );
INVx3_ASAP7_75t_L g767 ( .A(n_697), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_687), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_602), .A2(n_145), .B1(n_146), .B2(n_150), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_643), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_609), .A2(n_151), .B1(n_153), .B2(n_154), .Y(n_771) );
BUFx4_ASAP7_75t_SL g772 ( .A(n_609), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_645), .B(n_156), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_656), .Y(n_774) );
INVx2_ASAP7_75t_SL g775 ( .A(n_674), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_619), .B(n_169), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_609), .B(n_171), .Y(n_777) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_633), .A2(n_173), .B(n_175), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_L g779 ( .A1(n_620), .A2(n_177), .B(n_182), .C(n_183), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_630), .Y(n_780) );
AO31x2_ASAP7_75t_L g781 ( .A1(n_677), .A2(n_184), .A3(n_185), .B(n_186), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_693), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_SL g783 ( .A1(n_617), .A2(n_188), .B(n_189), .C(n_190), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_570), .B(n_195), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_686), .B(n_264), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_606), .A2(n_196), .B(n_197), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_637), .A2(n_200), .B1(n_201), .B2(n_203), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_634), .Y(n_788) );
AND2x4_ASAP7_75t_L g789 ( .A(n_588), .B(n_248), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_652), .B(n_204), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_660), .Y(n_791) );
BUFx3_ASAP7_75t_L g792 ( .A(n_626), .Y(n_792) );
NAND2xp33_ASAP7_75t_L g793 ( .A(n_642), .B(n_206), .Y(n_793) );
INVx2_ASAP7_75t_SL g794 ( .A(n_674), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_642), .A2(n_207), .B1(n_209), .B2(n_210), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_641), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_618), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_797) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_697), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_605), .B(n_220), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_660), .B(n_221), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_575), .A2(n_222), .B(n_223), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_656), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_607), .B(n_225), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_661), .Y(n_804) );
O2A1O1Ixp33_ASAP7_75t_L g805 ( .A1(n_685), .A2(n_230), .B(n_231), .C(n_232), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_659), .B(n_234), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_659), .B(n_236), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_L g808 ( .A1(n_690), .A2(n_237), .B(n_242), .C(n_244), .Y(n_808) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_697), .Y(n_809) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_616), .Y(n_810) );
A2O1A1Ixp33_ASAP7_75t_L g811 ( .A1(n_648), .A2(n_246), .B(n_247), .C(n_628), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_657), .Y(n_812) );
INVxp67_ASAP7_75t_L g813 ( .A(n_611), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_624), .A2(n_696), .B(n_675), .C(n_631), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_631), .B(n_632), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_664), .A2(n_676), .B(n_673), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_666), .A2(n_578), .B1(n_596), .B2(n_595), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_612), .A2(n_668), .B1(n_657), .B2(n_655), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_672), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_662), .A2(n_663), .B(n_653), .Y(n_820) );
A2O1A1Ixp33_ASAP7_75t_L g821 ( .A1(n_639), .A2(n_644), .B(n_597), .C(n_592), .Y(n_821) );
NAND3x1_ASAP7_75t_L g822 ( .A(n_644), .B(n_611), .C(n_589), .Y(n_822) );
A2O1A1Ixp33_ASAP7_75t_L g823 ( .A1(n_579), .A2(n_577), .B(n_683), .C(n_580), .Y(n_823) );
NAND2x1p5_ASAP7_75t_L g824 ( .A(n_672), .B(n_573), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_SL g825 ( .A1(n_658), .A2(n_502), .B(n_623), .C(n_669), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_625), .B(n_651), .Y(n_826) );
OR2x6_ASAP7_75t_L g827 ( .A(n_573), .B(n_524), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_635), .A2(n_574), .B(n_608), .Y(n_828) );
BUFx2_ASAP7_75t_L g829 ( .A(n_689), .Y(n_829) );
O2A1O1Ixp33_ASAP7_75t_SL g830 ( .A1(n_658), .A2(n_502), .B(n_623), .C(n_669), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g831 ( .A1(n_689), .A2(n_625), .B(n_493), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g832 ( .A1(n_577), .A2(n_580), .B(n_683), .C(n_688), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_828), .A2(n_830), .B(n_825), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_L g834 ( .A1(n_832), .A2(n_810), .B(n_725), .C(n_814), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_826), .A2(n_764), .B1(n_791), .B2(n_717), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_717), .B(n_700), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_831), .B(n_709), .Y(n_837) );
AO31x2_ASAP7_75t_L g838 ( .A1(n_712), .A2(n_823), .A3(n_703), .B(n_758), .Y(n_838) );
OAI21xp33_ASAP7_75t_SL g839 ( .A1(n_756), .A2(n_755), .B(n_711), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g840 ( .A1(n_747), .A2(n_701), .B1(n_743), .B2(n_730), .C(n_718), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_700), .B(n_711), .Y(n_841) );
INVx1_ASAP7_75t_SL g842 ( .A(n_713), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_754), .B(n_704), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_705), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_827), .B(n_770), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_761), .B(n_782), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_765), .A2(n_773), .B(n_815), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_737), .Y(n_848) );
OA21x2_ASAP7_75t_L g849 ( .A1(n_729), .A2(n_786), .B(n_762), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_714), .A2(n_736), .B1(n_719), .B2(n_746), .C(n_817), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_820), .A2(n_811), .B(n_793), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_816), .A2(n_721), .B(n_805), .Y(n_852) );
BUFx2_ASAP7_75t_L g853 ( .A(n_827), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_726), .A2(n_722), .B1(n_745), .B2(n_748), .C(n_760), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_749), .A2(n_777), .B1(n_727), .B2(n_720), .Y(n_855) );
OR2x6_ASAP7_75t_L g856 ( .A(n_727), .B(n_756), .Y(n_856) );
A2O1A1Ixp33_ASAP7_75t_L g857 ( .A1(n_757), .A2(n_779), .B(n_808), .C(n_803), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_716), .A2(n_699), .B1(n_789), .B2(n_829), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_780), .B(n_788), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_780), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_802), .B(n_706), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_796), .B(n_759), .Y(n_862) );
AO31x2_ASAP7_75t_L g863 ( .A1(n_708), .A2(n_753), .A3(n_797), .B(n_728), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_789), .A2(n_740), .B1(n_731), .B2(n_806), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_800), .A2(n_783), .B(n_702), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_739), .B(n_804), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_768), .B(n_799), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_724), .A2(n_778), .B(n_821), .Y(n_868) );
OA21x2_ASAP7_75t_L g869 ( .A1(n_766), .A2(n_750), .B(n_752), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_710), .Y(n_870) );
AO31x2_ASAP7_75t_L g871 ( .A1(n_707), .A2(n_795), .A3(n_787), .B(n_801), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_710), .Y(n_872) );
OA21x2_ASAP7_75t_L g873 ( .A1(n_763), .A2(n_769), .B(n_784), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_818), .B(n_767), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_784), .A2(n_785), .B(n_790), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_785), .A2(n_790), .B(n_751), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_738), .A2(n_776), .B1(n_813), .B2(n_771), .C(n_741), .Y(n_877) );
O2A1O1Ixp33_ASAP7_75t_L g878 ( .A1(n_819), .A2(n_812), .B(n_807), .C(n_775), .Y(n_878) );
AO21x2_ASAP7_75t_L g879 ( .A1(n_781), .A2(n_809), .B(n_723), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_798), .B(n_767), .Y(n_880) );
AOI33xp33_ASAP7_75t_L g881 ( .A1(n_794), .A2(n_733), .A3(n_772), .B1(n_744), .B2(n_710), .B3(n_742), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_774), .A2(n_792), .B1(n_824), .B2(n_732), .C(n_798), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_732), .B(n_723), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_723), .B(n_734), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_744), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_744), .B(n_734), .Y(n_886) );
BUFx2_ASAP7_75t_L g887 ( .A(n_822), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_734), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_742), .A2(n_826), .B1(n_542), .B2(n_621), .Y(n_889) );
BUFx3_ASAP7_75t_L g890 ( .A(n_781), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_781), .B(n_625), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_832), .A2(n_828), .B(n_635), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_713), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_827), .Y(n_894) );
BUFx3_ASAP7_75t_L g895 ( .A(n_741), .Y(n_895) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_764), .A2(n_534), .B(n_485), .Y(n_896) );
OAI221xp5_ASAP7_75t_SL g897 ( .A1(n_764), .A2(n_492), .B1(n_451), .B2(n_516), .C(n_532), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_715), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_832), .A2(n_828), .B(n_635), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_826), .B(n_524), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_715), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_713), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_826), .A2(n_450), .B1(n_534), .B2(n_472), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_717), .B(n_577), .Y(n_904) );
BUFx2_ASAP7_75t_L g905 ( .A(n_827), .Y(n_905) );
INVx3_ASAP7_75t_L g906 ( .A(n_727), .Y(n_906) );
AND2x2_ASAP7_75t_SL g907 ( .A(n_731), .B(n_586), .Y(n_907) );
AO31x2_ASAP7_75t_L g908 ( .A1(n_712), .A2(n_814), .A3(n_615), .B(n_823), .Y(n_908) );
OR2x6_ASAP7_75t_L g909 ( .A(n_727), .B(n_756), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_828), .A2(n_537), .B(n_608), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_715), .A2(n_492), .B1(n_627), .B2(n_651), .C(n_622), .Y(n_911) );
INVx3_ASAP7_75t_L g912 ( .A(n_727), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_715), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g914 ( .A1(n_828), .A2(n_537), .B(n_608), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_709), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_774), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_709), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_709), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_717), .B(n_577), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_713), .Y(n_920) );
A2O1A1Ixp33_ASAP7_75t_L g921 ( .A1(n_717), .A2(n_832), .B(n_577), .C(n_683), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_717), .B(n_700), .Y(n_922) );
AO21x2_ASAP7_75t_L g923 ( .A1(n_735), .A2(n_598), .B(n_828), .Y(n_923) );
INVx8_ASAP7_75t_L g924 ( .A(n_727), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_826), .B(n_524), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_826), .B(n_524), .Y(n_926) );
OR2x6_ASAP7_75t_L g927 ( .A(n_727), .B(n_756), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_826), .B(n_524), .Y(n_928) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_727), .A2(n_472), .B1(n_518), .B2(n_512), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_826), .B(n_524), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_709), .Y(n_931) );
INVx11_ASAP7_75t_L g932 ( .A(n_772), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_826), .B(n_458), .Y(n_933) );
INVx2_ASAP7_75t_SL g934 ( .A(n_772), .Y(n_934) );
INVx2_ASAP7_75t_L g935 ( .A(n_713), .Y(n_935) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_727), .A2(n_450), .B1(n_572), .B2(n_586), .Y(n_936) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_828), .A2(n_537), .B(n_608), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_832), .A2(n_828), .B(n_635), .Y(n_938) );
AO21x2_ASAP7_75t_L g939 ( .A1(n_833), .A2(n_884), .B(n_892), .Y(n_939) );
AO21x2_ASAP7_75t_L g940 ( .A1(n_884), .A2(n_938), .B(n_899), .Y(n_940) );
INVx3_ASAP7_75t_L g941 ( .A(n_922), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_856), .A2(n_909), .B1(n_927), .B2(n_903), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_841), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_924), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_841), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_911), .B(n_835), .Y(n_946) );
OA21x2_ASAP7_75t_L g947 ( .A1(n_892), .A2(n_899), .B(n_888), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_915), .Y(n_948) );
INVx3_ASAP7_75t_L g949 ( .A(n_922), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_836), .B(n_842), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_836), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_860), .Y(n_952) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_917), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_842), .B(n_859), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_870), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_880), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_859), .B(n_904), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_904), .B(n_919), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_872), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_893), .B(n_902), .Y(n_960) );
OAI31xp33_ASAP7_75t_L g961 ( .A1(n_897), .A2(n_896), .A3(n_929), .B(n_850), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_920), .B(n_935), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_844), .B(n_843), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_883), .B(n_880), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_911), .B(n_933), .Y(n_965) );
BUFx2_ASAP7_75t_L g966 ( .A(n_839), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_843), .B(n_848), .Y(n_967) );
OR2x6_ASAP7_75t_L g968 ( .A(n_875), .B(n_876), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_846), .B(n_921), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_883), .Y(n_970) );
BUFx3_ASAP7_75t_L g971 ( .A(n_924), .Y(n_971) );
AO21x2_ASAP7_75t_L g972 ( .A1(n_937), .A2(n_914), .B(n_910), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_852), .A2(n_851), .B(n_865), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_918), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_900), .B(n_925), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_898), .B(n_901), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_862), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_890), .Y(n_978) );
INVxp33_ASAP7_75t_L g979 ( .A(n_931), .Y(n_979) );
OR2x6_ASAP7_75t_L g980 ( .A(n_856), .B(n_927), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_879), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_840), .A2(n_936), .B1(n_850), .B2(n_854), .C(n_858), .Y(n_982) );
AO21x2_ASAP7_75t_L g983 ( .A1(n_886), .A2(n_923), .B(n_847), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_913), .B(n_862), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_866), .B(n_889), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_881), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_856), .Y(n_987) );
AOI22xp5_ASAP7_75t_L g988 ( .A1(n_840), .A2(n_927), .B1(n_909), .B2(n_928), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_923), .A2(n_868), .B(n_891), .Y(n_989) );
NOR2xp33_ASAP7_75t_SL g990 ( .A(n_934), .B(n_909), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_926), .B(n_930), .Y(n_991) );
HB1xp67_ASAP7_75t_L g992 ( .A(n_845), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_874), .Y(n_993) );
BUFx2_ASAP7_75t_L g994 ( .A(n_885), .Y(n_994) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_878), .Y(n_995) );
AO21x1_ASAP7_75t_SL g996 ( .A1(n_864), .A2(n_867), .B(n_855), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_845), .B(n_907), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_861), .B(n_894), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_834), .B(n_867), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_882), .B(n_905), .Y(n_1000) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_924), .Y(n_1001) );
INVxp67_ASAP7_75t_SL g1002 ( .A(n_837), .Y(n_1002) );
AO21x2_ASAP7_75t_L g1003 ( .A1(n_857), .A2(n_877), .B(n_908), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_908), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_869), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_853), .B(n_882), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_906), .B(n_912), .Y(n_1007) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_906), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_873), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_887), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_912), .B(n_871), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_869), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_932), .B(n_877), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_895), .A2(n_873), .B1(n_849), .B2(n_871), .C(n_863), .Y(n_1014) );
AO21x2_ASAP7_75t_L g1015 ( .A1(n_838), .A2(n_849), .B(n_863), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_838), .B(n_863), .Y(n_1016) );
INVx5_ASAP7_75t_SL g1017 ( .A(n_916), .Y(n_1017) );
INVxp67_ASAP7_75t_L g1018 ( .A(n_948), .Y(n_1018) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_980), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_954), .B(n_950), .Y(n_1020) );
NAND3xp33_ASAP7_75t_L g1021 ( .A(n_961), .B(n_982), .C(n_986), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_950), .B(n_957), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_994), .B(n_993), .Y(n_1023) );
NOR2x1_ASAP7_75t_L g1024 ( .A(n_980), .B(n_942), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_957), .B(n_958), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_994), .B(n_993), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_966), .A2(n_990), .B1(n_987), .B2(n_1000), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_1011), .B(n_964), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_976), .Y(n_1029) );
OR2x2_ASAP7_75t_SL g1030 ( .A(n_1010), .B(n_986), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_955), .Y(n_1031) );
INVx1_ASAP7_75t_SL g1032 ( .A(n_944), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_959), .Y(n_1033) );
AO21x2_ASAP7_75t_L g1034 ( .A1(n_973), .A2(n_1012), .B(n_1014), .Y(n_1034) );
INVx4_ASAP7_75t_L g1035 ( .A(n_980), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_963), .Y(n_1036) );
AO21x2_ASAP7_75t_L g1037 ( .A1(n_1012), .A2(n_972), .B(n_1005), .Y(n_1037) );
BUFx2_ASAP7_75t_SL g1038 ( .A(n_944), .Y(n_1038) );
AO21x2_ASAP7_75t_L g1039 ( .A1(n_972), .A2(n_1005), .B(n_981), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_963), .B(n_967), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_967), .B(n_1011), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_961), .A2(n_946), .B1(n_965), .B2(n_996), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1011), .B(n_999), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_976), .Y(n_1044) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_1011), .B(n_964), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_999), .B(n_970), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_970), .B(n_984), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_1013), .B(n_998), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_968), .B(n_952), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_988), .A2(n_980), .B1(n_966), .B2(n_941), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_980), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_978), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_996), .A2(n_988), .B1(n_968), .B2(n_1000), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_968), .B(n_952), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_968), .B(n_943), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_968), .B(n_945), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_941), .B(n_949), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_945), .B(n_962), .Y(n_1058) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_953), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_969), .A2(n_995), .B1(n_975), .B2(n_987), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_941), .B(n_949), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_960), .B(n_962), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_941), .A2(n_949), .B1(n_1006), .B2(n_951), .Y(n_1063) );
NAND2xp5_ASAP7_75t_SL g1064 ( .A(n_1010), .B(n_997), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1003), .B(n_969), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1066 ( .A(n_977), .B(n_940), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_974), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_991), .B(n_992), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_944), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1003), .B(n_985), .Y(n_1070) );
INVx1_ASAP7_75t_SL g1071 ( .A(n_971), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_979), .B(n_985), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1041), .B(n_1020), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1074 ( .A(n_1020), .B(n_940), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1031), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1031), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1041), .B(n_940), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1043), .B(n_947), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1043), .B(n_947), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_1042), .A2(n_1002), .B1(n_1017), .B2(n_1001), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1065), .B(n_947), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1037), .Y(n_1082) );
INVx3_ASAP7_75t_L g1083 ( .A(n_1039), .Y(n_1083) );
NAND2xp5_ASAP7_75t_SL g1084 ( .A(n_1069), .B(n_1017), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1025), .B(n_1003), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1025), .B(n_1004), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_1052), .Y(n_1087) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_1028), .B(n_1009), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1022), .B(n_939), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1062), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1055), .B(n_983), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1055), .B(n_983), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1056), .B(n_983), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1046), .B(n_939), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1033), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1046), .B(n_939), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1056), .B(n_983), .Y(n_1097) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_1021), .B(n_1016), .C(n_1007), .Y(n_1098) );
CKINVDCx16_ASAP7_75t_R g1099 ( .A(n_1038), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1070), .B(n_1015), .Y(n_1100) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_1045), .B(n_972), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1070), .B(n_1015), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1062), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1047), .B(n_1015), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1033), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1047), .B(n_1015), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1049), .B(n_989), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1049), .B(n_989), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1054), .B(n_989), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_1024), .A2(n_956), .B1(n_1007), .B2(n_1008), .Y(n_1110) );
NAND2x1p5_ASAP7_75t_L g1111 ( .A(n_1035), .B(n_956), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1079), .B(n_1045), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1079), .B(n_1040), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1090), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1103), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1079), .B(n_1040), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1086), .B(n_1029), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1086), .B(n_1044), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1078), .B(n_1034), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1075), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1078), .B(n_1034), .Y(n_1121) );
INVx2_ASAP7_75t_SL g1122 ( .A(n_1099), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1099), .B(n_1048), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1075), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1076), .Y(n_1125) );
INVxp67_ASAP7_75t_L g1126 ( .A(n_1087), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1082), .Y(n_1127) );
INVx6_ASAP7_75t_L g1128 ( .A(n_1088), .Y(n_1128) );
INVx1_ASAP7_75t_SL g1129 ( .A(n_1073), .Y(n_1129) );
NOR2xp67_ASAP7_75t_L g1130 ( .A(n_1098), .B(n_1018), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1074), .B(n_1023), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1104), .B(n_1036), .Y(n_1132) );
INVx1_ASAP7_75t_SL g1133 ( .A(n_1073), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1104), .B(n_1067), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1106), .B(n_1058), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1077), .B(n_1034), .Y(n_1136) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_1098), .B(n_1059), .C(n_1053), .Y(n_1137) );
BUFx2_ASAP7_75t_L g1138 ( .A(n_1087), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1095), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1087), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1106), .B(n_1058), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1077), .B(n_1066), .Y(n_1142) );
NOR3xp33_ASAP7_75t_L g1143 ( .A(n_1080), .B(n_1027), .C(n_1050), .Y(n_1143) );
INVx1_ASAP7_75t_SL g1144 ( .A(n_1084), .Y(n_1144) );
NAND2x1_ASAP7_75t_L g1145 ( .A(n_1110), .B(n_1035), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1081), .B(n_1066), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1105), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1105), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1094), .B(n_1026), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1120), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1127), .Y(n_1151) );
OAI221xp5_ASAP7_75t_SL g1152 ( .A1(n_1143), .A2(n_1060), .B1(n_1072), .B2(n_1085), .C(n_1074), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1114), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1113), .B(n_1081), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1113), .B(n_1100), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1116), .B(n_1100), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1116), .B(n_1100), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1120), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1124), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1142), .B(n_1102), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1142), .B(n_1102), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1124), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1129), .B(n_1089), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_1140), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_1137), .A2(n_1080), .B1(n_1101), .B2(n_1108), .Y(n_1165) );
INVx2_ASAP7_75t_SL g1166 ( .A(n_1122), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1115), .B(n_1102), .Y(n_1167) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_1130), .A2(n_1096), .B1(n_1094), .B2(n_1085), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1125), .Y(n_1169) );
AOI222xp33_ASAP7_75t_L g1170 ( .A1(n_1136), .A2(n_1092), .B1(n_1097), .B2(n_1091), .C1(n_1093), .C2(n_1108), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1138), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1146), .B(n_1091), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1133), .B(n_1089), .Y(n_1173) );
AOI211xp5_ASAP7_75t_L g1174 ( .A1(n_1122), .A2(n_1063), .B(n_1071), .C(n_1032), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1123), .A2(n_1030), .B1(n_1038), .B2(n_1069), .Y(n_1175) );
O2A1O1Ixp33_ASAP7_75t_L g1176 ( .A1(n_1134), .A2(n_1064), .B(n_1008), .C(n_1068), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1125), .Y(n_1177) );
INVxp67_ASAP7_75t_SL g1178 ( .A(n_1138), .Y(n_1178) );
INVx2_ASAP7_75t_SL g1179 ( .A(n_1166), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1150), .Y(n_1180) );
NAND3xp33_ASAP7_75t_SL g1181 ( .A(n_1174), .B(n_1145), .C(n_1144), .Y(n_1181) );
NAND2x1p5_ASAP7_75t_L g1182 ( .A(n_1166), .B(n_971), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1150), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1158), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1158), .Y(n_1185) );
NAND2xp5_ASAP7_75t_SL g1186 ( .A(n_1175), .B(n_1126), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1170), .B(n_1119), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1153), .B(n_1117), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_1163), .B(n_1131), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_1152), .A2(n_1119), .B1(n_1121), .B2(n_1136), .C(n_1118), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1164), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1159), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1159), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1172), .B(n_1121), .Y(n_1194) );
INVxp67_ASAP7_75t_L g1195 ( .A(n_1171), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1163), .B(n_1131), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1151), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1172), .B(n_1146), .Y(n_1198) );
NOR2xp33_ASAP7_75t_SL g1199 ( .A(n_1182), .B(n_1178), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_1190), .A2(n_1168), .B1(n_1165), .B2(n_1167), .Y(n_1200) );
AOI21xp33_ASAP7_75t_L g1201 ( .A1(n_1190), .A2(n_1176), .B(n_1145), .Y(n_1201) );
OAI322xp33_ASAP7_75t_L g1202 ( .A1(n_1187), .A2(n_1173), .A3(n_1160), .B1(n_1161), .B2(n_1157), .C1(n_1156), .C2(n_1155), .Y(n_1202) );
NOR2xp33_ASAP7_75t_SL g1203 ( .A(n_1182), .B(n_1181), .Y(n_1203) );
OAI21xp5_ASAP7_75t_L g1204 ( .A1(n_1181), .A2(n_1154), .B(n_1173), .Y(n_1204) );
OAI32xp33_ASAP7_75t_L g1205 ( .A1(n_1191), .A2(n_1154), .A3(n_1132), .B1(n_1149), .B2(n_1141), .Y(n_1205) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_1186), .A2(n_1128), .B1(n_1101), .B2(n_1112), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_1195), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1180), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1179), .B(n_1112), .Y(n_1209) );
INVxp67_ASAP7_75t_L g1210 ( .A(n_1188), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_1195), .A2(n_1101), .B1(n_1109), .B2(n_1108), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1202), .A2(n_1192), .B1(n_1184), .B2(n_1185), .C(n_1183), .Y(n_1212) );
AOI222xp33_ASAP7_75t_L g1213 ( .A1(n_1204), .A2(n_1193), .B1(n_1194), .B2(n_1198), .C1(n_1017), .C2(n_1169), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1207), .Y(n_1214) );
OAI21xp5_ASAP7_75t_L g1215 ( .A1(n_1203), .A2(n_1196), .B(n_1189), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1200), .A2(n_1101), .B1(n_1128), .B2(n_1107), .Y(n_1216) );
AOI21xp33_ASAP7_75t_L g1217 ( .A1(n_1207), .A2(n_1083), .B(n_1026), .Y(n_1217) );
NAND4xp25_ASAP7_75t_L g1218 ( .A(n_1201), .B(n_1001), .C(n_971), .D(n_1101), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_1206), .A2(n_1030), .B1(n_1128), .B2(n_1135), .Y(n_1219) );
AOI221x1_ASAP7_75t_L g1220 ( .A1(n_1208), .A2(n_1162), .B1(n_1177), .B2(n_1083), .C(n_1197), .Y(n_1220) );
NAND5xp2_ASAP7_75t_L g1221 ( .A(n_1213), .B(n_1199), .C(n_1211), .D(n_1111), .E(n_1210), .Y(n_1221) );
AND4x1_ASAP7_75t_L g1222 ( .A(n_1215), .B(n_1211), .C(n_1017), .D(n_1209), .Y(n_1222) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1214), .B(n_1205), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1218), .Y(n_1224) );
NOR2x1_ASAP7_75t_L g1225 ( .A(n_1219), .B(n_1001), .Y(n_1225) );
CKINVDCx16_ASAP7_75t_R g1226 ( .A(n_1216), .Y(n_1226) );
INVx5_ASAP7_75t_L g1227 ( .A(n_1226), .Y(n_1227) );
NAND4xp75_ASAP7_75t_L g1228 ( .A(n_1225), .B(n_1212), .C(n_1220), .D(n_1217), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1224), .Y(n_1229) );
NAND5xp2_ASAP7_75t_L g1230 ( .A(n_1223), .B(n_1111), .C(n_1017), .D(n_1109), .E(n_1107), .Y(n_1230) );
NOR3xp33_ASAP7_75t_L g1231 ( .A(n_1229), .B(n_1221), .C(n_1222), .Y(n_1231) );
OAI22xp5_ASAP7_75t_SL g1232 ( .A1(n_1227), .A2(n_1051), .B1(n_1019), .B2(n_1111), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1233 ( .A1(n_1231), .A2(n_1227), .B1(n_1228), .B2(n_1230), .C(n_1019), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1232), .Y(n_1234) );
INVx5_ASAP7_75t_L g1235 ( .A(n_1234), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_1233), .A2(n_1128), .B1(n_1177), .B2(n_1162), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1235), .Y(n_1237) );
AOI222xp33_ASAP7_75t_L g1238 ( .A1(n_1237), .A2(n_1236), .B1(n_1083), .B2(n_1148), .C1(n_1139), .C2(n_1147), .Y(n_1238) );
AOI22xp5_ASAP7_75t_L g1239 ( .A1(n_1238), .A2(n_1057), .B1(n_1061), .B2(n_1107), .Y(n_1239) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_1239), .A2(n_1092), .B1(n_1093), .B2(n_1097), .Y(n_1240) );
endmodule