module fake_jpeg_24929_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_1),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_23),
.B1(n_18),
.B2(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_42),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_16),
.C(n_28),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_51),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_16),
.B(n_28),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_34),
.B(n_29),
.C(n_27),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_26),
.B1(n_20),
.B2(n_33),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_26),
.B1(n_23),
.B2(n_35),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_64),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_33),
.B1(n_53),
.B2(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_17),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_36),
.B1(n_33),
.B2(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_72),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_43),
.B1(n_25),
.B2(n_53),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_81),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_40),
.B(n_34),
.C(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_36),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_40),
.C(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_91),
.B1(n_75),
.B2(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_64),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_69),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_92),
.B(n_102),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_38),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_62),
.B1(n_81),
.B2(n_61),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_38),
.B(n_35),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_38),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_3),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_4),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_91),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_111),
.B1(n_124),
.B2(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_121),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_58),
.B1(n_52),
.B2(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_58),
.B1(n_25),
.B2(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_30),
.B1(n_24),
.B2(n_22),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_78),
.B1(n_39),
.B2(n_32),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_80),
.B1(n_32),
.B2(n_39),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_13),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_14),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_3),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_94),
.C(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_11),
.B1(n_12),
.B2(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_105),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_7),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_101),
.C(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_98),
.B1(n_113),
.B2(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_138),
.B(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_115),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_146),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_120),
.C(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_120),
.C(n_112),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_135),
.C(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_117),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_154),
.B(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_139),
.C(n_130),
.Y(n_156)
);

OAI322xp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_121),
.A3(n_128),
.B1(n_124),
.B2(n_104),
.C1(n_92),
.C2(n_101),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_137),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_160),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_139),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_89),
.B(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_87),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_170),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_152),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_173),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_151),
.C(n_125),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_159),
.B1(n_135),
.B2(n_145),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_179),
.B(n_182),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_149),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_145),
.B1(n_136),
.B2(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_154),
.B1(n_162),
.B2(n_136),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_183),
.C(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_162),
.B1(n_160),
.B2(n_151),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g186 ( 
.A(n_183),
.B(n_172),
.CI(n_166),
.CON(n_186),
.SN(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.C(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_167),
.C(n_107),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_170),
.B(n_121),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_177),
.C(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_195),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_185),
.B1(n_184),
.B2(n_187),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_191),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_190),
.Y(n_198)
);

AOI311xp33_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_193),
.A3(n_107),
.B(n_9),
.C(n_8),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_200),
.A3(n_198),
.B1(n_197),
.B2(n_9),
.C1(n_8),
.C2(n_97),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_97),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_9),
.Y(n_203)
);


endmodule