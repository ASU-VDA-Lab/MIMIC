module fake_jpeg_14525_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_14),
.B1(n_9),
.B2(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_20),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_21),
.B2(n_23),
.Y(n_31)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_37),
.B(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_18),
.B1(n_22),
.B2(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_22),
.B1(n_20),
.B2(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_42),
.B1(n_23),
.B2(n_37),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_24),
.C(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_34),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_41),
.B(n_39),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_44),
.B(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_46),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_6),
.B2(n_49),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_0),
.C(n_49),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_0),
.Y(n_54)
);


endmodule