module fake_aes_8110_n_723 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_723);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_723;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_51), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_2), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_26), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_57), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_33), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_70), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_24), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_66), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_21), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_32), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_27), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_75), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_30), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_73), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_9), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_8), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_56), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_76), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_42), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_60), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_67), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_50), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_28), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_45), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_22), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_4), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_69), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_8), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_49), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_12), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_38), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_20), .Y(n_124) );
INVxp33_ASAP7_75t_SL g125 ( .A(n_17), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_95), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_91), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_127), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_82), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_109), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_111), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_123), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_84), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_103), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_88), .B(n_36), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_88), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_127), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_105), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_101), .B(n_0), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_97), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_93), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_99), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_98), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_99), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_106), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_79), .B(n_1), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_106), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_79), .B(n_1), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_102), .B(n_2), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_85), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_81), .B(n_3), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_161), .B(n_129), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_133), .B(n_113), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_133), .B(n_81), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_133), .B(n_90), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_131), .A2(n_125), .B1(n_116), .B2(n_117), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_115), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_161), .A2(n_108), .B1(n_87), .B2(n_120), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_147), .B(n_107), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_136), .B(n_96), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_130), .B(n_121), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_141), .B(n_98), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_138), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_141), .B(n_83), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_130), .Y(n_198) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_150), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_158), .B(n_83), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_120), .B1(n_87), .B2(n_117), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_142), .B(n_119), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_142), .B(n_144), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_129), .A2(n_126), .B1(n_119), .B2(n_114), .Y(n_208) );
INVx4_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_150), .B(n_112), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
INVxp67_ASAP7_75t_L g214 ( .A(n_143), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
INVxp33_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_138), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_159), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_144), .B(n_110), .Y(n_222) );
BUFx10_ASAP7_75t_L g223 ( .A(n_171), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_146), .B(n_86), .Y(n_224) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_145), .B(n_94), .Y(n_225) );
AO22x2_ASAP7_75t_L g226 ( .A1(n_146), .A2(n_126), .B1(n_114), .B2(n_113), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_151), .B(n_104), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_151), .A2(n_112), .B1(n_108), .B2(n_100), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_138), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_153), .Y(n_230) );
NAND3xp33_ASAP7_75t_L g231 ( .A(n_153), .B(n_100), .C(n_4), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_135), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_155), .B(n_3), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_155), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_156), .B(n_6), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g237 ( .A(n_167), .B(n_7), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_165), .B(n_10), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_166), .B(n_11), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_219), .B(n_139), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_178), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_234), .A2(n_166), .B(n_168), .C(n_169), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_229), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_178), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_178), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_229), .Y(n_249) );
INVxp67_ASAP7_75t_SL g250 ( .A(n_199), .Y(n_250) );
NOR3xp33_ASAP7_75t_SL g251 ( .A(n_182), .B(n_172), .C(n_169), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_230), .B(n_168), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_180), .B(n_172), .Y(n_255) );
INVx4_ASAP7_75t_L g256 ( .A(n_178), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_206), .B(n_167), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_206), .B(n_170), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_180), .B(n_237), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_180), .B(n_163), .Y(n_261) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_233), .B(n_164), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_206), .B(n_224), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_217), .B(n_164), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_239), .A2(n_164), .B(n_163), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_217), .B(n_145), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_239), .Y(n_272) );
OAI21xp33_ASAP7_75t_SL g273 ( .A1(n_176), .A2(n_164), .B(n_163), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_181), .B(n_145), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_233), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_176), .A2(n_140), .B1(n_145), .B2(n_148), .Y(n_277) );
BUFx4f_ASAP7_75t_L g278 ( .A(n_204), .Y(n_278) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_183), .B(n_163), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_209), .Y(n_280) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_223), .B(n_148), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_177), .B(n_148), .Y(n_282) );
CKINVDCx8_ASAP7_75t_R g283 ( .A(n_204), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_192), .B(n_148), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_233), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_192), .B(n_145), .Y(n_286) );
NOR3xp33_ASAP7_75t_SL g287 ( .A(n_188), .B(n_11), .C(n_13), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_185), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_208), .A2(n_145), .B1(n_149), .B2(n_157), .Y(n_289) );
NAND2xp33_ASAP7_75t_SL g290 ( .A(n_209), .B(n_152), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_200), .B(n_13), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_204), .Y(n_292) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_198), .Y(n_293) );
AND3x1_ASAP7_75t_SL g294 ( .A(n_203), .B(n_15), .C(n_16), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_190), .B(n_157), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_226), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_189), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_200), .B(n_16), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_185), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_226), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_195), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_226), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_193), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_223), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_191), .B(n_157), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_201), .B(n_149), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_202), .B(n_149), .Y(n_308) );
NOR2xp33_ASAP7_75t_R g309 ( .A(n_223), .B(n_47), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_204), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_196), .A2(n_137), .B1(n_132), .B2(n_152), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_208), .B(n_17), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_256), .B(n_195), .Y(n_314) );
BUFx10_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_305), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_241), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_262), .A2(n_208), .B1(n_214), .B2(n_240), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_309), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_298), .B(n_232), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_256), .B(n_195), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_256), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_255), .B(n_196), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_242), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_262), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_291), .B(n_240), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_250), .B(n_228), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_275), .A2(n_225), .B(n_195), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_264), .B(n_208), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_268), .B(n_238), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_301), .A2(n_204), .B1(n_227), .B2(n_235), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_255), .B(n_238), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_255), .B(n_236), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_262), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_266), .Y(n_337) );
BUFx2_ASAP7_75t_SL g338 ( .A(n_283), .Y(n_338) );
AND2x6_ASAP7_75t_L g339 ( .A(n_242), .B(n_204), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_291), .B(n_222), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_291), .B(n_195), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_301), .A2(n_231), .B1(n_194), .B2(n_227), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_269), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_269), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_260), .B(n_194), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_257), .B(n_227), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_278), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_245), .B(n_227), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_285), .A2(n_227), .B1(n_174), .B2(n_179), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_292), .Y(n_351) );
CKINVDCx8_ASAP7_75t_R g352 ( .A(n_299), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_272), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_271), .A2(n_174), .B(n_187), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_245), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_278), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_299), .B(n_227), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_299), .B(n_18), .Y(n_359) );
INVx3_ASAP7_75t_SL g360 ( .A(n_281), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_310), .B(n_18), .Y(n_361) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_284), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_248), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_246), .B(n_247), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_252), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_274), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_252), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_276), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_267), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_315), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_251), .B1(n_284), .B2(n_263), .C(n_282), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_327), .A2(n_277), .B1(n_260), .B2(n_313), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_283), .B1(n_276), .B2(n_258), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_352), .A2(n_273), .B(n_287), .C(n_279), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_327), .A2(n_260), .B1(n_313), .B2(n_286), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_334), .B(n_293), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
CKINVDCx6p67_ASAP7_75t_R g380 ( .A(n_360), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_329), .A2(n_285), .B(n_276), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_327), .A2(n_286), .B1(n_295), .B2(n_297), .Y(n_382) );
AO31x2_ASAP7_75t_L g383 ( .A1(n_319), .A2(n_295), .A3(n_297), .B(n_303), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_334), .B(n_284), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_327), .A2(n_303), .B1(n_294), .B2(n_261), .Y(n_386) );
AOI211xp5_ASAP7_75t_L g387 ( .A1(n_321), .A2(n_282), .B(n_243), .C(n_261), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_316), .Y(n_388) );
CKINVDCx8_ASAP7_75t_R g389 ( .A(n_318), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_317), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_358), .A2(n_270), .B1(n_286), .B2(n_246), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_347), .A2(n_289), .B(n_265), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_355), .A2(n_253), .B(n_259), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_330), .A2(n_261), .B1(n_282), .B2(n_270), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_359), .A2(n_278), .B1(n_247), .B2(n_311), .Y(n_395) );
CKINVDCx6p67_ASAP7_75t_R g396 ( .A(n_360), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_324), .B(n_259), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_358), .A2(n_311), .B1(n_292), .B2(n_249), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_335), .B(n_249), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_265), .B1(n_292), .B2(n_249), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_337), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_358), .A2(n_312), .B1(n_296), .B2(n_244), .Y(n_403) );
OAI21xp33_ASAP7_75t_SL g404 ( .A1(n_377), .A2(n_345), .B(n_343), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_337), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_386), .A2(n_330), .B1(n_344), .B2(n_328), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_390), .B(n_344), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_383), .B(n_336), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
HB1xp67_ASAP7_75t_SL g411 ( .A(n_389), .Y(n_411) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_386), .A2(n_361), .A3(n_331), .B1(n_340), .B2(n_318), .C1(n_369), .C2(n_358), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_372), .A2(n_354), .B1(n_367), .B2(n_365), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_390), .B(n_354), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_376), .A2(n_367), .B1(n_363), .B2(n_365), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_402), .B(n_335), .Y(n_416) );
OA21x2_ASAP7_75t_L g417 ( .A1(n_381), .A2(n_343), .B(n_345), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_371), .A2(n_361), .B1(n_328), .B2(n_340), .C(n_346), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_402), .B(n_336), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
NOR2x1_ASAP7_75t_L g422 ( .A(n_374), .B(n_348), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_320), .B(n_333), .C(n_326), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_384), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_378), .A2(n_362), .B1(n_326), .B2(n_341), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_378), .A2(n_362), .B1(n_341), .B2(n_368), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_399), .B(n_315), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_397), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_385), .A2(n_368), .B1(n_315), .B2(n_320), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_370), .B(n_360), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_410), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_411), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_406), .A2(n_388), .B1(n_399), .B2(n_382), .C(n_394), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_405), .B(n_383), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_413), .A2(n_392), .B(n_400), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_412), .B(n_306), .C(n_403), .D(n_393), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_410), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_432), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_412), .A2(n_395), .B(n_403), .C(n_391), .Y(n_443) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_370), .B1(n_396), .B2(n_380), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_420), .B(n_383), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_430), .A2(n_373), .B1(n_396), .B2(n_380), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_420), .B(n_383), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_430), .B(n_383), .Y(n_448) );
NOR2xp33_ASAP7_75t_R g449 ( .A(n_411), .B(n_389), .Y(n_449) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_409), .B(n_379), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_432), .Y(n_451) );
AOI33xp33_ASAP7_75t_L g452 ( .A1(n_426), .A2(n_137), .A3(n_215), .B1(n_187), .B2(n_184), .B3(n_179), .Y(n_452) );
OAI222xp33_ASAP7_75t_L g453 ( .A1(n_408), .A2(n_398), .B1(n_379), .B2(n_349), .C1(n_350), .C2(n_364), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_419), .A2(n_315), .B1(n_342), .B2(n_338), .Y(n_455) );
NAND2xp33_ASAP7_75t_SL g456 ( .A(n_408), .B(n_348), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_350), .B(n_137), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_308), .B1(n_307), .B2(n_254), .C(n_244), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_416), .A2(n_254), .B1(n_290), .B2(n_339), .C1(n_348), .C2(n_357), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_426), .A2(n_290), .B1(n_349), .B2(n_366), .C(n_332), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_423), .B(n_215), .C(n_184), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_19), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_418), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_416), .B(n_366), .Y(n_465) );
OAI33xp33_ASAP7_75t_L g466 ( .A1(n_415), .A2(n_207), .A3(n_213), .B1(n_211), .B2(n_197), .B3(n_193), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_423), .A2(n_213), .B(n_197), .C(n_211), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_418), .Y(n_468) );
OAI33xp33_ASAP7_75t_L g469 ( .A1(n_415), .A2(n_205), .A3(n_207), .B1(n_220), .B2(n_221), .B3(n_19), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
OAI21x1_ASAP7_75t_L g472 ( .A1(n_450), .A2(n_417), .B(n_422), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_463), .B(n_416), .Y(n_473) );
AOI322xp5_ASAP7_75t_L g474 ( .A1(n_444), .A2(n_427), .A3(n_431), .B1(n_405), .B2(n_407), .C1(n_414), .C2(n_422), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g475 ( .A1(n_446), .A2(n_431), .B(n_427), .Y(n_475) );
AOI33xp33_ASAP7_75t_L g476 ( .A1(n_463), .A2(n_445), .A3(n_447), .B1(n_437), .B2(n_436), .B3(n_405), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_437), .B(n_408), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_448), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_470), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_468), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_465), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_445), .B(n_407), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_447), .B(n_428), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_469), .A2(n_407), .B1(n_414), .B2(n_404), .C(n_429), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_442), .B(n_414), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_458), .B(n_425), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_470), .B(n_425), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_456), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_449), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_452), .B(n_428), .C(n_421), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_442), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_470), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_433), .B(n_425), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_433), .B(n_424), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_451), .B(n_424), .Y(n_503) );
OAI21xp5_ASAP7_75t_SL g504 ( .A1(n_435), .A2(n_429), .B(n_421), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_440), .B(n_424), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_440), .B(n_421), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_441), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_453), .B(n_429), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_441), .B(n_421), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_443), .B(n_421), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_456), .B(n_417), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_439), .B(n_21), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_455), .A2(n_349), .B1(n_351), .B2(n_332), .C(n_366), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_439), .B(n_22), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_450), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_438), .B(n_457), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_457), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_457), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_438), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_455), .B(n_417), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_493), .B(n_462), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_484), .B(n_23), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_495), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_483), .B(n_459), .Y(n_527) );
AND2x4_ASAP7_75t_SL g528 ( .A(n_485), .B(n_357), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_487), .B(n_23), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_471), .B(n_25), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_485), .B(n_417), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_488), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_485), .B(n_461), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_475), .B(n_466), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_467), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_477), .B(n_205), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_476), .B(n_221), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_503), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_473), .B(n_29), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_501), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_479), .B(n_220), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_479), .B(n_31), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_492), .B(n_34), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_480), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_516), .B(n_514), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_480), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_492), .B(n_35), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_494), .B(n_357), .C(n_351), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_510), .B(n_37), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_518), .B(n_39), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_474), .B(n_40), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_478), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_507), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_518), .B(n_41), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_488), .B(n_43), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_482), .B(n_44), .Y(n_557) );
AND4x1_ASAP7_75t_L g558 ( .A(n_486), .B(n_338), .C(n_48), .D(n_52), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_482), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_497), .B(n_46), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_497), .B(n_54), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_58), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_500), .B(n_59), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_478), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_512), .B(n_61), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_505), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_489), .B(n_62), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_504), .B(n_64), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_478), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_523), .B(n_65), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_489), .B(n_490), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_523), .B(n_68), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_506), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_506), .Y(n_575) );
INVx3_ASAP7_75t_SL g576 ( .A(n_506), .Y(n_576) );
NAND2xp33_ASAP7_75t_L g577 ( .A(n_522), .B(n_339), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_481), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_521), .B(n_77), .Y(n_579) );
NAND2xp33_ASAP7_75t_R g580 ( .A(n_513), .B(n_502), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_502), .B(n_78), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_366), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_545), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_535), .A2(n_522), .B(n_472), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_546), .B(n_522), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_539), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_522), .B1(n_508), .B2(n_511), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_572), .B(n_511), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_530), .B(n_522), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_529), .B(n_520), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_544), .B(n_513), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_576), .B(n_481), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_541), .B(n_520), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_525), .A2(n_515), .B(n_517), .C(n_519), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_559), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_536), .A2(n_517), .B1(n_496), .B2(n_519), .Y(n_599) );
OAI22xp33_ASAP7_75t_SL g600 ( .A1(n_576), .A2(n_507), .B1(n_496), .B2(n_491), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_569), .A2(n_472), .B(n_491), .C(n_509), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_563), .Y(n_602) );
OAI32xp33_ASAP7_75t_L g603 ( .A1(n_580), .A2(n_507), .A3(n_491), .B1(n_509), .B2(n_498), .Y(n_603) );
OAI21xp33_ASAP7_75t_SL g604 ( .A1(n_570), .A2(n_498), .B(n_349), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_577), .A2(n_332), .B1(n_349), .B2(n_357), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_567), .B(n_173), .Y(n_606) );
NOR2xp67_ASAP7_75t_L g607 ( .A(n_554), .B(n_173), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_538), .A2(n_527), .B1(n_552), .B2(n_550), .C(n_574), .Y(n_608) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_524), .B(n_339), .Y(n_609) );
A2O1A1Ixp33_ASAP7_75t_L g610 ( .A1(n_569), .A2(n_323), .B(n_356), .C(n_325), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_577), .A2(n_323), .B(n_356), .C(n_325), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_528), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_532), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_534), .B(n_173), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_550), .A2(n_173), .B(n_175), .C(n_186), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_536), .A2(n_332), .B1(n_339), .B2(n_351), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_575), .B(n_173), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_537), .B(n_175), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_537), .A2(n_175), .B1(n_186), .B2(n_210), .C(n_300), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_551), .B(n_175), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_528), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_578), .Y(n_624) );
NOR2x1p5_ASAP7_75t_L g625 ( .A(n_554), .B(n_323), .Y(n_625) );
NAND2xp33_ASAP7_75t_SL g626 ( .A(n_580), .B(n_339), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_544), .A2(n_364), .B(n_322), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_571), .A2(n_339), .B1(n_175), .B2(n_186), .C1(n_210), .C2(n_288), .Y(n_628) );
NAND3xp33_ASAP7_75t_SL g629 ( .A(n_558), .B(n_322), .C(n_314), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_566), .A2(n_186), .B1(n_210), .B2(n_300), .C(n_288), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_565), .B(n_186), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_544), .A2(n_364), .B1(n_314), .B2(n_322), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_555), .B(n_210), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_578), .Y(n_634) );
OAI322xp33_ASAP7_75t_L g635 ( .A1(n_588), .A2(n_540), .A3(n_557), .B1(n_582), .B2(n_543), .C1(n_553), .C2(n_542), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_586), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_613), .B(n_560), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_613), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_585), .B(n_573), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_585), .B(n_573), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_598), .Y(n_643) );
NOR4xp25_ASAP7_75t_SL g644 ( .A(n_626), .B(n_548), .C(n_549), .D(n_531), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_593), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_589), .B(n_562), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_602), .B(n_548), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_612), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_594), .A2(n_564), .B(n_561), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_592), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_596), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_624), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_625), .B(n_548), .Y(n_653) );
XNOR2xp5_ASAP7_75t_L g654 ( .A(n_623), .B(n_564), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_595), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_622), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_621), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_614), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_607), .Y(n_660) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_584), .B(n_531), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_614), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_599), .B(n_531), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_591), .B(n_561), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_591), .B(n_560), .Y(n_665) );
NOR3xp33_ASAP7_75t_SL g666 ( .A(n_629), .B(n_581), .C(n_556), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_618), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_636), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_644), .A2(n_603), .B(n_604), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_659), .A2(n_597), .B(n_608), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_654), .A2(n_594), .B1(n_605), .B2(n_601), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_646), .A2(n_605), .B1(n_601), .B2(n_632), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_649), .A2(n_587), .B1(n_609), .B2(n_616), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_639), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_641), .A2(n_616), .B1(n_600), .B2(n_628), .Y(n_676) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_648), .B(n_627), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_643), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_640), .B(n_606), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_650), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_651), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_645), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g683 ( .A1(n_653), .A2(n_610), .B(n_619), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_661), .A2(n_615), .B(n_620), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_652), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_656), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_666), .A2(n_611), .B(n_633), .C(n_630), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_666), .A2(n_568), .B1(n_579), .B2(n_617), .C(n_631), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_645), .Y(n_689) );
OA22x2_ASAP7_75t_L g690 ( .A1(n_677), .A2(n_657), .B1(n_660), .B2(n_663), .Y(n_690) );
NOR2x1p5_ASAP7_75t_L g691 ( .A(n_679), .B(n_663), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_680), .B(n_662), .Y(n_692) );
OAI321xp33_ASAP7_75t_L g693 ( .A1(n_671), .A2(n_642), .A3(n_641), .B1(n_665), .B2(n_664), .C(n_647), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_670), .A2(n_660), .B(n_657), .C(n_642), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_681), .B(n_655), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_672), .A2(n_658), .B(n_667), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_685), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_682), .B(n_637), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_689), .B(n_635), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_669), .A2(n_210), .B(n_339), .C(n_280), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_674), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_669), .A2(n_304), .B(n_280), .C(n_302), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_675), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_678), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_687), .B(n_302), .C(n_364), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_673), .A2(n_314), .B1(n_676), .B2(n_684), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_683), .A2(n_687), .B(n_668), .C(n_684), .Y(n_707) );
OAI221xp5_ASAP7_75t_SL g708 ( .A1(n_688), .A2(n_649), .B1(n_676), .B2(n_673), .C(n_669), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_686), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_709), .B(n_706), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_707), .B(n_696), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_699), .Y(n_712) );
AOI221x1_ASAP7_75t_L g713 ( .A1(n_705), .A2(n_704), .B1(n_703), .B2(n_701), .C(n_697), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_690), .Y(n_714) );
NOR2xp67_ASAP7_75t_L g715 ( .A(n_710), .B(n_694), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_711), .B(n_708), .C(n_693), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_712), .A2(n_693), .B(n_690), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_716), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_715), .A2(n_712), .B1(n_717), .B2(n_714), .Y(n_719) );
OR3x1_ASAP7_75t_L g720 ( .A(n_718), .B(n_713), .C(n_702), .Y(n_720) );
INVx3_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_700), .B1(n_692), .B2(n_691), .C1(n_695), .C2(n_698), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_721), .B(n_720), .Y(n_723) );
endmodule