module fake_jpeg_16064_n_357 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_357);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_12),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_39),
.B(n_49),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_55),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_56),
.Y(n_115)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_58),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_14),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_16),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_22),
.B1(n_14),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_71),
.A2(n_75),
.B1(n_77),
.B2(n_88),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_74),
.B(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_47),
.B1(n_41),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_108),
.B1(n_13),
.B2(n_29),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_14),
.B1(n_20),
.B2(n_22),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_20),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_79),
.A2(n_82),
.B(n_0),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_98),
.B1(n_103),
.B2(n_2),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_14),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_112),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_14),
.B1(n_20),
.B2(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_28),
.B1(n_35),
.B2(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_20),
.B1(n_35),
.B2(n_31),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_104),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_36),
.B1(n_30),
.B2(n_18),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_30),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_29),
.C(n_13),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_18),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_37),
.B(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_37),
.B(n_29),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_117),
.B(n_142),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_16),
.B1(n_13),
.B2(n_29),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_125),
.B1(n_143),
.B2(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_158),
.B1(n_100),
.B2(n_132),
.Y(n_203)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

OA22x2_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_127),
.A2(n_102),
.B1(n_91),
.B2(n_100),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_150),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_5),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_132),
.A2(n_135),
.B(n_77),
.Y(n_179)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_8),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_89),
.C(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_88),
.A2(n_3),
.B(n_9),
.C(n_10),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_9),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_10),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_151),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_0),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_1),
.B1(n_2),
.B2(n_97),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_155),
.B(n_70),
.Y(n_167)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_157),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_82),
.B(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_2),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_76),
.A2(n_110),
.B1(n_80),
.B2(n_97),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_87),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_115),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_72),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_200),
.B(n_141),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_184),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_121),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_71),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_174),
.B(n_172),
.C(n_179),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_191),
.Y(n_234)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_107),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_115),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_68),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_115),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_186),
.B(n_194),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_123),
.B(n_68),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_196),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_140),
.A2(n_114),
.B1(n_69),
.B2(n_102),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_207),
.B1(n_162),
.B2(n_136),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_69),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_114),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_91),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_126),
.B1(n_120),
.B2(n_154),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_154),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_119),
.B1(n_135),
.B2(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_211),
.A2(n_218),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_163),
.B1(n_135),
.B2(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_221),
.B1(n_223),
.B2(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_220),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_149),
.B(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_137),
.B1(n_127),
.B2(n_117),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_198),
.B(n_174),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_160),
.B1(n_151),
.B2(n_164),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_127),
.B(n_153),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_224),
.A2(n_236),
.B(n_206),
.Y(n_263)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_227),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_244),
.C(n_184),
.Y(n_253)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_206),
.B1(n_207),
.B2(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_189),
.B(n_148),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_122),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_237),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_136),
.B(n_118),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_238),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_242),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_191),
.B(n_128),
.CI(n_159),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_241),
.B(n_200),
.Y(n_271)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_246),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_268),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_255),
.C(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_170),
.C(n_199),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_271),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_199),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_266),
.B(n_274),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_211),
.A2(n_200),
.B1(n_171),
.B2(n_193),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_196),
.B1(n_188),
.B2(n_176),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_200),
.B(n_168),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_192),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_273),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_171),
.B1(n_192),
.B2(n_175),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_212),
.B1(n_210),
.B2(n_240),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_215),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_234),
.A2(n_223),
.B(n_231),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_238),
.B1(n_218),
.B2(n_229),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_276),
.A2(n_283),
.B1(n_287),
.B2(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_230),
.C(n_226),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_282),
.C(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_230),
.C(n_234),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_227),
.B1(n_225),
.B2(n_220),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_269),
.C(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_235),
.C(n_209),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_217),
.B1(n_175),
.B2(n_205),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_247),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_251),
.B(n_166),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_294),
.C(n_297),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_293),
.A2(n_300),
.B1(n_256),
.B2(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_169),
.C(n_176),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_173),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_267),
.B(n_228),
.C(n_188),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_248),
.B(n_268),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_250),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_250),
.A2(n_266),
.B1(n_263),
.B2(n_271),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_300),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_257),
.B1(n_246),
.B2(n_249),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_308),
.B1(n_310),
.B2(n_314),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_256),
.B1(n_260),
.B2(n_264),
.Y(n_308)
);

OAI32xp33_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_261),
.A3(n_258),
.B1(n_270),
.B2(n_254),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_313),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_264),
.B1(n_258),
.B2(n_260),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_316),
.C(n_296),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_317),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_254),
.B(n_259),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_259),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_245),
.B1(n_275),
.B2(n_261),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_288),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_278),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_278),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_292),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_324),
.C(n_326),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_279),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_306),
.B(n_296),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_295),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_331),
.C(n_323),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_299),
.C(n_295),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_287),
.A3(n_283),
.B1(n_277),
.B2(n_245),
.C(n_177),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_332),
.B(n_315),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_317),
.B1(n_307),
.B2(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_335),
.B(n_338),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_314),
.B(n_303),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_340),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_308),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_326),
.B(n_331),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_301),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_324),
.B(n_320),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_337),
.A2(n_321),
.B1(n_330),
.B2(n_314),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_344),
.C(n_348),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_177),
.B(n_190),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_334),
.C(n_336),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_336),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_353),
.C(n_349),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_335),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_354),
.A2(n_345),
.B(n_334),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_341),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_345),
.B1(n_339),
.B2(n_340),
.Y(n_357)
);


endmodule