module fake_jpeg_16568_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_54),
.B1(n_31),
.B2(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_17),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_29),
.B1(n_32),
.B2(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_40),
.B1(n_29),
.B2(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_37),
.B1(n_25),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_17),
.B1(n_32),
.B2(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_24),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_78),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_39),
.B(n_2),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_19),
.B(n_27),
.C(n_37),
.Y(n_88)
);

NAND2x1_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_37),
.Y(n_75)
);

NAND2x1_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_39),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_34),
.B1(n_33),
.B2(n_38),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_58),
.B1(n_63),
.B2(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_39),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_60),
.B(n_72),
.Y(n_119)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_91),
.Y(n_130)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_69),
.B1(n_58),
.B2(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_74),
.B1(n_56),
.B2(n_63),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_127),
.B1(n_67),
.B2(n_39),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_112),
.A2(n_116),
.B1(n_118),
.B2(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_60),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_123),
.B(n_132),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_59),
.B1(n_73),
.B2(n_78),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_93),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_73),
.B1(n_77),
.B2(n_81),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_124),
.B(n_88),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_73),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_62),
.B(n_68),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_64),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_83),
.C(n_66),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_92),
.C(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_33),
.B1(n_34),
.B2(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_84),
.B1(n_101),
.B2(n_104),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_39),
.B1(n_67),
.B2(n_19),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_39),
.B(n_2),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_134),
.B(n_92),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_135),
.B(n_100),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_97),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_142),
.C(n_146),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_106),
.B(n_105),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_149),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_151),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_97),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_86),
.C(n_96),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.C(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_86),
.C(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_107),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_154),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_88),
.B1(n_109),
.B2(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_127),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_84),
.B1(n_93),
.B2(n_39),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_14),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_115),
.B1(n_112),
.B2(n_123),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_172),
.B1(n_178),
.B2(n_179),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_118),
.C(n_110),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_132),
.C(n_114),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_119),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_111),
.C(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_176),
.C(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_111),
.C(n_131),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_131),
.B1(n_128),
.B2(n_121),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_183),
.B(n_152),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_39),
.C(n_28),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_155),
.CI(n_149),
.CON(n_187),
.SN(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_193),
.B(n_198),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_137),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_27),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_158),
.B1(n_5),
.B2(n_8),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_196),
.B1(n_168),
.B2(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_28),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_16),
.C(n_19),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_199),
.C(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_16),
.C(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_11),
.C(n_12),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_164),
.C(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_176),
.C(n_184),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_9),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_212),
.B1(n_214),
.B2(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_201),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_196),
.C(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_189),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_218),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_223),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_224),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_203),
.C(n_202),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_187),
.B(n_186),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_186),
.B1(n_199),
.B2(n_197),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_225),
.B(n_217),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_213),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_210),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_207),
.B(n_209),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_240),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_222),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_230),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_244),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_246),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_248),
.B(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_11),
.Y(n_252)
);


endmodule