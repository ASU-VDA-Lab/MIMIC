module fake_netlist_6_33_n_474 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_474);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_474;

wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_111;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_109;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_402;
wire n_352;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_92;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_406;
wire n_102;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_464;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_277;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_85;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_24),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_31),
.B(n_29),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_22),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_25),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_14),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_37),
.B(n_63),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_27),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_10),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_6),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_44),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_4),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_11),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_16),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_13),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_33),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_17),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_40),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_39),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_23),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_38),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_5),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_66),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_78),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_18),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_26),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_19),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_3),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_3),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_115),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_91),
.A2(n_6),
.B(n_7),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_7),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_99),
.B(n_147),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_28),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx8_ASAP7_75t_R g180 ( 
.A(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_94),
.B(n_9),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_12),
.B(n_13),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_96),
.B(n_21),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_128),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_12),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_102),
.B(n_32),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_35),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_109),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_41),
.B(n_58),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_150),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_70),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_151),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_176),
.B(n_85),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_159),
.Y(n_225)
);

CKINVDCx6p67_ASAP7_75t_R g226 ( 
.A(n_183),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_87),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_88),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_200),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_92),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_190),
.B(n_93),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_139),
.B1(n_135),
.B2(n_122),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_198),
.B(n_95),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_97),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g250 ( 
.A1(n_165),
.A2(n_107),
.B(n_100),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_180),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_168),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_178),
.B(n_108),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_111),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_166),
.B(n_211),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_196),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_196),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_216),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_174),
.C(n_201),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_216),
.B1(n_201),
.B2(n_186),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_226),
.B(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_202),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_202),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_172),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_212),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_250),
.A2(n_173),
.B1(n_195),
.B2(n_208),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_222),
.A2(n_203),
.B(n_162),
.C(n_181),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_201),
.C(n_169),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_114),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_251),
.B(n_213),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_L g286 ( 
.A(n_224),
.B(n_116),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_R g287 ( 
.A(n_241),
.B(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_221),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_182),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_241),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_242),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_182),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_262),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_185),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_242),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_265),
.B(n_272),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_253),
.B(n_209),
.C(n_220),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_117),
.B1(n_121),
.B2(n_129),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g301 ( 
.A(n_291),
.Y(n_301)
);

AO22x1_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_206),
.B1(n_169),
.B2(n_187),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_185),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_SL g304 ( 
.A(n_266),
.B(n_132),
.C(n_133),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_207),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_136),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_255),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_259),
.B(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_287),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_167),
.B(n_218),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_188),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

OA22x2_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_184),
.B1(n_175),
.B2(n_167),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_281),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_207),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_141),
.C(n_143),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_264),
.B(n_146),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_206),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_278),
.A2(n_152),
.B1(n_153),
.B2(n_195),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_235),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_258),
.A2(n_205),
.B(n_204),
.C(n_255),
.Y(n_325)
);

NOR2x1p5_ASAP7_75t_SL g326 ( 
.A(n_273),
.B(n_239),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_205),
.B(n_229),
.C(n_194),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_268),
.B(n_206),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_217),
.Y(n_329)
);

CKINVDCx10_ASAP7_75t_R g330 ( 
.A(n_282),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_265),
.A2(n_173),
.B1(n_191),
.B2(n_194),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_289),
.A2(n_229),
.B(n_194),
.C(n_191),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_191),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_260),
.A2(n_249),
.B(n_247),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_199),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_199),
.Y(n_338)
);

AO31x2_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_248),
.A3(n_210),
.B(n_214),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_199),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_210),
.B1(n_214),
.B2(n_217),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_320),
.A2(n_210),
.B(n_214),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_214),
.Y(n_343)
);

AO31x2_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_217),
.A3(n_331),
.B(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_309),
.Y(n_348)
);

AO21x2_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_304),
.B(n_324),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_333),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_332),
.B(n_313),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_300),
.B(n_307),
.Y(n_354)
);

AOI221x1_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_329),
.B1(n_325),
.B2(n_322),
.C(n_327),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_R g356 ( 
.A(n_305),
.B(n_318),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_312),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_293),
.A2(n_294),
.B1(n_328),
.B2(n_316),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_311),
.B(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_326),
.A2(n_308),
.B(n_293),
.C(n_294),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_293),
.A2(n_330),
.B(n_302),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_296),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_298),
.A2(n_310),
.B(n_274),
.C(n_265),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_296),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_296),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_271),
.B1(n_289),
.B2(n_274),
.Y(n_369)
);

OR2x6_ASAP7_75t_L g370 ( 
.A(n_315),
.B(n_291),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_296),
.B(n_306),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_298),
.A2(n_272),
.B1(n_265),
.B2(n_261),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_296),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_297),
.A2(n_274),
.B(n_266),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_367),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

AO31x2_ASAP7_75t_L g382 ( 
.A1(n_366),
.A2(n_375),
.A3(n_357),
.B(n_355),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_376),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g384 ( 
.A1(n_360),
.A2(n_337),
.B(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_370),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_343),
.B(n_342),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_369),
.A2(n_340),
.B(n_358),
.C(n_354),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_341),
.B(n_363),
.Y(n_393)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_370),
.Y(n_395)
);

AO21x2_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_339),
.B(n_344),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_339),
.A2(n_344),
.B(n_352),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_339),
.A2(n_359),
.B(n_374),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_356),
.B(n_347),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_365),
.B(n_372),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_365),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_364),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_374),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_383),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_383),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_401),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_399),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_392),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_399),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_382),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_388),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_398),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_396),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_382),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_412),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_419),
.B(n_382),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_406),
.A2(n_402),
.B1(n_395),
.B2(n_391),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_396),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_389),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_407),
.B(n_400),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_389),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_417),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_431),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_415),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_407),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_427),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

AOI211xp5_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_428),
.B(n_433),
.C(n_434),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_427),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_421),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_443),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_436),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_440),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_445),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_449),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_453),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_447),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_451),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_456),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_459),
.A2(n_456),
.B(n_448),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_456),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_425),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_SL g464 ( 
.A(n_462),
.B(n_444),
.C(n_455),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_463),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_458),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_467),
.A2(n_466),
.B1(n_465),
.B2(n_432),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_457),
.B1(n_455),
.B2(n_450),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_468),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_469),
.B(n_410),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_413),
.B(n_393),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_413),
.B(n_384),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_394),
.B1(n_404),
.B2(n_409),
.Y(n_474)
);


endmodule