module real_jpeg_6046_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_525;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_0),
.A2(n_74),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_0),
.A2(n_74),
.B1(n_204),
.B2(n_394),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_0),
.A2(n_74),
.B1(n_361),
.B2(n_407),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_1),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_1),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_2),
.A2(n_170),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_205),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_2),
.A2(n_205),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_2),
.A2(n_205),
.B1(n_434),
.B2(n_436),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_3),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_3),
.Y(n_435)
);

INVx6_ASAP7_75t_L g437 ( 
.A(n_3),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_49),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_4),
.A2(n_77),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_4),
.A2(n_77),
.B1(n_165),
.B2(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_4),
.A2(n_77),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_5),
.A2(n_130),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_5),
.A2(n_172),
.B1(n_191),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_172),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_5),
.A2(n_71),
.B1(n_172),
.B2(n_357),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_61),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_6),
.A2(n_61),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_6),
.A2(n_61),
.B1(n_129),
.B2(n_417),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_8),
.Y(n_540)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_12),
.Y(n_543)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_14),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_132),
.C(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_14),
.B(n_96),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_14),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_14),
.B(n_143),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_14),
.B(n_106),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_15),
.A2(n_182),
.B1(n_183),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_15),
.A2(n_129),
.B1(n_187),
.B2(n_249),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_15),
.A2(n_187),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_15),
.A2(n_187),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_16),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_16),
.A2(n_30),
.B1(n_51),
.B2(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_16),
.A2(n_51),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_16),
.A2(n_51),
.B1(n_220),
.B2(n_387),
.Y(n_386)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_18),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_18),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_18),
.A2(n_204),
.B1(n_270),
.B2(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_18),
.A2(n_270),
.B1(n_403),
.B2(n_405),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_18),
.A2(n_270),
.B1(n_325),
.B2(n_434),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_538),
.B(n_541),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_64),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_52),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_24),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_24),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_25),
.B(n_167),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_25),
.A2(n_53),
.B1(n_410),
.B2(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_26),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_28),
.Y(n_261)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_28),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_29),
.Y(n_333)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_29),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_29),
.Y(n_407)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_30),
.A2(n_322),
.A3(n_326),
.B1(n_328),
.B2(n_334),
.Y(n_321)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_34),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_35),
.A2(n_353),
.B(n_354),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_35),
.B(n_356),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_53),
.B1(n_54),
.B2(n_62),
.Y(n_52)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_48),
.Y(n_357)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_52),
.B(n_66),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_62),
.B1(n_70),
.B2(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_75),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_53),
.A2(n_355),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_53),
.A2(n_62),
.B1(n_70),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_60),
.B(n_167),
.Y(n_334)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_60),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_62),
.A2(n_433),
.B(n_464),
.Y(n_474)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_152),
.B(n_537),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_148),
.C(n_149),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_67),
.A2(n_68),
.B1(n_533),
.B2(n_534),
.Y(n_532)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_78),
.C(n_114),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_69),
.B(n_525),
.Y(n_524)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_72),
.A2(n_167),
.B(n_334),
.Y(n_353)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_73),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_78),
.A2(n_114),
.B1(n_115),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_78),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_79),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_79),
.A2(n_109),
.B1(n_296),
.B2(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_79),
.A2(n_109),
.B1(n_402),
.B2(n_408),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_79),
.A2(n_105),
.B1(n_109),
.B2(n_514),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_96),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_83),
.Y(n_279)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx6_ASAP7_75t_L g366 ( 
.A(n_88),
.Y(n_366)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_94),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_95),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_95),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_96),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_96),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

AOI22x1_ASAP7_75t_L g438 ( 
.A1(n_96),
.A2(n_150),
.B1(n_303),
.B2(n_439),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_96),
.A2(n_150),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_100),
.Y(n_282)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_100),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_102),
.Y(n_399)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_109),
.B(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_109),
.A2(n_296),
.B(n_302),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_114),
.A2(n_115),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_114),
.B(n_509),
.C(n_512),
.Y(n_520)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_142),
.B(n_144),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_162),
.B(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_116),
.A2(n_142),
.B1(n_202),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_116),
.A2(n_168),
.B(n_248),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_116),
.A2(n_142),
.B1(n_368),
.B2(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_117),
.B(n_169),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_117),
.A2(n_143),
.B1(n_393),
.B2(n_397),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_117),
.A2(n_143),
.B1(n_397),
.B2(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_117),
.A2(n_143),
.B1(n_416),
.B2(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_131),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_125),
.B2(n_129),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_121),
.Y(n_251)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_131),
.A2(n_202),
.B(n_206),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_136),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_138),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_138),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_139),
.Y(n_391)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_142),
.A2(n_206),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_144),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_147),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_148),
.B(n_149),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_150),
.A2(n_254),
.B(n_258),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_150),
.B(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_150),
.A2(n_258),
.B(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_531),
.B(n_536),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_503),
.B(n_528),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_372),
.A3(n_479),
.B1(n_497),
.C1(n_498),
.Y(n_154)
);

AOI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_315),
.B(n_371),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_287),
.B(n_314),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_242),
.B(n_286),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_209),
.B(n_241),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_179),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_160),
.B(n_179),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_173),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_161),
.A2(n_173),
.B1(n_174),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_188),
.B(n_194),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_167),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_170),
.Y(n_277)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_178),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_178),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_199),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_200),
.C(n_208),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_188),
.B(n_194),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_188),
.A2(n_337),
.B1(n_338),
.B2(n_341),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_188),
.A2(n_378),
.B1(n_383),
.B2(n_386),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_188),
.A2(n_386),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_189),
.A2(n_268),
.B1(n_307),
.B2(n_312),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_189),
.A2(n_342),
.B1(n_422),
.B2(n_430),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_193),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_208),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_231),
.B(n_240),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_217),
.B(n_230),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_215),
.Y(n_340)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_215),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_229),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_229),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_225),
.B(n_228),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_267),
.B(n_274),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_238),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_244),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_265),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_252),
.C(n_265),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_251),
.Y(n_419)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_276),
.A3(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_275),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_288),
.B(n_289),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_313),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_293),
.C(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_304),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_305),
.C(n_306),
.Y(n_347)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_307),
.Y(n_337)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_316),
.B(n_317),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_350),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_318)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_335),
.B2(n_336),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_321),
.B(n_335),
.Y(n_475)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx6_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_347),
.B(n_348),
.C(n_350),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_358),
.B2(n_370),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_351),
.B(n_359),
.C(n_367),
.Y(n_488)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_358),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_367),
.Y(n_358)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_465),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_373),
.A2(n_465),
.B(n_499),
.C(n_502),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_440),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_374),
.B(n_440),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_413),
.C(n_425),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_375),
.B(n_413),
.CI(n_425),
.CON(n_478),
.SN(n_478)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_400),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_401),
.C(n_409),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_392),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_377),
.B(n_392),
.Y(n_471)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_409),
.Y(n_400)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_402),
.Y(n_439)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_420),
.B2(n_424),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_420),
.Y(n_458)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_424),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_420),
.A2(n_458),
.B(n_461),
.Y(n_506)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.C(n_438),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_427),
.B(n_429),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_431),
.A2(n_432),
.B1(n_438),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_438),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_441),
.B(n_444),
.C(n_456),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_456),
.B2(n_457),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_452),
.B(n_455),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_453),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

FAx1_ASAP7_75t_SL g505 ( 
.A(n_455),
.B(n_506),
.CI(n_507),
.CON(n_505),
.SN(n_505)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_506),
.C(n_507),
.Y(n_527)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_478),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_478),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.C(n_472),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_467),
.A2(n_468),
.B1(n_471),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_471),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.C(n_476),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_473),
.A2(n_474),
.B1(n_476),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_476),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_478),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_492),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_481),
.A2(n_500),
.B(n_501),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_489),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_489),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.C(n_488),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_495),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_488),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_494),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_517),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_516),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_516),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_505),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_509),
.B1(n_511),
.B2(n_515),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_508),
.A2(n_509),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_519),
.C(n_523),
.Y(n_535)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_511),
.Y(n_515)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_517),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_527),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_527),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_532),
.B(n_535),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

BUFx4f_ASAP7_75t_SL g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_539),
.Y(n_542)
);

INVx13_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);


endmodule