module real_aes_2345_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g237 ( .A(n_0), .B(n_158), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_1), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_2), .B(n_142), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_3), .B(n_160), .Y(n_510) );
INVx1_ASAP7_75t_L g149 ( .A(n_4), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_5), .B(n_142), .Y(n_141) );
NAND2xp33_ASAP7_75t_SL g228 ( .A(n_6), .B(n_148), .Y(n_228) );
INVx1_ASAP7_75t_L g209 ( .A(n_7), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_8), .Y(n_120) );
AND2x2_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
XNOR2xp5_ASAP7_75t_L g127 ( .A(n_10), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g520 ( .A(n_10), .B(n_225), .Y(n_520) );
AND2x2_ASAP7_75t_L g512 ( .A(n_11), .B(n_199), .Y(n_512) );
INVx2_ASAP7_75t_L g138 ( .A(n_12), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_13), .B(n_160), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_14), .B(n_482), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
AOI221x1_ASAP7_75t_L g222 ( .A1(n_16), .A2(n_151), .B1(n_223), .B2(n_225), .C(n_227), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_17), .B(n_142), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_18), .B(n_142), .Y(n_543) );
INVx1_ASAP7_75t_L g116 ( .A(n_19), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_20), .A2(n_91), .B1(n_142), .B2(n_210), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_21), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_22), .A2(n_151), .B(n_156), .Y(n_150) );
AOI221xp5_ASAP7_75t_SL g186 ( .A1(n_23), .A2(n_36), .B1(n_142), .B2(n_151), .C(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_24), .B(n_158), .Y(n_157) );
OR2x2_ASAP7_75t_L g139 ( .A(n_25), .B(n_90), .Y(n_139) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_25), .A2(n_90), .B(n_138), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_26), .B(n_160), .Y(n_198) );
INVxp67_ASAP7_75t_L g221 ( .A(n_27), .Y(n_221) );
AND2x2_ASAP7_75t_L g182 ( .A(n_28), .B(n_172), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_29), .A2(n_151), .B(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_30), .A2(n_225), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_31), .B(n_160), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_32), .A2(n_151), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_33), .B(n_160), .Y(n_538) );
AND2x2_ASAP7_75t_L g148 ( .A(n_34), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g152 ( .A(n_34), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g217 ( .A(n_34), .Y(n_217) );
OR2x6_ASAP7_75t_L g114 ( .A(n_35), .B(n_115), .Y(n_114) );
XOR2xp5_ASAP7_75t_L g480 ( .A(n_37), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_38), .B(n_142), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_39), .A2(n_83), .B1(n_151), .B2(n_215), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_40), .B(n_160), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_41), .A2(n_75), .B1(n_467), .B2(n_468), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_41), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_42), .B(n_142), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_43), .B(n_158), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_44), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_45), .A2(n_151), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_46), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g240 ( .A(n_47), .B(n_172), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_48), .B(n_158), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_49), .B(n_172), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_50), .B(n_142), .Y(n_526) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_51), .A2(n_465), .B1(n_466), .B2(n_469), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_51), .Y(n_469) );
INVx1_ASAP7_75t_L g145 ( .A(n_52), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_52), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_53), .B(n_160), .Y(n_518) );
AND2x2_ASAP7_75t_L g554 ( .A(n_54), .B(n_172), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_55), .B(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_56), .B(n_158), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_57), .B(n_158), .Y(n_537) );
AND2x2_ASAP7_75t_L g173 ( .A(n_58), .B(n_172), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_59), .B(n_142), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_60), .B(n_160), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_61), .B(n_142), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_62), .A2(n_151), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_63), .B(n_158), .Y(n_169) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_64), .B(n_137), .Y(n_201) );
AND2x2_ASAP7_75t_L g549 ( .A(n_65), .B(n_137), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_66), .A2(n_151), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_67), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_68), .B(n_199), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_69), .B(n_158), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_70), .B(n_158), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_71), .A2(n_94), .B1(n_151), .B2(n_215), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_72), .B(n_160), .Y(n_546) );
INVx1_ASAP7_75t_L g147 ( .A(n_73), .Y(n_147) );
INVx1_ASAP7_75t_L g153 ( .A(n_73), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_74), .B(n_158), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_75), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_76), .A2(n_151), .B(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_77), .A2(n_151), .B(n_500), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_78), .A2(n_151), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g540 ( .A(n_79), .B(n_137), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_80), .B(n_172), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_81), .B(n_142), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_82), .A2(n_85), .B1(n_142), .B2(n_210), .Y(n_251) );
INVx1_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_86), .B(n_158), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_87), .B(n_158), .Y(n_189) );
AND2x2_ASAP7_75t_L g503 ( .A(n_88), .B(n_199), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_89), .A2(n_151), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_92), .B(n_160), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_93), .A2(n_151), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_95), .B(n_160), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_96), .A2(n_103), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_96), .Y(n_483) );
INVxp67_ASAP7_75t_L g224 ( .A(n_97), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_98), .B(n_142), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_99), .B(n_160), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_100), .A2(n_151), .B(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g548 ( .A(n_101), .Y(n_548) );
BUFx2_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_102), .B(n_474), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_103), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_121), .B(n_799), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_107), .B(n_800), .Y(n_799) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_109), .B(n_118), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g473 ( .A(n_111), .Y(n_473) );
BUFx3_ASAP7_75t_L g477 ( .A(n_111), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x6_ASAP7_75t_SL g489 ( .A(n_112), .B(n_114), .Y(n_489) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_112), .B(n_113), .Y(n_791) );
OR2x2_ASAP7_75t_L g798 ( .A(n_112), .B(n_114), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OA22x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_126), .B1(n_478), .B2(n_479), .Y(n_121) );
CKINVDCx11_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_470), .B(n_474), .Y(n_126) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B1(n_463), .B2(n_464), .Y(n_128) );
OAI22x1_ASAP7_75t_L g793 ( .A1(n_129), .A2(n_486), .B1(n_791), .B2(n_794), .Y(n_793) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_130), .A2(n_486), .B1(n_490), .B2(n_789), .Y(n_485) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_374), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_296), .C(n_346), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_263), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_183), .B1(n_202), .B2(n_245), .C(n_255), .Y(n_133) );
INVx1_ASAP7_75t_SL g345 ( .A(n_134), .Y(n_345) );
AND2x4_ASAP7_75t_SL g134 ( .A(n_135), .B(n_163), .Y(n_134) );
INVx2_ASAP7_75t_L g267 ( .A(n_135), .Y(n_267) );
OR2x2_ASAP7_75t_L g289 ( .A(n_135), .B(n_280), .Y(n_289) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_135), .Y(n_304) );
INVx5_ASAP7_75t_L g311 ( .A(n_135), .Y(n_311) );
AND2x4_ASAP7_75t_L g317 ( .A(n_135), .B(n_175), .Y(n_317) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_135), .B(n_247), .Y(n_320) );
OR2x2_ASAP7_75t_L g329 ( .A(n_135), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g336 ( .A(n_135), .B(n_164), .Y(n_336) );
AND2x2_ASAP7_75t_L g437 ( .A(n_135), .B(n_174), .Y(n_437) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g162 ( .A(n_138), .B(n_139), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_162), .Y(n_140) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
INVx1_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
AND2x6_ASAP7_75t_L g158 ( .A(n_144), .B(n_153), .Y(n_158) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g160 ( .A(n_146), .B(n_155), .Y(n_160) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
AND2x2_ASAP7_75t_L g154 ( .A(n_149), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
BUFx3_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
INVx2_ASAP7_75t_L g219 ( .A(n_153), .Y(n_219) );
AND2x4_ASAP7_75t_L g215 ( .A(n_154), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_158), .B(n_548), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_161), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_161), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_161), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_161), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_161), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_161), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_161), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_161), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_161), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_161), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_161), .A2(n_559), .B(n_560), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_162), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_162), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_162), .B(n_224), .Y(n_223) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_162), .B(n_228), .C(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_162), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_162), .A2(n_556), .B(n_557), .Y(n_555) );
INVx3_ASAP7_75t_SL g288 ( .A(n_163), .Y(n_288) );
AND2x2_ASAP7_75t_L g332 ( .A(n_163), .B(n_247), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_163), .A2(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g373 ( .A(n_163), .B(n_311), .Y(n_373) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_174), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_164), .B(n_175), .Y(n_254) );
OR2x2_ASAP7_75t_L g258 ( .A(n_164), .B(n_175), .Y(n_258) );
INVx1_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_164), .Y(n_278) );
INVx2_ASAP7_75t_L g286 ( .A(n_164), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_164), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g395 ( .A(n_164), .B(n_280), .Y(n_395) );
AND2x2_ASAP7_75t_L g410 ( .A(n_164), .B(n_247), .Y(n_410) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_171), .B(n_173), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_171), .A2(n_176), .B(n_182), .Y(n_175) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_171), .A2(n_176), .B(n_182), .Y(n_330) );
AOI21x1_ASAP7_75t_L g505 ( .A1(n_171), .A2(n_506), .B(n_512), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_172), .A2(n_186), .B(n_190), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_172), .A2(n_498), .B(n_499), .Y(n_497) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_172), .A2(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g279 ( .A(n_175), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_175), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_183), .B(n_403), .Y(n_402) );
NOR2x1p5_ASAP7_75t_L g183 ( .A(n_184), .B(n_191), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g231 ( .A(n_185), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_185), .B(n_192), .Y(n_261) );
INVx1_ASAP7_75t_L g271 ( .A(n_185), .Y(n_271) );
INVx2_ASAP7_75t_L g294 ( .A(n_185), .Y(n_294) );
INVx2_ASAP7_75t_L g300 ( .A(n_185), .Y(n_300) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_185), .Y(n_370) );
OR2x2_ASAP7_75t_L g401 ( .A(n_185), .B(n_192), .Y(n_401) );
OR2x2_ASAP7_75t_L g417 ( .A(n_191), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_SL g205 ( .A(n_192), .B(n_206), .Y(n_205) );
AND2x4_ASAP7_75t_L g243 ( .A(n_192), .B(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g281 ( .A(n_192), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g293 ( .A(n_192), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_192), .B(n_272), .Y(n_306) );
OR2x2_ASAP7_75t_L g314 ( .A(n_192), .B(n_206), .Y(n_314) );
INVx2_ASAP7_75t_L g341 ( .A(n_192), .Y(n_341) );
INVx1_ASAP7_75t_L g359 ( .A(n_192), .Y(n_359) );
NOR2xp33_ASAP7_75t_R g392 ( .A(n_192), .B(n_232), .Y(n_392) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_199), .Y(n_193) );
INVx2_ASAP7_75t_SL g249 ( .A(n_199), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_199), .A2(n_543), .B(n_544), .Y(n_542) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g226 ( .A(n_200), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_203), .B(n_241), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_203), .A2(n_284), .B1(n_287), .B2(n_290), .Y(n_283) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_230), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g298 ( .A(n_205), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g333 ( .A(n_205), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g412 ( .A(n_205), .B(n_390), .Y(n_412) );
INVx3_ASAP7_75t_L g244 ( .A(n_206), .Y(n_244) );
AND2x4_ASAP7_75t_L g272 ( .A(n_206), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_206), .B(n_232), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_206), .B(n_294), .Y(n_339) );
AND2x2_ASAP7_75t_L g344 ( .A(n_206), .B(n_341), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_206), .B(n_231), .Y(n_381) );
INVx1_ASAP7_75t_L g451 ( .A(n_206), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_206), .B(n_369), .Y(n_462) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_222), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B1(n_215), .B2(n_220), .Y(n_207) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
NOR2x1p5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g533 ( .A(n_225), .Y(n_533) );
INVx4_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_226), .A2(n_234), .B(n_240), .Y(n_233) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_226), .A2(n_514), .B(n_520), .Y(n_513) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g242 ( .A(n_232), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_232), .B(n_244), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_232), .Y(n_273) );
AND2x2_ASAP7_75t_L g299 ( .A(n_232), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g315 ( .A(n_232), .B(n_294), .Y(n_315) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_232), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_232), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g404 ( .A(n_232), .Y(n_404) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_239), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_242), .B(n_271), .Y(n_282) );
AOI221x1_ASAP7_75t_SL g376 ( .A1(n_243), .A2(n_377), .B1(n_380), .B2(n_382), .C(n_386), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_243), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g434 ( .A(n_243), .B(n_299), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_243), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g365 ( .A(n_244), .B(n_293), .Y(n_365) );
AND2x2_ASAP7_75t_L g403 ( .A(n_244), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
AND2x2_ASAP7_75t_L g256 ( .A(n_247), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g351 ( .A(n_247), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_247), .B(n_267), .Y(n_356) );
AND2x4_ASAP7_75t_L g385 ( .A(n_247), .B(n_286), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_247), .B(n_317), .Y(n_421) );
OR2x2_ASAP7_75t_L g439 ( .A(n_247), .B(n_370), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_247), .B(n_330), .Y(n_449) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
AOI21x1_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_253), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g305 ( .A(n_254), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_254), .A2(n_313), .B1(n_316), .B2(n_318), .Y(n_312) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_259), .Y(n_255) );
INVx2_ASAP7_75t_L g268 ( .A(n_256), .Y(n_268) );
AND2x2_ASAP7_75t_L g407 ( .A(n_257), .B(n_267), .Y(n_407) );
AND2x2_ASAP7_75t_L g453 ( .A(n_257), .B(n_320), .Y(n_453) );
AND2x2_ASAP7_75t_L g458 ( .A(n_257), .B(n_309), .Y(n_458) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AOI32xp33_ASAP7_75t_L g427 ( .A1(n_259), .A2(n_329), .A3(n_409), .B1(n_428), .B2(n_430), .Y(n_427) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
AOI211xp5_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_269), .B(n_274), .C(n_283), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_266), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_267), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g447 ( .A(n_267), .Y(n_447) );
AND2x2_ASAP7_75t_L g357 ( .A(n_269), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_270), .B(n_272), .Y(n_269) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_270), .Y(n_457) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_271), .Y(n_326) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_271), .Y(n_426) );
INVx1_ASAP7_75t_L g323 ( .A(n_272), .Y(n_323) );
AND2x2_ASAP7_75t_L g389 ( .A(n_272), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_272), .B(n_400), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_281), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_276), .A2(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g285 ( .A(n_280), .B(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_285), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g416 ( .A(n_285), .Y(n_416) );
AND2x2_ASAP7_75t_L g446 ( .A(n_285), .B(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_286), .Y(n_423) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_288), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g363 ( .A(n_289), .Y(n_363) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g322 ( .A(n_293), .B(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_294), .Y(n_390) );
AND2x2_ASAP7_75t_L g399 ( .A(n_295), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_319), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_306), .B2(n_307), .C(n_312), .Y(n_297) );
INVx1_ASAP7_75t_L g418 ( .A(n_299), .Y(n_418) );
INVxp33_ASAP7_75t_SL g450 ( .A(n_299), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_301), .A2(n_397), .B(n_405), .Y(n_396) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_305), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
AND2x2_ASAP7_75t_L g353 ( .A(n_306), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g372 ( .A(n_306), .B(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g433 ( .A1(n_306), .A2(n_434), .B1(n_435), .B2(n_438), .Y(n_433) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OR2x2_ASAP7_75t_L g328 ( .A(n_309), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_309), .B(n_317), .Y(n_367) );
AND2x4_ASAP7_75t_L g384 ( .A(n_311), .B(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_311), .B(n_385), .Y(n_431) );
AND2x2_ASAP7_75t_L g443 ( .A(n_311), .B(n_395), .Y(n_443) );
NAND2xp33_ASAP7_75t_L g428 ( .A(n_313), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_SL g371 ( .A(n_314), .Y(n_371) );
INVx1_ASAP7_75t_L g442 ( .A(n_315), .Y(n_442) );
INVx2_ASAP7_75t_SL g394 ( .A(n_317), .Y(n_394) );
AOI211xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_321), .B(n_324), .C(n_342), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B(n_331), .C(n_335), .Y(n_324) );
OR2x6_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g354 ( .A(n_326), .Y(n_354) );
INVx1_ASAP7_75t_SL g379 ( .A(n_329), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_329), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_334), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_338), .A2(n_421), .B1(n_422), .B2(n_424), .Y(n_420) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
OAI211xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_352), .B(n_355), .C(n_360), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B1(n_366), .B2(n_368), .C(n_372), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g452 ( .A1(n_371), .A2(n_453), .B1(n_454), .B2(n_458), .C1(n_459), .C2(n_461), .Y(n_452) );
INVx2_ASAP7_75t_L g387 ( .A(n_373), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_413), .C(n_432), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_396), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_384), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_385), .B(n_447), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_393), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVxp33_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_394), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_402), .A2(n_406), .B1(n_408), .B2(n_411), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_417), .B(n_419), .C(n_427), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_440), .C(n_452), .Y(n_432) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_451), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_448), .B(n_450), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVxp33_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
CKINVDCx11_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
AO221x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_485), .B1(n_792), .B2(n_793), .C(n_795), .Y(n_479) );
INVx1_ASAP7_75t_L g792 ( .A(n_480), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g794 ( .A(n_490), .Y(n_794) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_693), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_618), .C(n_654), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_592), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_521), .B(n_550), .C(n_575), .Y(n_493) );
AND2x2_ASAP7_75t_L g683 ( .A(n_494), .B(n_552), .Y(n_683) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_495), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g716 ( .A(n_495), .B(n_598), .Y(n_716) );
AND2x2_ASAP7_75t_L g732 ( .A(n_495), .B(n_567), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_495), .B(n_742), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g765 ( .A(n_495), .B(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_SL g562 ( .A(n_496), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_577), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_496), .B(n_504), .Y(n_653) );
BUFx2_ASAP7_75t_L g658 ( .A(n_496), .Y(n_658) );
AND2x2_ASAP7_75t_L g702 ( .A(n_496), .B(n_513), .Y(n_702) );
AND2x4_ASAP7_75t_L g774 ( .A(n_496), .B(n_775), .Y(n_774) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_496), .B(n_566), .Y(n_786) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_504), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g705 ( .A(n_504), .Y(n_705) );
BUFx2_ASAP7_75t_L g754 ( .A(n_504), .Y(n_754) );
INVx1_ASAP7_75t_L g776 ( .A(n_504), .Y(n_776) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx3_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_505), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
INVx2_ASAP7_75t_L g566 ( .A(n_513), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_513), .B(n_563), .Y(n_567) );
INVx2_ASAP7_75t_L g642 ( .A(n_513), .Y(n_642) );
OR2x2_ASAP7_75t_L g649 ( .A(n_513), .B(n_598), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AND2x2_ASAP7_75t_L g604 ( .A(n_521), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_601), .Y(n_638) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
AND2x2_ASAP7_75t_L g674 ( .A(n_522), .B(n_573), .Y(n_674) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g631 ( .A(n_523), .B(n_532), .Y(n_631) );
AND2x2_ASAP7_75t_L g750 ( .A(n_523), .B(n_541), .Y(n_750) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g572 ( .A(n_524), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g646 ( .A(n_524), .B(n_532), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_524), .B(n_553), .Y(n_651) );
OR2x2_ASAP7_75t_L g714 ( .A(n_524), .B(n_541), .Y(n_714) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
AND2x2_ASAP7_75t_L g552 ( .A(n_531), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g591 ( .A(n_531), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g531 ( .A(n_532), .B(n_541), .Y(n_531) );
AO21x1_ASAP7_75t_SL g532 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_532) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_533), .A2(n_534), .B(n_540), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
AND2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g617 ( .A(n_541), .Y(n_617) );
NAND2x1_ASAP7_75t_L g627 ( .A(n_541), .B(n_553), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_570), .Y(n_632) );
BUFx2_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
AND2x2_ASAP7_75t_L g724 ( .A(n_541), .B(n_603), .Y(n_724) );
AND2x2_ASAP7_75t_L g735 ( .A(n_541), .B(n_573), .Y(n_735) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_561), .B1(n_567), .B2(n_568), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_552), .A2(n_732), .B1(n_782), .B2(n_787), .Y(n_781) );
INVx4_ASAP7_75t_L g570 ( .A(n_553), .Y(n_570) );
INVx2_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_553), .Y(n_672) );
OR2x2_ASAP7_75t_L g687 ( .A(n_553), .B(n_573), .Y(n_687) );
OR2x2_ASAP7_75t_SL g713 ( .A(n_553), .B(n_714), .Y(n_713) );
OR2x6_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_SL g594 ( .A(n_562), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_562), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g662 ( .A(n_562), .B(n_610), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_562), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g584 ( .A(n_563), .Y(n_584) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
AND2x2_ASAP7_75t_L g665 ( .A(n_563), .B(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g775 ( .A(n_563), .Y(n_775) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_565), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_565), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g583 ( .A(n_566), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_567), .B(n_716), .Y(n_715) );
AOI321xp33_ASAP7_75t_L g737 ( .A1(n_568), .A2(n_639), .A3(n_707), .B1(n_738), .B2(n_739), .C(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_569), .Y(n_636) );
AND2x2_ASAP7_75t_L g661 ( .A(n_569), .B(n_590), .Y(n_661) );
AND2x2_ASAP7_75t_L g736 ( .A(n_569), .B(n_646), .Y(n_736) );
INVx1_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
BUFx2_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_570), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g660 ( .A(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
BUFx2_ASAP7_75t_L g667 ( .A(n_572), .Y(n_667) );
INVx2_ASAP7_75t_L g603 ( .A(n_573), .Y(n_603) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_573), .Y(n_626) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI21xp33_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_585), .B(n_588), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_576), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx3_ASAP7_75t_L g610 ( .A(n_578), .Y(n_610) );
AND2x2_ASAP7_75t_L g641 ( .A(n_578), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g598 ( .A(n_579), .B(n_580), .Y(n_598) );
INVx1_ASAP7_75t_L g681 ( .A(n_583), .Y(n_681) );
INVx1_ASAP7_75t_SL g766 ( .A(n_584), .Y(n_766) );
INVxp33_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_587), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g692 ( .A(n_587), .B(n_649), .Y(n_692) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g696 ( .A(n_589), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_589), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_627), .Y(n_682) );
NOR4xp25_ASAP7_75t_L g777 ( .A(n_590), .B(n_621), .C(n_778), .D(n_779), .Y(n_777) );
OR2x2_ASAP7_75t_L g745 ( .A(n_591), .B(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_599), .B1(n_604), .B2(n_606), .C(n_611), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g620 ( .A(n_595), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g677 ( .A(n_597), .Y(n_677) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g700 ( .A(n_598), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_598), .B(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g644 ( .A(n_601), .B(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_603), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx2_ASAP7_75t_L g621 ( .A(n_608), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_608), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g613 ( .A(n_610), .Y(n_613) );
OAI321xp33_ASAP7_75t_L g725 ( .A1(n_610), .A2(n_718), .A3(n_726), .B1(n_731), .B2(n_733), .C(n_737), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g680 ( .A(n_613), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g780 ( .A(n_616), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g760 ( .A(n_617), .B(n_631), .Y(n_760) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_633), .C(n_637), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g729 ( .A(n_626), .Y(n_729) );
INVx3_ASAP7_75t_L g668 ( .A(n_627), .Y(n_668) );
OR2x2_ASAP7_75t_L g771 ( .A(n_627), .B(n_645), .Y(n_771) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_629), .A2(n_713), .B1(n_715), .B2(n_717), .Y(n_712) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g711 ( .A(n_632), .Y(n_711) );
OR2x2_ASAP7_75t_L g788 ( .A(n_632), .B(n_645), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_641), .B(n_658), .Y(n_757) );
AND2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g708 ( .A(n_642), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B1(n_650), .B2(n_652), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_645), .A2(n_688), .B(n_690), .C(n_692), .Y(n_689) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_648), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_648), .B(n_740), .Y(n_762) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g734 ( .A(n_651), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_685), .B(n_688), .C(n_689), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_655), .B(n_669), .C(n_684), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_661), .B2(n_662), .C1(n_663), .C2(n_666), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g718 ( .A(n_658), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_691), .Y(n_744) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g678 ( .A(n_665), .Y(n_678) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g783 ( .A(n_667), .B(n_700), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_668), .A2(n_759), .B1(n_761), .B2(n_763), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI21xp5_ASAP7_75t_SL g743 ( .A1(n_676), .A2(n_744), .B(n_745), .Y(n_743) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g691 ( .A(n_677), .Y(n_691) );
AND2x2_ASAP7_75t_L g785 ( .A(n_677), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g769 ( .A(n_681), .Y(n_769) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g698 ( .A(n_687), .B(n_688), .Y(n_698) );
INVx1_ASAP7_75t_L g751 ( .A(n_687), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_725), .C(n_747), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_701), .C(n_706), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_696), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_712), .C(n_719), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g730 ( .A(n_713), .Y(n_730) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_714), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_716), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g778 ( .A(n_716), .Y(n_778) );
AND2x2_ASAP7_75t_L g768 ( .A(n_718), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g746 ( .A(n_722), .Y(n_746) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_734), .A2(n_768), .B1(n_770), .B2(n_772), .C(n_777), .Y(n_767) );
OAI21xp33_ASAP7_75t_SL g782 ( .A1(n_739), .A2(n_783), .B(n_784), .Y(n_782) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_758), .C(n_767), .D(n_781), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B1(n_755), .B2(n_756), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
BUFx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
endmodule