module fake_jpeg_30862_n_473 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_54),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_18),
.B(n_8),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_57),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_46),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_63),
.B(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_0),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_22),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_76),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_6),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_29),
.B(n_6),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_81),
.B(n_36),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_29),
.B(n_6),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_6),
.Y(n_90)
);

BUFx6f_ASAP7_75t_SL g91 ( 
.A(n_44),
.Y(n_91)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_95),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_96),
.B(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_48),
.A2(n_16),
.B1(n_32),
.B2(n_41),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_118),
.A2(n_125),
.B1(n_131),
.B2(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_16),
.B1(n_43),
.B2(n_36),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_81),
.B1(n_76),
.B2(n_24),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_52),
.A2(n_32),
.B1(n_41),
.B2(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_140),
.Y(n_194)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_57),
.B1(n_93),
.B2(n_56),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_43),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_51),
.Y(n_153)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_49),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_50),
.A2(n_32),
.B1(n_44),
.B2(n_24),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_32),
.B1(n_44),
.B2(n_24),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_72),
.B1(n_44),
.B2(n_91),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_162),
.Y(n_197)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_156),
.A2(n_171),
.B1(n_118),
.B2(n_26),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_65),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_65),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_186),
.Y(n_206)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_150),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_173),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_98),
.A2(n_92),
.B1(n_86),
.B2(n_70),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_189),
.B1(n_147),
.B2(n_105),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_181),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_109),
.A2(n_53),
.B1(n_67),
.B2(n_71),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_104),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_180),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_107),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_100),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_188),
.B1(n_195),
.B2(n_137),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_89),
.A3(n_44),
.B1(n_55),
.B2(n_41),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_151),
.A3(n_55),
.B1(n_105),
.B2(n_47),
.Y(n_223)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_193),
.Y(n_213)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_127),
.A2(n_68),
.B1(n_87),
.B2(n_78),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_26),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_191),
.Y(n_232)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_110),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_110),
.A2(n_69),
.B1(n_74),
.B2(n_21),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_127),
.B1(n_148),
.B2(n_146),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_SL g200 ( 
.A(n_159),
.B(n_144),
.C(n_131),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_200),
.A2(n_165),
.B(n_154),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_211),
.B1(n_212),
.B2(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_89),
.C(n_141),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_222),
.C(n_224),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_137),
.B1(n_108),
.B2(n_125),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_135),
.B1(n_148),
.B2(n_146),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_66),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_217),
.B1(n_200),
.B2(n_230),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_152),
.B(n_47),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_106),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_106),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_220),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_235),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_249),
.B1(n_252),
.B2(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_156),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_244),
.Y(n_280)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_243),
.A2(n_260),
.B(n_225),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_164),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_186),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_209),
.C(n_199),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_161),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_253),
.Y(n_282)
);

A2O1A1O1Ixp25_ASAP7_75t_L g248 ( 
.A1(n_197),
.A2(n_206),
.B(n_223),
.C(n_222),
.D(n_226),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_21),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_189),
.B1(n_130),
.B2(n_135),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_187),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_228),
.Y(n_268)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_256),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_130),
.B1(n_62),
.B2(n_64),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_176),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_182),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_161),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_157),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_262),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_208),
.A2(n_173),
.B(n_183),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_204),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_160),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_202),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_175),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_221),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_235),
.B1(n_234),
.B2(n_238),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_268),
.B(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_233),
.A2(n_215),
.B1(n_229),
.B2(n_61),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_275),
.B1(n_277),
.B2(n_252),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_243),
.B(n_227),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_233),
.A2(n_229),
.B1(n_196),
.B2(n_163),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_257),
.A2(n_77),
.B1(n_209),
.B2(n_174),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_199),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_284),
.B(n_289),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_287),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_246),
.B(n_157),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_241),
.B(n_236),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_291),
.B(n_234),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_192),
.B1(n_188),
.B2(n_214),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_262),
.B1(n_261),
.B2(n_264),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_169),
.A3(n_193),
.B1(n_218),
.B2(n_219),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_259),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_201),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_297),
.B(n_301),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_308),
.B(n_287),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_315),
.B1(n_317),
.B2(n_269),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_306),
.B(n_310),
.Y(n_351)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_245),
.B(n_242),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_314),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_253),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_319),
.B1(n_320),
.B2(n_97),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_271),
.A2(n_237),
.B1(n_248),
.B2(n_250),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_321),
.B1(n_278),
.B2(n_292),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_254),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_313),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_280),
.B1(n_274),
.B2(n_290),
.Y(n_317)
);

AOI22x1_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_251),
.B1(n_262),
.B2(n_260),
.Y(n_319)
);

AOI22x1_ASAP7_75t_L g320 ( 
.A1(n_265),
.A2(n_251),
.B1(n_247),
.B2(n_214),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_239),
.B1(n_225),
.B2(n_202),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_324),
.Y(n_348)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_303),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_289),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_329),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_281),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_276),
.C(n_285),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_341),
.C(n_342),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_332),
.A2(n_343),
.B1(n_321),
.B2(n_305),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_307),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_334),
.B(n_338),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_336),
.A2(n_355),
.B1(n_319),
.B2(n_320),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_25),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_316),
.B(n_278),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_346),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_273),
.C(n_268),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_280),
.C(n_286),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_277),
.B1(n_286),
.B2(n_293),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_295),
.C(n_219),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_330),
.C(n_329),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_323),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_353),
.Y(n_362)
);

NOR3xp33_ASAP7_75t_SL g346 ( 
.A(n_302),
.B(n_201),
.C(n_151),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_308),
.A2(n_267),
.B(n_170),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_324),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_298),
.A2(n_239),
.B1(n_190),
.B2(n_167),
.Y(n_350)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_352),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_201),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_298),
.A2(n_167),
.B1(n_102),
.B2(n_97),
.Y(n_354)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_350),
.B1(n_333),
.B2(n_354),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_360),
.A2(n_379),
.B1(n_343),
.B2(n_328),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_311),
.B1(n_312),
.B2(n_319),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_336),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_369),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_11),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_201),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_371),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_320),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_376),
.C(n_381),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_352),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_375),
.B(n_377),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_335),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_333),
.A2(n_155),
.B1(n_145),
.B2(n_121),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_339),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_342),
.B(n_121),
.C(n_42),
.Y(n_381)
);

BUFx8_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_383),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_13),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_360),
.A2(n_347),
.B(n_332),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_393),
.B(n_402),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_351),
.C(n_346),
.Y(n_389)
);

OAI221xp5_ASAP7_75t_L g404 ( 
.A1(n_389),
.A2(n_356),
.B1(n_371),
.B2(n_380),
.C(n_381),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_79),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_392),
.A2(n_398),
.B1(n_13),
.B2(n_14),
.Y(n_416)
);

NAND2x1_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_353),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_344),
.C(n_345),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_397),
.C(n_23),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_326),
.C(n_42),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_367),
.A2(n_358),
.B1(n_370),
.B2(n_368),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_73),
.B1(n_42),
.B2(n_0),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_401),
.B(n_370),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_12),
.B(n_14),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_404),
.A2(n_411),
.B1(n_416),
.B2(n_396),
.Y(n_424)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_357),
.C(n_373),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_405),
.B(n_415),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g406 ( 
.A(n_390),
.B(n_362),
.CI(n_373),
.CON(n_406),
.SN(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_408),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_362),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_21),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_410),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_23),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_418),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_13),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_13),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_34),
.C(n_28),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_399),
.C(n_400),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_37),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_419),
.A2(n_384),
.B1(n_395),
.B2(n_402),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_414),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_423),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_427),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_34),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_420),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_416),
.A2(n_385),
.B1(n_389),
.B2(n_387),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_407),
.A2(n_400),
.B(n_393),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_432),
.A2(n_12),
.B(n_11),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_415),
.A2(n_392),
.B1(n_398),
.B2(n_383),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_433),
.A2(n_436),
.B1(n_37),
.B2(n_35),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_434),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_418),
.A2(n_406),
.B(n_409),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_435),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_417),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_401),
.Y(n_438)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_438),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_432),
.A2(n_405),
.B1(n_14),
.B2(n_4),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_442),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_443),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_429),
.A2(n_14),
.B(n_12),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_28),
.C(n_34),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_447),
.C(n_423),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_435),
.A2(n_5),
.B(n_28),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_0),
.B(n_1),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_438),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_456),
.B1(n_437),
.B2(n_442),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_439),
.A2(n_430),
.B(n_425),
.Y(n_451)
);

AOI21x1_ASAP7_75t_L g462 ( 
.A1(n_451),
.A2(n_452),
.B(n_455),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_449),
.A2(n_422),
.B(n_426),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_442),
.Y(n_461)
);

A2O1A1O1Ixp25_ASAP7_75t_L g455 ( 
.A1(n_444),
.A2(n_433),
.B(n_5),
.C(n_35),
.D(n_37),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_448),
.C(n_440),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_459),
.B(n_460),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_447),
.C(n_443),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_461),
.A2(n_462),
.B(n_458),
.Y(n_465)
);

NAND2x1_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_464),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_458),
.A2(n_445),
.B(n_35),
.Y(n_464)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_465),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_461),
.A2(n_455),
.B(n_1),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_1),
.B(n_34),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_467),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_466),
.B(n_469),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_34),
.Y(n_473)
);


endmodule