module real_jpeg_31377_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_6;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_13),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_11),
.Y(n_10)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AOI211xp5_ASAP7_75t_L g5 ( 
.A1(n_6),
.A2(n_14),
.B(n_21),
.C(n_25),
.Y(n_5)
);

AOI22xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_13),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_15),
.B1(n_19),
.B2(n_20),
.Y(n_14)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_23),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_18),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);


endmodule