module fake_jpeg_11898_n_394 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_0),
.CON(n_57),
.SN(n_57)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_77),
.B(n_0),
.Y(n_113)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_64),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_15),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_71),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_39),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_1),
.Y(n_77)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_92),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_14),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_1),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_25),
.B(n_2),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_101),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_108),
.Y(n_159)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_32),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_47),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_3),
.B(n_12),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_42),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_44),
.B(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_3),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_23),
.B(n_14),
.C(n_12),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_50),
.C(n_45),
.Y(n_160)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_97),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_113),
.B(n_175),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_46),
.B1(n_28),
.B2(n_42),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_121),
.A2(n_125),
.B1(n_130),
.B2(n_170),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_124),
.A2(n_130),
.B(n_142),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_58),
.A2(n_46),
.B1(n_28),
.B2(n_42),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_127),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_59),
.A2(n_47),
.B1(n_53),
.B2(n_24),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_133),
.A2(n_162),
.B1(n_152),
.B2(n_150),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_54),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_134),
.B(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_51),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_91),
.A2(n_38),
.B1(n_49),
.B2(n_24),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_77),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_153),
.B(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_93),
.A2(n_38),
.B1(n_26),
.B2(n_49),
.Y(n_162)
);

INVx2_ASAP7_75t_R g164 ( 
.A(n_57),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_66),
.B(n_26),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_34),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_81),
.A2(n_53),
.B1(n_34),
.B2(n_40),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_173),
.B1(n_73),
.B2(n_87),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_40),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_145),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_68),
.A2(n_0),
.B1(n_29),
.B2(n_106),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_83),
.B(n_80),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_171),
.Y(n_194)
);

OR2x2_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_80),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_R g233 ( 
.A(n_176),
.B(n_184),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_61),
.C(n_63),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_202),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_179),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_180),
.A2(n_181),
.B1(n_195),
.B2(n_222),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_73),
.B1(n_79),
.B2(n_82),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_117),
.A2(n_86),
.B1(n_88),
.B2(n_94),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_199),
.B1(n_181),
.B2(n_178),
.Y(n_238)
);

NAND2x1_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_87),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_185),
.Y(n_248)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_194),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_227),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_197),
.A2(n_214),
.B1(n_218),
.B2(n_202),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_136),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_200),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_121),
.A2(n_125),
.B1(n_159),
.B2(n_175),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_146),
.B(n_112),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_203),
.B(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_114),
.B(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_126),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_211),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_131),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_216),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_144),
.B1(n_116),
.B2(n_123),
.Y(n_214)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_215),
.Y(n_230)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_116),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_217),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_144),
.A2(n_123),
.B1(n_152),
.B2(n_143),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_122),
.B(n_151),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_219),
.B(n_220),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_122),
.B(n_151),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_147),
.B(n_148),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_221),
.B(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_151),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_147),
.B(n_148),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_228),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_154),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_154),
.A2(n_161),
.B1(n_153),
.B2(n_164),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_184),
.B1(n_176),
.B2(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_236),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_182),
.B1(n_180),
.B2(n_195),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_177),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_240),
.B(n_256),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_183),
.B1(n_201),
.B2(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_250),
.B1(n_254),
.B2(n_268),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_201),
.B1(n_226),
.B2(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_188),
.B(n_192),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_212),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_260),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_189),
.B(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_196),
.B(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_189),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_230),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_179),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_249),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_179),
.A2(n_228),
.B1(n_199),
.B2(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_288),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_244),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_269),
.B1(n_252),
.B2(n_238),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_258),
.B1(n_267),
.B2(n_266),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_234),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_282),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_292),
.C(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_295),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_239),
.B(n_253),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_246),
.B(n_235),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_301),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_264),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_247),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_263),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_249),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_298),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_260),
.B(n_236),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_299),
.A2(n_266),
.B(n_271),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_243),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_275),
.C(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_309),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_242),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.C(n_275),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_242),
.B1(n_230),
.B2(n_261),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_313),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_277),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_316),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_258),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_324),
.B1(n_291),
.B2(n_283),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_287),
.A2(n_270),
.B1(n_231),
.B2(n_237),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_321),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_292),
.C(n_275),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_331),
.C(n_338),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_300),
.Y(n_331)
);

OAI322xp33_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_273),
.A3(n_280),
.B1(n_294),
.B2(n_288),
.C1(n_276),
.C2(n_299),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_332),
.B(n_340),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_273),
.C(n_280),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_314),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g334 ( 
.A1(n_323),
.A2(n_290),
.B1(n_289),
.B2(n_279),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_336),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_310),
.A2(n_278),
.B(n_245),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_278),
.B(n_310),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_301),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_341),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_315),
.B1(n_313),
.B2(n_309),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_349),
.C(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_303),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_339),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_330),
.A2(n_306),
.B1(n_316),
.B2(n_317),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_352),
.A2(n_325),
.B1(n_329),
.B2(n_341),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_338),
.C(n_326),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_334),
.A2(n_304),
.B1(n_310),
.B2(n_324),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_355),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_363)
);

AOI31xp67_ASAP7_75t_L g357 ( 
.A1(n_351),
.A2(n_304),
.A3(n_326),
.B(n_334),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_358),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_331),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_345),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_364),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_350),
.B1(n_344),
.B2(n_322),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_366),
.C(n_352),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_363),
.A2(n_355),
.B1(n_347),
.B2(n_343),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_367),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_354),
.B(n_353),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_342),
.A2(n_319),
.B(n_272),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_365),
.C(n_367),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_349),
.C(n_342),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_372),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_318),
.B(n_286),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_360),
.A2(n_343),
.B1(n_350),
.B2(n_344),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_373),
.B(n_375),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_297),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_379),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_372),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_381),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_384),
.A2(n_386),
.B(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_376),
.C(n_368),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_385),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_373),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_389),
.C(n_383),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_318),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g391 ( 
.A1(n_388),
.A2(n_369),
.B(n_271),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_391),
.A2(n_270),
.B(n_255),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.Y(n_394)
);


endmodule