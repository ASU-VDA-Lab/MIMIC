module fake_jpeg_31131_n_536 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_536);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_62),
.B(n_65),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_68),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_90),
.Y(n_130)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_2),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_88),
.Y(n_108)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_29),
.B(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_2),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_102),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_99),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_103),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_50),
.C(n_31),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_107),
.B(n_140),
.C(n_2),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_62),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_125),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_40),
.C(n_24),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_56),
.B(n_38),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_152),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_63),
.A2(n_44),
.B1(n_34),
.B2(n_38),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_40),
.B1(n_46),
.B2(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_42),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_42),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_32),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_80),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_91),
.B(n_52),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_52),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_76),
.A2(n_51),
.B1(n_44),
.B2(n_30),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_94),
.B1(n_51),
.B2(n_44),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_168),
.A2(n_212),
.B(n_133),
.Y(n_232)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_124),
.A2(n_82),
.B1(n_78),
.B2(n_30),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_179),
.B1(n_191),
.B2(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_176),
.B(n_184),
.Y(n_247)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_105),
.B1(n_104),
.B2(n_89),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_116),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_108),
.B(n_80),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_145),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_37),
.Y(n_188)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_116),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_193),
.A2(n_199),
.B1(n_207),
.B2(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_79),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_194),
.B(n_201),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_195),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_139),
.B1(n_118),
.B2(n_112),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_204),
.B1(n_150),
.B2(n_156),
.Y(n_240)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_142),
.A2(n_79),
.B1(n_73),
.B2(n_61),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_135),
.A2(n_77),
.B1(n_73),
.B2(n_61),
.Y(n_200)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_99),
.B1(n_32),
.B2(n_6),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_123),
.A2(n_32),
.B1(n_5),
.B2(n_7),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_214),
.Y(n_249)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_218),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_136),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_5),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_120),
.B(n_5),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_139),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_210),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_174),
.A2(n_144),
.B1(n_160),
.B2(n_156),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g286 ( 
.A1(n_226),
.A2(n_242),
.B1(n_212),
.B2(n_137),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_125),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_243),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_240),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_232),
.B(n_249),
.Y(n_263)
);

AOI22x1_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_163),
.B1(n_115),
.B2(n_165),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_151),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_146),
.C(n_111),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_180),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_167),
.A2(n_115),
.B(n_155),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_167),
.B(n_180),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_168),
.A2(n_121),
.B(n_122),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_260),
.B(n_167),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_198),
.A2(n_121),
.B(n_143),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_251),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_263),
.A2(n_265),
.B(n_237),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_220),
.A2(n_160),
.B1(n_150),
.B2(n_191),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_264),
.A2(n_214),
.B1(n_206),
.B2(n_203),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_208),
.B1(n_210),
.B2(n_172),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_266),
.A2(n_259),
.B1(n_238),
.B2(n_234),
.Y(n_311)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_236),
.B(n_224),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_187),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_189),
.B1(n_179),
.B2(n_177),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_286),
.B1(n_236),
.B2(n_231),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_285),
.B(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_198),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_275),
.B(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_229),
.B(n_183),
.Y(n_278)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_197),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_281),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_186),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_282),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_208),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_202),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_229),
.B(n_182),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_292),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_227),
.B(n_209),
.Y(n_292)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_253),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_261),
.B(n_227),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_296),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_211),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_260),
.B(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_189),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_324),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_298),
.B(n_286),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_255),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_305),
.C(n_333),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_255),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_310),
.A2(n_316),
.B1(n_328),
.B2(n_270),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_314),
.A2(n_318),
.B1(n_325),
.B2(n_270),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_272),
.A2(n_242),
.B1(n_234),
.B2(n_254),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_264),
.A2(n_242),
.B1(n_178),
.B2(n_169),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_320),
.B(n_323),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_275),
.B(n_258),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_283),
.A2(n_259),
.B1(n_238),
.B2(n_195),
.Y(n_325)
);

XOR2x2_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_257),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_327),
.B(n_279),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_223),
.B1(n_246),
.B2(n_245),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g356 ( 
.A1(n_329),
.A2(n_291),
.B(n_278),
.C(n_290),
.D(n_284),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_245),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_256),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_363),
.B1(n_325),
.B2(n_314),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_307),
.A2(n_286),
.B(n_273),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_355),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_269),
.B(n_265),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_336),
.A2(n_347),
.B(n_356),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_337),
.B(n_354),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_342),
.B1(n_343),
.B2(n_367),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_285),
.B1(n_295),
.B2(n_286),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_285),
.B1(n_286),
.B2(n_262),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_280),
.C(n_292),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_299),
.C(n_320),
.Y(n_373)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_349),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_329),
.A2(n_296),
.B(n_267),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_357),
.B(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_308),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_353),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_293),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_274),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_276),
.B(n_293),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_308),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_364),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_359),
.B(n_316),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_279),
.Y(n_360)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_366),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_282),
.Y(n_362)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_282),
.B1(n_268),
.B2(n_235),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_268),
.B(n_246),
.Y(n_365)
);

INVx6_ASAP7_75t_SL g366 ( 
.A(n_301),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_305),
.A2(n_235),
.B1(n_277),
.B2(n_216),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_360),
.B(n_315),
.Y(n_369)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_306),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_382),
.C(n_392),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_376),
.A2(n_383),
.B1(n_338),
.B2(n_343),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_322),
.Y(n_377)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_377),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_333),
.C(n_332),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_338),
.A2(n_327),
.B1(n_311),
.B2(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_322),
.Y(n_385)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_315),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_360),
.B(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_391),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_355),
.B(n_331),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_328),
.C(n_326),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_336),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_340),
.B(n_303),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_303),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_397),
.B(n_335),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_399),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_326),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_401),
.A2(n_410),
.B1(n_388),
.B2(n_375),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_363),
.B1(n_369),
.B2(n_390),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_402),
.A2(n_424),
.B1(n_372),
.B2(n_309),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_406),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_407),
.B(n_416),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_373),
.B(n_345),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_422),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_393),
.A2(n_335),
.B(n_351),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_409),
.A2(n_384),
.B(n_379),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_339),
.B1(n_341),
.B2(n_367),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_368),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_393),
.A2(n_387),
.B(n_398),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_429),
.Y(n_436)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_347),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_359),
.C(n_357),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_426),
.C(n_427),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_383),
.A2(n_334),
.B1(n_356),
.B2(n_361),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_419),
.A2(n_381),
.B1(n_387),
.B2(n_378),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_352),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_381),
.A2(n_350),
.B1(n_364),
.B2(n_319),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_319),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_377),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_313),
.C(n_301),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_309),
.C(n_216),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_387),
.A2(n_349),
.B(n_346),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_435),
.Y(n_454)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_415),
.Y(n_434)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_400),
.C(n_385),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_439),
.C(n_453),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_400),
.C(n_399),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_370),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_442),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_368),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_443),
.Y(n_462)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_444),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_445),
.A2(n_409),
.B(n_417),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_376),
.B1(n_379),
.B2(n_374),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_449),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_452),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_423),
.B(n_375),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_451),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_374),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_372),
.C(n_277),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_413),
.B(n_429),
.Y(n_455)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_468),
.Y(n_473)
);

XOR2x2_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_422),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_433),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_427),
.C(n_407),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_472),
.C(n_438),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_417),
.B(n_414),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_439),
.B(n_420),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_451),
.Y(n_481)
);

BUFx12_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_419),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_424),
.C(n_425),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_475),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_433),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_453),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_477),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_440),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_441),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_482),
.Y(n_498)
);

AOI31xp33_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_405),
.A3(n_442),
.B(n_421),
.Y(n_479)
);

OAI21x1_ASAP7_75t_SL g494 ( 
.A1(n_479),
.A2(n_457),
.B(n_468),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_430),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_483),
.B(n_484),
.Y(n_492)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_490),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_438),
.C(n_401),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_11),
.C(n_12),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_128),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_460),
.B(n_8),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_472),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_467),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_456),
.A2(n_117),
.B(n_137),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_480),
.A2(n_466),
.B(n_457),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_491),
.A2(n_495),
.B(n_11),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_494),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_483),
.A2(n_470),
.B(n_463),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_500),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_473),
.A2(n_458),
.B1(n_471),
.B2(n_467),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_476),
.B(n_9),
.Y(n_501)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

MAJx2_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_9),
.C(n_10),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_13),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_503),
.B(n_12),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_492),
.C(n_498),
.Y(n_506)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_493),
.A2(n_473),
.B(n_482),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_504),
.A2(n_477),
.B(n_475),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_508),
.B(n_511),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_510),
.B(n_512),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_11),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_513),
.B(n_515),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_13),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_493),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_517),
.B(n_505),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_506),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_514),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_526),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_519),
.A2(n_512),
.B(n_503),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_527),
.B(n_523),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_521),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_531),
.C(n_509),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_529),
.C(n_522),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_520),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_505),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_13),
.Y(n_536)
);


endmodule