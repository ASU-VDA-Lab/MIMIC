module fake_jpeg_22579_n_271 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_61),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.C(n_25),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_68),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_24),
.Y(n_64)
);

AO22x2_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_37),
.B1(n_34),
.B2(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_19),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_32),
.B1(n_21),
.B2(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_77),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_44),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_100),
.C(n_86),
.Y(n_114)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_52),
.B1(n_58),
.B2(n_56),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_103),
.B1(n_56),
.B2(n_42),
.Y(n_121)
);

AO21x1_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_65),
.B(n_44),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_60),
.B1(n_78),
.B2(n_48),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_54),
.B1(n_58),
.B2(n_40),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_85),
.B1(n_52),
.B2(n_75),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_0),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_53),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_54),
.B1(n_40),
.B2(n_39),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_51),
.B(n_55),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_87),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_69),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_90),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_118),
.B1(n_120),
.B2(n_123),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_97),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_84),
.B1(n_75),
.B2(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_82),
.C(n_41),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_102),
.B1(n_99),
.B2(n_96),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_125),
.B1(n_134),
.B2(n_92),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_87),
.B1(n_74),
.B2(n_69),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_131),
.B(n_21),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_87),
.B1(n_74),
.B2(n_49),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_94),
.B1(n_46),
.B2(n_106),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_22),
.B(n_24),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_27),
.B1(n_22),
.B2(n_16),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_34),
.C(n_48),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_143),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_154),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_110),
.B1(n_105),
.B2(n_100),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_158),
.B(n_160),
.Y(n_170)
);

OAI22x1_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_94),
.B1(n_100),
.B2(n_97),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_100),
.B1(n_98),
.B2(n_90),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_161),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_107),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_113),
.B1(n_112),
.B2(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_149),
.B1(n_154),
.B2(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_45),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_128),
.B(n_79),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_111),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_169),
.B1(n_174),
.B2(n_186),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_115),
.B1(n_133),
.B2(n_126),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_171),
.B1(n_151),
.B2(n_144),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_176),
.C(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_133),
.B1(n_122),
.B2(n_126),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_122),
.B1(n_26),
.B2(n_20),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_45),
.B1(n_79),
.B2(n_46),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_128),
.C(n_45),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_185),
.B(n_147),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_0),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_31),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_128),
.B(n_79),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_153),
.B1(n_160),
.B2(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_176),
.C(n_167),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_165),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_196),
.B(n_199),
.Y(n_219)
);

OAI31xp33_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_158),
.A3(n_151),
.B(n_161),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_203),
.B1(n_171),
.B2(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_151),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_205),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_10),
.C(n_15),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_20),
.B1(n_0),
.B2(n_1),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_170),
.C(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_170),
.C(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_213),
.B(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_178),
.B1(n_179),
.B2(n_1),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_31),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_5),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_204),
.B1(n_193),
.B2(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_196),
.B(n_2),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_229),
.B(n_232),
.Y(n_241)
);

AO221x1_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_31),
.B1(n_1),
.B2(n_3),
.C(n_4),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_227),
.B(n_236),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_1),
.B(n_15),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_2),
.B(n_4),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_4),
.B(n_5),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_11),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_7),
.B(n_10),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_246),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_223),
.B(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_244),
.B(n_13),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_220),
.B1(n_217),
.B2(n_208),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_224),
.B1(n_227),
.B2(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_12),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_221),
.C(n_215),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_13),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_11),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_231),
.B1(n_230),
.B2(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_250),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_252),
.B(n_237),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_212),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_253),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_254),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_241),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_238),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_264),
.B(n_258),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_263),
.B(n_247),
.C(n_14),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_268),
.B(n_13),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_269),
.B(n_14),
.CI(n_241),
.CON(n_270),
.SN(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_14),
.Y(n_271)
);


endmodule