module real_jpeg_11232_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_310, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_310;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_143),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_3),
.A2(n_27),
.B1(n_35),
.B2(n_143),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_45),
.B(n_56),
.C(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_32),
.B(n_43),
.C(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_9),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_152),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_9),
.A2(n_27),
.B1(n_35),
.B2(n_152),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_10),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_10),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_11),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_12),
.A2(n_27),
.B1(n_35),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_91),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_91),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_91),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_62),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_15),
.A2(n_45),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_45),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_15),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_81),
.B1(n_84),
.B2(n_161),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_32),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_15),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_15),
.A2(n_29),
.B(n_33),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_15),
.A2(n_27),
.B1(n_35),
.B2(n_163),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_16),
.A2(n_27),
.B1(n_35),
.B2(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_16),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_17),
.A2(n_27),
.B1(n_35),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_125),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_125),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_64),
.C(n_77),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_23),
.A2(n_64),
.B1(n_65),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_23),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_24),
.A2(n_25),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_53),
.C(n_63),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_26),
.A2(n_31),
.B1(n_37),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_26),
.A2(n_31),
.B1(n_90),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_26),
.A2(n_31),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_26),
.A2(n_31),
.B1(n_124),
.B2(n_259),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_28),
.B(n_163),
.C(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_31),
.Y(n_208)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_42),
.A2(n_44),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_42),
.A2(n_44),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_42),
.A2(n_44),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_44),
.B1(n_188),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_42),
.A2(n_44),
.B1(n_204),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_42),
.A2(n_44),
.B1(n_243),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_42),
.A2(n_44),
.B1(n_128),
.B2(n_255),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_44),
.B(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_45),
.B(n_47),
.Y(n_192)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_46),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_54),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_57),
.B1(n_73),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_55),
.A2(n_57),
.B1(n_87),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_55),
.A2(n_57),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_55),
.A2(n_57),
.B1(n_151),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_55),
.A2(n_57),
.B1(n_176),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_55),
.A2(n_57),
.B1(n_184),
.B2(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_55),
.A2(n_57),
.B1(n_121),
.B2(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_56),
.Y(n_156)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_57),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_58),
.B(n_60),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_58),
.B(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_59),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_66),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_74),
.A2(n_76),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_88),
.B(n_89),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_79),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_88),
.B1(n_89),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_290),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_85),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_81),
.A2(n_84),
.B1(n_142),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_81),
.A2(n_84),
.B1(n_145),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_81),
.A2(n_84),
.B1(n_178),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_81),
.A2(n_84),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_81),
.A2(n_84),
.B1(n_119),
.B2(n_231),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_83),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_82),
.A2(n_83),
.B1(n_196),
.B2(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_163),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_86),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_132),
.B(n_308),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_129),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_108),
.B(n_129),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_115),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_109),
.Y(n_295)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_115),
.A2(n_116),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_126),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_117),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_118),
.B(n_120),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI321xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_284),
.A3(n_296),
.B1(n_302),
.B2(n_307),
.C(n_310),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_249),
.C(n_280),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_220),
.B(n_248),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_198),
.B(n_219),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_180),
.B(n_197),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_170),
.B(n_179),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_158),
.B(n_169),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_157),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_157),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_171),
.B(n_172),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.C(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.CI(n_189),
.CON(n_182),
.SN(n_182)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_194),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_199),
.B(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_212),
.B2(n_213),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_215),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_211),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_222),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_235),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_224),
.B(n_234),
.C(n_235),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_244),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_241),
.C(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_250),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_251),
.B(n_267),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.C(n_266),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_261),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_256),
.B1(n_257),
.B2(n_260),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_266),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_264),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_278),
.B2(n_279),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_271),
.C(n_279),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_282),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);


endmodule