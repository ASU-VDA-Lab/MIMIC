module real_jpeg_5198_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_0),
.B(n_61),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_0),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_0),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_0),
.B(n_307),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_0),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_0),
.B(n_399),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_0),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_1),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_1),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_1),
.B(n_105),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_1),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_1),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_1),
.B(n_426),
.Y(n_425)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_2),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_2),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_3),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_3),
.B(n_91),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_108),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_3),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_328),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_3),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_4),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_4),
.B(n_61),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_4),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_4),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_4),
.B(n_284),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_4),
.B(n_423),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_6),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_6),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_6),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_7),
.B(n_68),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_7),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_7),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_7),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_7),
.B(n_273),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_9),
.Y(n_544)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_10),
.Y(n_301)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_12),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_13),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_13),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_13),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_13),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_13),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_13),
.B(n_115),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_13),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_13),
.B(n_420),
.Y(n_419)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_14),
.Y(n_547)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_16),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_16),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_16),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_16),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_16),
.B(n_140),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_16),
.B(n_397),
.Y(n_396)
);

AND2x4_ASAP7_75t_SL g412 ( 
.A(n_16),
.B(n_413),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_17),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_17),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_17),
.B(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_19),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_19),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_19),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_19),
.B(n_140),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_19),
.B(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_542),
.B(n_545),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_43),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_30),
.B1(n_37),
.B2(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_47),
.C(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_32),
.Y(n_397)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_33),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_33),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_72),
.C(n_74),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_44),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_62),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_45),
.B(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_54),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_47),
.A2(n_53),
.B1(n_67),
.B2(n_118),
.Y(n_122)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_49),
.Y(n_399)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_51),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_51),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_63),
.C(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_62),
.Y(n_125)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_64),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_67),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_514)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_69),
.Y(n_228)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_70),
.Y(n_368)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_71),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_71),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_71),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_129),
.B(n_541),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_126),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_79),
.B(n_126),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_123),
.C(n_124),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_80),
.A2(n_81),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_106),
.C(n_119),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_82),
.A2(n_83),
.B1(n_518),
.B2(n_520),
.Y(n_517)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_89),
.C(n_93),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_94),
.B(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_509)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_106),
.A2(n_119),
.B1(n_120),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_106),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_118),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_107),
.B(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_112),
.B1(n_207),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_112),
.B(n_204),
.C(n_207),
.Y(n_515)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_116),
.Y(n_331)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_117),
.Y(n_424)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_123),
.B(n_124),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_535),
.B(n_540),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_502),
.B(n_532),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_310),
.B(n_501),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_256),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_133),
.B(n_256),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_201),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_134),
.B(n_202),
.C(n_231),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_173),
.C(n_183),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_135),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.C(n_157),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_136),
.B(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_139),
.C(n_141),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_140),
.Y(n_288)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_144),
.A2(n_145),
.B1(n_157),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_154),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_146),
.B(n_154),
.Y(n_477)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_147),
.Y(n_414)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_149),
.B(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_153),
.Y(n_352)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_153),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_157),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_158),
.Y(n_242)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_164),
.B(n_169),
.C(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_168),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_169),
.A2(n_170),
.B1(n_207),
.B2(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_207),
.C(n_235),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_172),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_183),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_179),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_179),
.A2(n_181),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_180),
.C(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_179),
.B(n_248),
.C(n_252),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.C(n_198),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_184),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.C(n_192),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_185),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_187),
.B(n_192),
.Y(n_268)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_191),
.Y(n_343)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_191),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_194),
.B(n_198),
.Y(n_291)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_197),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_231),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_203),
.B(n_212),
.C(n_230),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_207),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_222),
.B1(n_229),
.B2(n_230),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.C(n_219),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_219),
.Y(n_244)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_223),
.B(n_225),
.C(n_226),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_245),
.B2(n_246),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_232),
.B(n_247),
.C(n_254),
.Y(n_527)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.C(n_243),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_258),
.B(n_261),
.Y(n_497)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_263),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_289),
.C(n_292),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_265),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_278),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_266),
.A2(n_267),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_269),
.A2(n_270),
.B(n_274),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_269),
.B(n_278),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.C(n_286),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_445)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_286),
.B(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_287),
.B(n_308),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_292),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_306),
.C(n_309),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_294),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_302),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_295),
.B(n_457),
.Y(n_456)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_298),
.A2(n_302),
.B1(n_303),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_298),
.Y(n_458)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_306),
.B(n_309),
.Y(n_479)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_495),
.B(n_500),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_482),
.B(n_494),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_464),
.B(n_481),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_438),
.B(n_463),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_403),
.B(n_437),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_374),
.B(n_402),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_354),
.B(n_373),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_337),
.B(n_353),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_332),
.B(n_336),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_326),
.Y(n_338)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_339),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_346),
.B2(n_347),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_349),
.C(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_372),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_372),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_363),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_363),
.C(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_361),
.Y(n_379)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_389),
.C(n_390),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_377),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_378),
.B(n_388),
.C(n_391),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_381),
.C(n_382),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_382)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_386),
.Y(n_407)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_398),
.C(n_400),
.Y(n_435)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.Y(n_395)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_396),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_398),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_436),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_436),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_416),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_406),
.B(n_415),
.C(n_462),
.Y(n_461)
);

XNOR2x1_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_452),
.C(n_453),
.Y(n_451)
);

XNOR2x1_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_412),
.Y(n_408)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_412),
.Y(n_453)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_427),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_429),
.C(n_434),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_422),
.C(n_425),
.Y(n_449)
);

INVx6_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_434),
.B2(n_435),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_433),
.Y(n_448)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_461),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_461),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_450),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_442),
.C(n_450),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_447),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_473),
.C(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_448),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_455),
.C(n_460),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_459),
.B2(n_460),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_480),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_480),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_470),
.C(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_476),
.C(n_478),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_492),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_492),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_489),
.C(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_498),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_528),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g532 ( 
.A1(n_503),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_522),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_522),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_511),
.B2(n_521),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_512),
.C(n_517),
.Y(n_539)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.C(n_510),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_524),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_510),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_511),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_517),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_515),
.C(n_516),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_516),
.Y(n_526)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_518),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.C(n_527),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_525),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_530),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_531),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_536),
.B(n_539),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_539),
.Y(n_540)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx13_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_544),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);


endmodule