module fake_jpeg_12621_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_51),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_48),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_53),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_62),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_67),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_93),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_65),
.B1(n_56),
.B2(n_58),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_71),
.B1(n_58),
.B2(n_61),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_92),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_55),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_104),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_4),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_99),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_81),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_50),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_102),
.B(n_3),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_115),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_116),
.Y(n_121)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_64),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_64),
.C(n_28),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_136),
.C(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_24),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_25),
.B(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_14),
.B1(n_16),
.B2(n_19),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_32),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_115),
.C(n_106),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_20),
.C(n_21),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_147),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_22),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_131),
.B1(n_119),
.B2(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_148),
.B1(n_127),
.B2(n_120),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_29),
.B(n_30),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_157),
.B(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_140),
.B1(n_137),
.B2(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_156),
.C(n_150),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

AO221x1_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_124),
.B1(n_125),
.B2(n_146),
.C(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_160),
.A2(n_153),
.B1(n_154),
.B2(n_138),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_161),
.B(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_162),
.B(n_163),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_38),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_39),
.Y(n_168)
);


endmodule