module real_aes_15538_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g37 ( .A(n_1), .Y(n_37) );
AOI21xp33_ASAP7_75t_SL g9 ( .A1(n_2), .A2(n_10), .B(n_23), .Y(n_9) );
INVx2_ASAP7_75t_L g41 ( .A(n_3), .Y(n_41) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_5), .Y(n_18) );
INVx1_ASAP7_75t_L g22 ( .A(n_6), .Y(n_22) );
INVx2_ASAP7_75t_L g40 ( .A(n_7), .Y(n_40) );
BUFx3_ASAP7_75t_L g33 ( .A(n_8), .Y(n_33) );
INVxp67_ASAP7_75t_SL g10 ( .A(n_11), .Y(n_10) );
NOR2xp33_ASAP7_75t_SL g11 ( .A(n_12), .B(n_19), .Y(n_11) );
INVxp33_ASAP7_75t_SL g12 ( .A(n_13), .Y(n_12) );
NOR3xp33_ASAP7_75t_L g13 ( .A(n_14), .B(n_17), .C(n_18), .Y(n_13) );
INVx2_ASAP7_75t_SL g14 ( .A(n_15), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g27 ( .A(n_17), .Y(n_27) );
INVx1_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_21), .B(n_27), .Y(n_26) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
INVx2_ASAP7_75t_SL g23 ( .A(n_24), .Y(n_23) );
OR2x6_ASAP7_75t_L g24 ( .A(n_25), .B(n_28), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
AND2x2_ASAP7_75t_L g28 ( .A(n_29), .B(n_42), .Y(n_28) );
NAND3xp33_ASAP7_75t_L g29 ( .A(n_30), .B(n_34), .C(n_38), .Y(n_29) );
AND2x6_ASAP7_75t_L g43 ( .A(n_30), .B(n_44), .Y(n_43) );
INVx3_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
BUFx6f_ASAP7_75t_L g32 ( .A(n_33), .Y(n_32) );
INVx2_ASAP7_75t_SL g34 ( .A(n_35), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
INVx3_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
BUFx2_ASAP7_75t_L g38 ( .A(n_39), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g39 ( .A(n_40), .B(n_41), .Y(n_39) );
INVx1_ASAP7_75t_L g46 ( .A(n_40), .Y(n_46) );
INVx3_ASAP7_75t_L g45 ( .A(n_41), .Y(n_45) );
INVx4_ASAP7_75t_L g42 ( .A(n_43), .Y(n_42) );
AND2x4_ASAP7_75t_L g44 ( .A(n_45), .B(n_46), .Y(n_44) );
endmodule