module fake_netlist_6_1023_n_1146 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1146);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1146;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_1078;
wire n_314;
wire n_923;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_844;
wire n_953;
wire n_1017;
wire n_1094;
wire n_1004;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1041;
wire n_279;
wire n_686;
wire n_796;
wire n_1000;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_1075;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_267;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_70),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_81),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_67),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_154),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_202),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_163),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_116),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_82),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_49),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_32),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_131),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_91),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_47),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_103),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_80),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_21),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_21),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_113),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_60),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_196),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_177),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_153),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_99),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_191),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_166),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_184),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_110),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_76),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_107),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_135),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_28),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_159),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_102),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_133),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_104),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_210),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_117),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_171),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_54),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_243),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_229),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_254),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_232),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_223),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_263),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_226),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_249),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_230),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_227),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_336),
.Y(n_344)
);

CKINVDCx6p67_ASAP7_75t_R g345 ( 
.A(n_331),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_336),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_231),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

CKINVDCx11_ASAP7_75t_R g351 ( 
.A(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_340),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_228),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_290),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_338),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_293),
.A2(n_281),
.B1(n_224),
.B2(n_262),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_293),
.A2(n_262),
.B1(n_284),
.B2(n_283),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_292),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_234),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_297),
.A2(n_246),
.B1(n_286),
.B2(n_282),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_33),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_342),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_241),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_312),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_327),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_289),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_297),
.A2(n_279),
.B1(n_277),
.B2(n_276),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_292),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_321),
.B(n_242),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_302),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_294),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_302),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_332),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_351),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_376),
.B(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_L g403 ( 
.A1(n_374),
.A2(n_307),
.B1(n_308),
.B2(n_296),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_359),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_358),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_376),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_325),
.C(n_307),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_366),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_333),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_389),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_385),
.C(n_377),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_380),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_359),
.Y(n_429)
);

AO21x2_ASAP7_75t_L g430 ( 
.A1(n_380),
.A2(n_305),
.B(n_303),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_339),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_308),
.C(n_341),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_353),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

OA22x2_ASAP7_75t_L g440 ( 
.A1(n_391),
.A2(n_299),
.B1(n_305),
.B2(n_310),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_303),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_383),
.B(n_310),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_392),
.Y(n_447)
);

AO21x2_ASAP7_75t_L g448 ( 
.A1(n_392),
.A2(n_334),
.B(n_329),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_383),
.B(n_364),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_343),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_346),
.B(n_329),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_351),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_371),
.B(n_244),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_353),
.B(n_298),
.C(n_299),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_362),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_362),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_348),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

CKINVDCx6p67_ASAP7_75t_R g465 ( 
.A(n_345),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_371),
.B(n_247),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_345),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_346),
.B(n_294),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_362),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_348),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_394),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_409),
.B(n_362),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_250),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_363),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_339),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_413),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_417),
.Y(n_483)
);

XNOR2x2_ASAP7_75t_L g484 ( 
.A(n_429),
.B(n_0),
.Y(n_484)
);

OR2x6_ASAP7_75t_L g485 ( 
.A(n_410),
.B(n_347),
.Y(n_485)
);

XOR2x2_ASAP7_75t_L g486 ( 
.A(n_432),
.B(n_0),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_433),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_401),
.B(n_256),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_R g490 ( 
.A(n_436),
.B(n_2),
.Y(n_490)
);

NOR2x1p5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_258),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_401),
.B(n_260),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

XNOR2x2_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_2),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_430),
.B(n_363),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_468),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_440),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_433),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_399),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_464),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_411),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_428),
.A2(n_378),
.B(n_354),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_416),
.B(n_264),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_412),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_414),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_415),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_428),
.B(n_347),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_425),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_363),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_437),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_448),
.A2(n_355),
.B(n_354),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_448),
.B(n_363),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_418),
.B(n_355),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_408),
.B(n_375),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_444),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_445),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_445),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_446),
.A2(n_378),
.B(n_267),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_419),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_266),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_454),
.B(n_373),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_447),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_439),
.B(n_373),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_408),
.B(n_375),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_403),
.B(n_270),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_458),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_460),
.B(n_274),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_405),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_458),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_431),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_470),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_536),
.B(n_470),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_506),
.B(n_471),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_515),
.B(n_420),
.Y(n_563)
);

O2A1O1Ixp5_ASAP7_75t_L g564 ( 
.A1(n_473),
.A2(n_459),
.B(n_466),
.C(n_472),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_503),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_449),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_472),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_459),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_493),
.B(n_449),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_528),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_509),
.Y(n_572)
);

AOI221xp5_ASAP7_75t_L g573 ( 
.A1(n_554),
.A2(n_436),
.B1(n_275),
.B2(n_466),
.C(n_400),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_493),
.B(n_514),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_L g575 ( 
.A(n_476),
.B(n_488),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_552),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_507),
.B(n_439),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_497),
.B(n_420),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_497),
.B(n_420),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_554),
.B(n_543),
.C(n_520),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_487),
.B(n_469),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_481),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_509),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_441),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_488),
.B(n_424),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_480),
.A2(n_461),
.B(n_456),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_492),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_474),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_520),
.A2(n_452),
.B1(n_404),
.B2(n_462),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_485),
.A2(n_404),
.B1(n_450),
.B2(n_465),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_475),
.B(n_404),
.Y(n_593)
);

O2A1O1Ixp5_ASAP7_75t_L g594 ( 
.A1(n_519),
.A2(n_452),
.B(n_378),
.C(n_450),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_511),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_477),
.B(n_452),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_478),
.B(n_479),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_485),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_482),
.B(n_452),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_483),
.A2(n_452),
.B1(n_378),
.B2(n_463),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_424),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_489),
.B(n_452),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_495),
.A2(n_378),
.B1(n_375),
.B2(n_396),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_424),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_481),
.B(n_463),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_522),
.B(n_540),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_543),
.A2(n_463),
.B1(n_396),
.B2(n_390),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_496),
.A2(n_373),
.B1(n_396),
.B2(n_390),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_556),
.B(n_373),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_508),
.B(n_400),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_540),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_486),
.A2(n_396),
.B1(n_390),
.B2(n_375),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_534),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_510),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_501),
.B(n_3),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_502),
.B(n_390),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_557),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_518),
.A2(n_405),
.B1(n_453),
.B2(n_5),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_490),
.A2(n_453),
.B1(n_4),
.B2(n_6),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_531),
.B(n_3),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_4),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_505),
.B(n_35),
.Y(n_624)
);

AO22x1_ASAP7_75t_L g625 ( 
.A1(n_490),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_523),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_512),
.B(n_7),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_559),
.B(n_557),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_524),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_578),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_481),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_615),
.B(n_588),
.Y(n_634)
);

INVx6_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_626),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_565),
.Y(n_637)
);

AOI21xp33_ASAP7_75t_L g638 ( 
.A1(n_581),
.A2(n_526),
.B(n_525),
.Y(n_638)
);

NAND2x1p5_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_599),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_563),
.B(n_484),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_619),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_569),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_589),
.B(n_527),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

NOR2x1_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_491),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_SL g647 ( 
.A(n_573),
.B(n_541),
.C(n_516),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

NOR2x2_ASAP7_75t_L g649 ( 
.A(n_607),
.B(n_494),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_575),
.A2(n_558),
.B1(n_555),
.B2(n_553),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_571),
.B(n_529),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_584),
.Y(n_652)
);

AND2x6_ASAP7_75t_SL g653 ( 
.A(n_607),
.B(n_513),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_577),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_570),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_592),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_568),
.A2(n_539),
.B(n_530),
.C(n_532),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_595),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_603),
.B(n_498),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_598),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_627),
.A2(n_535),
.B1(n_538),
.B2(n_544),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_612),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_597),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_561),
.B(n_546),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_617),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_606),
.B(n_547),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_567),
.B(n_533),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_616),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_606),
.B(n_533),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_600),
.B(n_500),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_579),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_617),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_624),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_SL g678 ( 
.A(n_621),
.B(n_545),
.C(n_9),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_560),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_614),
.B(n_549),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_627),
.B(n_550),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_623),
.B(n_548),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_SL g684 ( 
.A(n_621),
.B(n_9),
.C(n_10),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_622),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_582),
.B(n_548),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_562),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_593),
.B(n_11),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_608),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_620),
.Y(n_690)
);

BUFx8_ASAP7_75t_SL g691 ( 
.A(n_596),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_614),
.B(n_12),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_585),
.B(n_36),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_620),
.B(n_13),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_654),
.B(n_609),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_670),
.A2(n_587),
.B(n_594),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_653),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_657),
.A2(n_594),
.B(n_564),
.Y(n_698)
);

AOI21xp33_ASAP7_75t_L g699 ( 
.A1(n_690),
.A2(n_604),
.B(n_601),
.Y(n_699)
);

OA21x2_ASAP7_75t_L g700 ( 
.A1(n_638),
.A2(n_564),
.B(n_611),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_666),
.B(n_605),
.Y(n_701)
);

AOI21x1_ASAP7_75t_SL g702 ( 
.A1(n_672),
.A2(n_625),
.B(n_591),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

NAND2x1_ASAP7_75t_L g704 ( 
.A(n_629),
.B(n_590),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_668),
.B(n_618),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_682),
.B(n_602),
.Y(n_706)
);

AOI21x1_ASAP7_75t_L g707 ( 
.A1(n_693),
.A2(n_610),
.B(n_605),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_693),
.A2(n_38),
.B(n_37),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_634),
.B(n_636),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_663),
.B(n_14),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_679),
.B(n_14),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_689),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_630),
.A2(n_40),
.B(n_39),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_644),
.A2(n_43),
.B(n_42),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_686),
.A2(n_45),
.B(n_44),
.Y(n_715)
);

OA21x2_ASAP7_75t_L g716 ( 
.A1(n_638),
.A2(n_48),
.B(n_46),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_675),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_631),
.Y(n_718)
);

OA21x2_ASAP7_75t_L g719 ( 
.A1(n_681),
.A2(n_51),
.B(n_50),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_663),
.B(n_15),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_15),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_650),
.A2(n_55),
.B(n_52),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_655),
.Y(n_723)
);

OAI21x1_ASAP7_75t_SL g724 ( 
.A1(n_687),
.A2(n_58),
.B(n_57),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_SL g725 ( 
.A1(n_647),
.A2(n_61),
.B(n_59),
.Y(n_725)
);

O2A1O1Ixp5_ASAP7_75t_L g726 ( 
.A1(n_688),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_726)
);

OA22x2_ASAP7_75t_L g727 ( 
.A1(n_692),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_635),
.Y(n_728)
);

OAI21x1_ASAP7_75t_SL g729 ( 
.A1(n_683),
.A2(n_134),
.B(n_219),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_650),
.A2(n_132),
.B(n_217),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_667),
.A2(n_130),
.B(n_216),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_632),
.B(n_19),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_652),
.Y(n_734)
);

NAND2x1p5_ASAP7_75t_L g735 ( 
.A(n_654),
.B(n_62),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_694),
.A2(n_19),
.B(n_20),
.C(n_22),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_641),
.B(n_20),
.Y(n_737)
);

AOI21x1_ASAP7_75t_L g738 ( 
.A1(n_660),
.A2(n_220),
.B(n_136),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_662),
.A2(n_648),
.B(n_637),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_662),
.A2(n_127),
.B(n_214),
.Y(n_740)
);

OA21x2_ASAP7_75t_L g741 ( 
.A1(n_658),
.A2(n_126),
.B(n_213),
.Y(n_741)
);

OA22x2_ASAP7_75t_L g742 ( 
.A1(n_655),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_659),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_642),
.Y(n_744)
);

AOI21x1_ASAP7_75t_SL g745 ( 
.A1(n_680),
.A2(n_24),
.B(n_25),
.Y(n_745)
);

OAI21x1_ASAP7_75t_SL g746 ( 
.A1(n_646),
.A2(n_139),
.B(n_211),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_659),
.B(n_640),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_651),
.A2(n_137),
.B(n_209),
.Y(n_748)
);

NOR2x1_ASAP7_75t_L g749 ( 
.A(n_633),
.B(n_63),
.Y(n_749)
);

CKINVDCx11_ASAP7_75t_R g750 ( 
.A(n_633),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_677),
.A2(n_125),
.B(n_208),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_656),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_661),
.A2(n_123),
.B(n_207),
.Y(n_753)
);

AO31x2_ASAP7_75t_L g754 ( 
.A1(n_665),
.A2(n_25),
.A3(n_26),
.B(n_27),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_628),
.B(n_26),
.Y(n_755)
);

AOI21xp33_ASAP7_75t_L g756 ( 
.A1(n_677),
.A2(n_27),
.B(n_28),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_671),
.A2(n_29),
.B1(n_31),
.B2(n_64),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_639),
.A2(n_143),
.B(n_65),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_673),
.A2(n_144),
.B(n_66),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_718),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_709),
.B(n_678),
.Y(n_761)
);

OAI21x1_ASAP7_75t_L g762 ( 
.A1(n_696),
.A2(n_691),
.B(n_649),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_736),
.A2(n_684),
.B(n_633),
.C(n_673),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_743),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_698),
.A2(n_653),
.B(n_677),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_701),
.A2(n_674),
.B(n_645),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_712),
.B(n_669),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_740),
.A2(n_674),
.A3(n_645),
.B(n_29),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_SL g770 ( 
.A1(n_755),
.A2(n_664),
.B1(n_674),
.B2(n_635),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_722),
.A2(n_645),
.B(n_69),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_747),
.B(n_215),
.Y(n_772)
);

BUFx4_ASAP7_75t_SL g773 ( 
.A(n_728),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_710),
.A2(n_68),
.B(n_71),
.C(n_72),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_723),
.B(n_206),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_730),
.A2(n_73),
.B(n_74),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_704),
.A2(n_700),
.B(n_759),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_SL g778 ( 
.A(n_726),
.B(n_75),
.C(n_77),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_706),
.A2(n_78),
.B1(n_79),
.B2(n_83),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_718),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_756),
.B(n_84),
.C(n_85),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_739),
.A2(n_86),
.B(n_87),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_732),
.B(n_88),
.Y(n_783)
);

AOI22x1_ASAP7_75t_L g784 ( 
.A1(n_695),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_705),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_727),
.B(n_96),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_205),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_699),
.A2(n_97),
.B(n_98),
.Y(n_788)
);

BUFx6f_ASAP7_75t_SL g789 ( 
.A(n_743),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_735),
.B(n_744),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_732),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_100),
.B(n_101),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_750),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_734),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_753),
.A2(n_105),
.B(n_106),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_707),
.A2(n_108),
.B(n_109),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_SL g797 ( 
.A1(n_720),
.A2(n_111),
.B(n_112),
.C(n_114),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_700),
.A2(n_204),
.B(n_118),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_713),
.A2(n_203),
.B(n_119),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_734),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_752),
.Y(n_801)
);

OAI21x1_ASAP7_75t_SL g802 ( 
.A1(n_746),
.A2(n_115),
.B(n_120),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_721),
.B(n_201),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_731),
.A2(n_121),
.B(n_122),
.Y(n_805)
);

NOR2x1_ASAP7_75t_R g806 ( 
.A(n_697),
.B(n_140),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_SL g807 ( 
.A1(n_757),
.A2(n_141),
.B(n_145),
.C(n_146),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_714),
.A2(n_147),
.B(n_148),
.C(n_149),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_725),
.A2(n_200),
.B(n_152),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_SL g810 ( 
.A1(n_749),
.A2(n_151),
.B(n_155),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_738),
.A2(n_157),
.B(n_158),
.Y(n_811)
);

BUFx12f_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_703),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_715),
.A2(n_198),
.B(n_161),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_748),
.A2(n_160),
.B(n_164),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_165),
.B(n_167),
.C(n_168),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_703),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_697),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_741),
.A2(n_197),
.B(n_175),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_754),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_697),
.B(n_173),
.Y(n_821)
);

AOI31xp67_ASAP7_75t_L g822 ( 
.A1(n_745),
.A2(n_176),
.A3(n_178),
.B(n_179),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_SL g823 ( 
.A(n_733),
.B(n_180),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_L g824 ( 
.A(n_737),
.B(n_181),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_742),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_741),
.A2(n_719),
.B(n_716),
.Y(n_827)
);

AOI21xp33_ASAP7_75t_L g828 ( 
.A1(n_724),
.A2(n_182),
.B(n_183),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_765),
.B(n_719),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_791),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_761),
.A2(n_716),
.B1(n_702),
.B2(n_754),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_760),
.Y(n_832)
);

CKINVDCx6p67_ASAP7_75t_R g833 ( 
.A(n_789),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_780),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_800),
.B(n_754),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_823),
.A2(n_729),
.B1(n_186),
.B2(n_187),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_804),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_794),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_801),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_789),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_767),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_817),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_812),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_786),
.A2(n_185),
.B1(n_188),
.B2(n_192),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_820),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_770),
.A2(n_193),
.B1(n_194),
.B2(n_810),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_764),
.Y(n_847)
);

INVx6_ASAP7_75t_L g848 ( 
.A(n_764),
.Y(n_848)
);

BUFx8_ASAP7_75t_SL g849 ( 
.A(n_793),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_SL g851 ( 
.A1(n_825),
.A2(n_784),
.B1(n_788),
.B2(n_781),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_SL g852 ( 
.A1(n_805),
.A2(n_815),
.B1(n_818),
.B2(n_785),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_764),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_769),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_824),
.A2(n_778),
.B1(n_772),
.B2(n_779),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_762),
.B(n_826),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_773),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_768),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_779),
.A2(n_763),
.B1(n_824),
.B2(n_787),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_790),
.Y(n_860)
);

BUFx12f_ASAP7_75t_L g861 ( 
.A(n_790),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_775),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_806),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_SL g864 ( 
.A1(n_774),
.A2(n_809),
.B(n_828),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_769),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_777),
.Y(n_866)
);

INVx6_ASAP7_75t_L g867 ( 
.A(n_806),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_822),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_803),
.Y(n_869)
);

INVx6_ASAP7_75t_L g870 ( 
.A(n_766),
.Y(n_870)
);

CKINVDCx11_ASAP7_75t_R g871 ( 
.A(n_821),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_782),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_799),
.A2(n_814),
.B1(n_819),
.B2(n_776),
.Y(n_874)
);

INVx6_ASAP7_75t_L g875 ( 
.A(n_821),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_783),
.A2(n_798),
.B1(n_771),
.B2(n_796),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_792),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_811),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_783),
.A2(n_795),
.B1(n_827),
.B2(n_807),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_816),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_797),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_SL g882 ( 
.A1(n_808),
.A2(n_581),
.B(n_694),
.Y(n_882)
);

CKINVDCx11_ASAP7_75t_R g883 ( 
.A(n_813),
.Y(n_883)
);

OAI22xp33_ASAP7_75t_L g884 ( 
.A1(n_825),
.A2(n_690),
.B1(n_694),
.B2(n_727),
.Y(n_884)
);

OAI22xp33_ASAP7_75t_L g885 ( 
.A1(n_779),
.A2(n_690),
.B1(n_581),
.B2(n_694),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_761),
.A2(n_690),
.B1(n_694),
.B2(n_620),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_760),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_760),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_789),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_813),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_760),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_845),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_832),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_834),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_835),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_861),
.Y(n_896)
);

INVx6_ASAP7_75t_L g897 ( 
.A(n_840),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_865),
.B(n_835),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_887),
.Y(n_899)
);

NOR2x1_ASAP7_75t_SL g900 ( 
.A(n_831),
.B(n_854),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_888),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_891),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_866),
.A2(n_852),
.B(n_864),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_860),
.Y(n_904)
);

AO21x2_ASAP7_75t_L g905 ( 
.A1(n_868),
.A2(n_866),
.B(n_872),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_837),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_839),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_830),
.B(n_838),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_831),
.B(n_842),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_856),
.B(n_829),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_885),
.A2(n_852),
.B1(n_859),
.B2(n_880),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_829),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_856),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_878),
.Y(n_914)
);

OA21x2_ASAP7_75t_L g915 ( 
.A1(n_879),
.A2(n_864),
.B(n_882),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_877),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_870),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_870),
.Y(n_918)
);

OAI21x1_ASAP7_75t_L g919 ( 
.A1(n_876),
.A2(n_881),
.B(n_859),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_873),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_847),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_SL g922 ( 
.A1(n_882),
.A2(n_886),
.B(n_846),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_869),
.B(n_858),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_875),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_875),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_848),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_840),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_851),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_851),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_874),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_841),
.B(n_855),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_862),
.B(n_874),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_889),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_844),
.B(n_843),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_886),
.B(n_884),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_884),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_836),
.A2(n_871),
.B(n_889),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_863),
.B(n_867),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_833),
.B(n_848),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_863),
.A2(n_867),
.B(n_850),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_883),
.B(n_890),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_849),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_857),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_845),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_913),
.B(n_914),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_898),
.B(n_895),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_892),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_941),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_892),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_909),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_893),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_921),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_945),
.Y(n_954)
);

AO31x2_ASAP7_75t_L g955 ( 
.A1(n_900),
.A2(n_903),
.A3(n_912),
.B(n_931),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_908),
.B(n_903),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_922),
.A2(n_911),
.B(n_936),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_909),
.B(n_894),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_945),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_910),
.B(n_919),
.Y(n_961)
);

AO21x2_ASAP7_75t_L g962 ( 
.A1(n_900),
.A2(n_905),
.B(n_931),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_910),
.B(n_919),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_939),
.B(n_924),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_901),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_905),
.A2(n_912),
.B(n_922),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_914),
.B(n_902),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_941),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_941),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_916),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_952),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_952),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_948),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_956),
.B(n_933),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_951),
.B(n_913),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_957),
.A2(n_933),
.B1(n_936),
.B2(n_930),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_958),
.B(n_916),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_967),
.B(n_906),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_953),
.B(n_907),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_899),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_960),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_947),
.B(n_907),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_970),
.B(n_899),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_947),
.B(n_908),
.Y(n_984)
);

BUFx6f_ASAP7_75t_SL g985 ( 
.A(n_949),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_960),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_948),
.A2(n_920),
.A3(n_929),
.B(n_930),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_952),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_965),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_950),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_967),
.B(n_915),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_946),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_961),
.B(n_915),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_971),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_971),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_949),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_980),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_981),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_981),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_972),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_986),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_972),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_988),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_988),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_991),
.B(n_955),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_977),
.B(n_969),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_986),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_991),
.B(n_955),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_980),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_1006),
.B(n_993),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_1006),
.B(n_993),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1002),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_998),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_998),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_996),
.B(n_968),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_997),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_997),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_999),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1010),
.B(n_975),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1010),
.B(n_975),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_996),
.B(n_977),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1013),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1014),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1015),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_996),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1022),
.B(n_996),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1020),
.B(n_976),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_1018),
.B(n_999),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_1030),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_SL g1032 ( 
.A(n_1026),
.B(n_942),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_1029),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1024),
.B(n_1017),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_SL g1035 ( 
.A(n_1026),
.B(n_942),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_1030),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_1030),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1036),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1031),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1031),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1035),
.A2(n_1027),
.B(n_1025),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1037),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1033),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_1032),
.B(n_943),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1036),
.B(n_1023),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1046),
.A2(n_1028),
.B1(n_1005),
.B2(n_1009),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1047),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1045),
.A2(n_1023),
.B(n_939),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1047),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_1011),
.Y(n_1052)
);

AOI221x1_ASAP7_75t_L g1053 ( 
.A1(n_1039),
.A2(n_1016),
.B1(n_943),
.B2(n_934),
.C(n_928),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_1038),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1040),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1054),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1054),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1052),
.B(n_1041),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1055),
.B(n_1043),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1049),
.B(n_1042),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

NOR2x1p5_ASAP7_75t_L g1062 ( 
.A(n_1050),
.B(n_896),
.Y(n_1062)
);

AOI221x1_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_1048),
.B1(n_1016),
.B2(n_1053),
.C(n_1013),
.Y(n_1063)
);

AOI21xp33_ASAP7_75t_L g1064 ( 
.A1(n_1057),
.A2(n_896),
.B(n_934),
.Y(n_1064)
);

AOI332xp33_ASAP7_75t_L g1065 ( 
.A1(n_1061),
.A2(n_944),
.A3(n_929),
.B1(n_1016),
.B2(n_928),
.B3(n_934),
.C1(n_924),
.C2(n_1001),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1060),
.B(n_968),
.Y(n_1066)
);

OAI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1060),
.A2(n_896),
.B1(n_897),
.B2(n_944),
.C(n_964),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1064),
.B(n_1059),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1066),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_1065),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_1063),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_1067),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1066),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_1058),
.C(n_1062),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_SL g1075 ( 
.A(n_1071),
.B(n_944),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_1071),
.B(n_940),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1069),
.Y(n_1077)
);

OA22x2_ASAP7_75t_L g1078 ( 
.A1(n_1070),
.A2(n_934),
.B1(n_928),
.B2(n_940),
.Y(n_1078)
);

AOI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1073),
.A2(n_928),
.B(n_969),
.C(n_968),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_R g1080 ( 
.A1(n_1077),
.A2(n_1072),
.B(n_1008),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1074),
.B(n_1011),
.Y(n_1081)
);

NOR2x1p5_ASAP7_75t_L g1082 ( 
.A(n_1076),
.B(n_1075),
.Y(n_1082)
);

XOR2x2_ASAP7_75t_L g1083 ( 
.A(n_1078),
.B(n_1012),
.Y(n_1083)
);

OAI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1079),
.A2(n_1012),
.B(n_1009),
.C(n_1005),
.Y(n_1084)
);

NAND4xp75_ASAP7_75t_L g1085 ( 
.A(n_1081),
.B(n_1021),
.C(n_1020),
.D(n_926),
.Y(n_1085)
);

AOI221x1_ASAP7_75t_L g1086 ( 
.A1(n_1080),
.A2(n_1082),
.B1(n_1083),
.B2(n_1084),
.C(n_1001),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_1081),
.B(n_969),
.C(n_968),
.Y(n_1087)
);

NAND5xp2_ASAP7_75t_L g1088 ( 
.A(n_1081),
.B(n_932),
.C(n_935),
.D(n_937),
.E(n_925),
.Y(n_1088)
);

OAI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1081),
.A2(n_968),
.B(n_969),
.C(n_926),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_1081),
.B(n_974),
.C(n_925),
.Y(n_1090)
);

OAI211xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1080),
.A2(n_897),
.B(n_937),
.C(n_920),
.Y(n_1091)
);

NAND4xp75_ASAP7_75t_L g1092 ( 
.A(n_1081),
.B(n_1021),
.C(n_932),
.D(n_935),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_1086),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_1088),
.B(n_987),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1091),
.B(n_938),
.C(n_904),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1087),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1085),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_1089),
.B(n_1008),
.Y(n_1098)
);

XNOR2x1_ASAP7_75t_L g1099 ( 
.A(n_1092),
.B(n_904),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_1090),
.B(n_938),
.C(n_904),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1086),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_SL g1102 ( 
.A(n_1097),
.B(n_897),
.C(n_979),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1093),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1101),
.B(n_938),
.C(n_897),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_1096),
.B(n_1099),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1095),
.B(n_1007),
.Y(n_1106)
);

AND4x1_ASAP7_75t_L g1107 ( 
.A(n_1100),
.B(n_897),
.C(n_985),
.D(n_983),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1094),
.B(n_987),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1098),
.B(n_969),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1093),
.Y(n_1110)
);

OR4x1_ASAP7_75t_L g1111 ( 
.A(n_1101),
.B(n_973),
.C(n_990),
.D(n_946),
.Y(n_1111)
);

AND3x4_ASAP7_75t_L g1112 ( 
.A(n_1096),
.B(n_918),
.C(n_927),
.Y(n_1112)
);

NOR2x1_ASAP7_75t_L g1113 ( 
.A(n_1101),
.B(n_1002),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1093),
.Y(n_1114)
);

XNOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_1105),
.B(n_918),
.Y(n_1115)
);

AOI222xp33_ASAP7_75t_L g1116 ( 
.A1(n_1103),
.A2(n_985),
.B1(n_995),
.B2(n_994),
.C1(n_1000),
.C2(n_1004),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1109),
.C(n_1104),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_1106),
.A2(n_1000),
.B(n_1004),
.C(n_995),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1111),
.Y(n_1119)
);

NAND5xp2_ASAP7_75t_L g1120 ( 
.A(n_1102),
.B(n_985),
.C(n_921),
.D(n_923),
.E(n_983),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1113),
.B(n_1107),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_L g1122 ( 
.A(n_1108),
.B(n_994),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1112),
.A2(n_1007),
.B1(n_1002),
.B2(n_1003),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1115),
.Y(n_1124)
);

AO22x1_ASAP7_75t_L g1125 ( 
.A1(n_1119),
.A2(n_1007),
.B1(n_1002),
.B2(n_1003),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1117),
.A2(n_1007),
.B1(n_1003),
.B2(n_927),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1121),
.A2(n_1003),
.B1(n_927),
.B2(n_918),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_982),
.B1(n_989),
.B2(n_917),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1120),
.A2(n_917),
.B1(n_963),
.B2(n_961),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1124),
.B(n_1122),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1127),
.Y(n_1131)
);

AOI311xp33_ASAP7_75t_L g1132 ( 
.A1(n_1129),
.A2(n_1116),
.A3(n_1118),
.B(n_923),
.C(n_950),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1130),
.B(n_1126),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1133),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_1128),
.B2(n_1125),
.Y(n_1135)
);

AOI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_1132),
.B(n_917),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1135),
.A2(n_966),
.B1(n_962),
.B2(n_963),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1136),
.A2(n_963),
.B1(n_961),
.B2(n_984),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1135),
.A2(n_963),
.B1(n_961),
.B2(n_978),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_987),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1139),
.B(n_987),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1137),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1142),
.B(n_978),
.Y(n_1143)
);

AO21x2_ASAP7_75t_L g1144 ( 
.A1(n_1141),
.A2(n_962),
.B(n_966),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1143),
.A2(n_1140),
.B1(n_959),
.B2(n_954),
.C(n_962),
.Y(n_1145)
);

AOI211xp5_ASAP7_75t_L g1146 ( 
.A1(n_1145),
.A2(n_1144),
.B(n_959),
.C(n_954),
.Y(n_1146)
);


endmodule