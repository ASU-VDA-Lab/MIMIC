module fake_netlist_6_2498_n_1547 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1547);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1547;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_859;
wire n_570;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_142),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_99),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_67),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_245),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_182),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_320),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_113),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_26),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_200),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_46),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_108),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_89),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_231),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_199),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_178),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_87),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_128),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_195),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_137),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_174),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_210),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_248),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_327),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_308),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_90),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_295),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_267),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_258),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_234),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_1),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_139),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_293),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_238),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_83),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_40),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_219),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_91),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_56),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_156),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_179),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_169),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_204),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_340),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_41),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_242),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_311),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_294),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_192),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_101),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_316),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_220),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_100),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_244),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_167),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_275),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_164),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_41),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_49),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_254),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_193),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_224),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_201),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_63),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_168),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_225),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_32),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_270),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_158),
.Y(n_426)
);

BUFx2_ASAP7_75t_SL g427 ( 
.A(n_33),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_166),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_286),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_344),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_290),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_12),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_150),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_230),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_312),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_229),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_235),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_343),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_226),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_190),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_21),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_326),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_313),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_132),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_227),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_57),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_196),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_301),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_39),
.B(n_102),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_66),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_7),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_46),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_151),
.Y(n_454)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_253),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_104),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_80),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_268),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_197),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_217),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_283),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_133),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_162),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_223),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_144),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_345),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_111),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_97),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_143),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_191),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_322),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_105),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_155),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_333),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_261),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_221),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_265),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_276),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_291),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_13),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_239),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_71),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_25),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_323),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_277),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_82),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_44),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_49),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_138),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_228),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_161),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_208),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_305),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_98),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_24),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_110),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_184),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_207),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_76),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_16),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_257),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_189),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_252),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_285),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_289),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_72),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_22),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_337),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_8),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_88),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_240),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_94),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_318),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_317),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_60),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_70),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_39),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_33),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_124),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_75),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_339),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_331),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_173),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_175),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_259),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_58),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_121),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_271),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_214),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_274),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_310),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_118),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_163),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_183),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_282),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_50),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_47),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_202),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_188),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_48),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_303),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_172),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_255),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_126),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_279),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_116),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_122),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_185),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_236),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_86),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_42),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_324),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_11),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_314),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_9),
.B(n_69),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_153),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_145),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_160),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_332),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_170),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_23),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_77),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_140),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_319),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_30),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_148),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_325),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_109),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_335),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_107),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_392),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_422),
.B(n_0),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_351),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_513),
.B(n_1),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_568),
.B(n_2),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_553),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_351),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_392),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_553),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_551),
.B(n_2),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_553),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_351),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_487),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_551),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_351),
.Y(n_587)
);

BUFx12f_ASAP7_75t_L g588 ( 
.A(n_480),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_513),
.B(n_3),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_400),
.A2(n_4),
.B(n_5),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_480),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g593 ( 
.A1(n_400),
.A2(n_6),
.B(n_7),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_354),
.Y(n_594)
);

BUFx6f_ASAP7_75t_SL g595 ( 
.A(n_394),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_401),
.B(n_9),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_389),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_561),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_424),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_477),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_356),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_389),
.Y(n_603)
);

BUFx8_ASAP7_75t_SL g604 ( 
.A(n_397),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_455),
.B(n_10),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_422),
.B(n_10),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_431),
.B(n_11),
.Y(n_607)
);

OAI22x1_ASAP7_75t_R g608 ( 
.A1(n_377),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_447),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_389),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_14),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_389),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_389),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_447),
.Y(n_615)
);

BUFx12f_ASAP7_75t_L g616 ( 
.A(n_379),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_522),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_386),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_431),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_522),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_564),
.B(n_15),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_415),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_389),
.Y(n_624)
);

BUFx12f_ASAP7_75t_L g625 ( 
.A(n_416),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_433),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_401),
.B(n_353),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_470),
.B(n_15),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_522),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_442),
.Y(n_630)
);

CKINVDCx6p67_ASAP7_75t_R g631 ( 
.A(n_470),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_452),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_507),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_348),
.A2(n_359),
.B(n_349),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_483),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_363),
.B(n_17),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_549),
.B(n_18),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_518),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_540),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_549),
.B(n_19),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_552),
.B(n_19),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_523),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_388),
.B(n_20),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_360),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_488),
.B(n_20),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_500),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_364),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_523),
.B(n_53),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_366),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_423),
.B(n_22),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_525),
.B(n_23),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_369),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_24),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_523),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_368),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_560),
.B(n_25),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_535),
.Y(n_660)
);

BUFx8_ASAP7_75t_SL g661 ( 
.A(n_376),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g662 ( 
.A(n_450),
.B(n_55),
.Y(n_662)
);

CKINVDCx6p67_ASAP7_75t_R g663 ( 
.A(n_427),
.Y(n_663)
);

BUFx8_ASAP7_75t_SL g664 ( 
.A(n_404),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_385),
.B(n_27),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_347),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_457),
.B(n_468),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_438),
.B(n_27),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_372),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_509),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_517),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_535),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_350),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_535),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_494),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_352),
.Y(n_677)
);

OA21x2_ASAP7_75t_L g678 ( 
.A1(n_381),
.A2(n_28),
.B(n_29),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_393),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_502),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_511),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_398),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_402),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_28),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_456),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_403),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_407),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_355),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_408),
.B(n_59),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_357),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_380),
.B(n_29),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_536),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_537),
.Y(n_694)
);

BUFx12f_ASAP7_75t_L g695 ( 
.A(n_565),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_532),
.B(n_30),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_358),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_441),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_473),
.B(n_34),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_409),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_410),
.B(n_35),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_414),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_361),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_421),
.B(n_35),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_362),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_432),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_436),
.Y(n_707)
);

OA21x2_ASAP7_75t_L g708 ( 
.A1(n_445),
.A2(n_36),
.B(n_37),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_471),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_449),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_365),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_451),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_454),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_367),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_462),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_478),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_515),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_467),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_469),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_474),
.B(n_43),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_475),
.B(n_43),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_476),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_485),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_490),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_491),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_573),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_576),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_661),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_664),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_604),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_666),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_674),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_658),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_677),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_580),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_689),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_703),
.B(n_493),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_709),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_691),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_685),
.B(n_496),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_602),
.B(n_370),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_616),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_573),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_578),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_625),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_647),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_577),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_671),
.Y(n_750)
);

BUFx8_ASAP7_75t_L g751 ( 
.A(n_595),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_580),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_694),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_595),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_695),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_685),
.B(n_505),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_631),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_618),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_703),
.B(n_506),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_663),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_R g762 ( 
.A(n_670),
.B(n_527),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_697),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_582),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_714),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_571),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_584),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_579),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_705),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_705),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_670),
.B(n_371),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_705),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_711),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_711),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_711),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_588),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_592),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_577),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_635),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_577),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_648),
.B(n_373),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_583),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_583),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_632),
.B(n_374),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_679),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_620),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_615),
.B(n_44),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_683),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_609),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_583),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_693),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_587),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_686),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_687),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_685),
.B(n_531),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_706),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_692),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_725),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_581),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_575),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_615),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_688),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_688),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_715),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_651),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_611),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_654),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_682),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_605),
.B(n_375),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_688),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_R g814 ( 
.A(n_690),
.B(n_533),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_680),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_642),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_707),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_680),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_680),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_681),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_594),
.B(n_378),
.Y(n_821)
);

INVx8_ASAP7_75t_L g822 ( 
.A(n_690),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_681),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_681),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_587),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_759),
.B(n_622),
.C(n_767),
.Y(n_826)
);

INVxp33_ASAP7_75t_L g827 ( 
.A(n_799),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_799),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_817),
.B(n_653),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_808),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_812),
.B(n_676),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_821),
.B(n_702),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_773),
.B(n_676),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_803),
.B(n_699),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_759),
.B(n_590),
.C(n_574),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_810),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_767),
.B(n_667),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_760),
.B(n_676),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_763),
.B(n_765),
.Y(n_839)
);

BUFx5_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_802),
.B(n_717),
.C(n_698),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_786),
.B(n_643),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_811),
.Y(n_843)
);

NOR3xp33_ASAP7_75t_L g844 ( 
.A(n_781),
.B(n_696),
.C(n_668),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_815),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_793),
.B(n_627),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_783),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_726),
.B(n_643),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_744),
.B(n_672),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_742),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_746),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_762),
.B(n_656),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_820),
.B(n_656),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_824),
.B(n_667),
.Y(n_856)
);

AO221x1_ASAP7_75t_L g857 ( 
.A1(n_766),
.A2(n_543),
.B1(n_544),
.B2(n_541),
.C(n_534),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_741),
.B(n_672),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_816),
.B(n_636),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_745),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_782),
.B(n_659),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_770),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_788),
.B(n_572),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_792),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_789),
.Y(n_865)
);

NAND3xp33_ASAP7_75t_L g866 ( 
.A(n_738),
.B(n_596),
.C(n_641),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_780),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_757),
.A2(n_665),
.B(n_701),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_825),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_819),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_823),
.B(n_730),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_736),
.B(n_634),
.Y(n_872)
);

NAND2xp33_ASAP7_75t_L g873 ( 
.A(n_814),
.B(n_690),
.Y(n_873)
);

INVxp33_ASAP7_75t_L g874 ( 
.A(n_787),
.Y(n_874)
);

BUFx6f_ASAP7_75t_SL g875 ( 
.A(n_755),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_752),
.B(n_634),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_809),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_791),
.B(n_572),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_754),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_732),
.B(n_606),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_797),
.B(n_724),
.Y(n_881)
);

AOI221xp5_ASAP7_75t_L g882 ( 
.A1(n_801),
.A2(n_586),
.B1(n_684),
.B2(n_646),
.C(n_652),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_822),
.A2(n_684),
.B1(n_720),
.B2(n_704),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_764),
.B(n_704),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_790),
.B(n_644),
.C(n_607),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_768),
.B(n_720),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_769),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_733),
.B(n_735),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_761),
.B(n_650),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_780),
.B(n_721),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_737),
.B(n_606),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_780),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_804),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_780),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_795),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_784),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_796),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_740),
.A2(n_690),
.B1(n_637),
.B2(n_640),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_771),
.B(n_650),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_784),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_798),
.B(n_724),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_806),
.B(n_637),
.C(n_628),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_784),
.B(n_640),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_805),
.B(n_645),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_784),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_785),
.B(n_657),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_813),
.B(n_645),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_785),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_785),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_785),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_758),
.B(n_382),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_755),
.B(n_383),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_794),
.B(n_673),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_822),
.A2(n_669),
.B(n_712),
.C(n_649),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_728),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_807),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_863),
.B(n_830),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_837),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_847),
.B(n_772),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_867),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_867),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_863),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_867),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_836),
.B(n_843),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_915),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_895),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_851),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_903),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_897),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_890),
.Y(n_930)
);

AND2x6_ASAP7_75t_SL g931 ( 
.A(n_839),
.B(n_608),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_916),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_856),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_888),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_871),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_L g936 ( 
.A(n_829),
.B(n_882),
.C(n_826),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_877),
.B(n_626),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_883),
.B(n_822),
.Y(n_938)
);

NOR2x1p5_ASAP7_75t_L g939 ( 
.A(n_835),
.B(n_779),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_875),
.B(n_729),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_905),
.Y(n_941)
);

CKINVDCx16_ASAP7_75t_R g942 ( 
.A(n_860),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_832),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_827),
.B(n_800),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_872),
.A2(n_708),
.B(n_678),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_846),
.B(n_774),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_850),
.A2(n_662),
.B1(n_387),
.B2(n_390),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_877),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_879),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_859),
.B(n_775),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_877),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_904),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_842),
.B(n_776),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_853),
.B(n_777),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_887),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_844),
.B(n_778),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_868),
.B(n_558),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_841),
.B(n_716),
.C(n_669),
.Y(n_959)
);

NOR3xp33_ASAP7_75t_L g960 ( 
.A(n_834),
.B(n_731),
.C(n_743),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_876),
.A2(n_708),
.B1(n_678),
.B2(n_593),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_828),
.B(n_747),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_862),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_861),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_905),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_902),
.A2(n_391),
.B1(n_395),
.B2(n_384),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_865),
.B(n_734),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_905),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_907),
.A2(n_650),
.B1(n_563),
.B2(n_566),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_866),
.B(n_562),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_864),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_SL g972 ( 
.A(n_880),
.B(n_396),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_869),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_900),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_874),
.B(n_748),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_891),
.B(n_750),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_906),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_845),
.B(n_633),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_857),
.A2(n_593),
.B1(n_591),
.B2(n_650),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_833),
.B(n_567),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_898),
.A2(n_570),
.B(n_712),
.C(n_649),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_840),
.B(n_591),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_889),
.B(n_753),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_840),
.B(n_884),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_886),
.A2(n_603),
.B1(n_610),
.B2(n_597),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_913),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_885),
.A2(n_612),
.B1(n_624),
.B2(n_614),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_862),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_855),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_854),
.B(n_756),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_900),
.A2(n_894),
.B(n_892),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_878),
.B(n_739),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_831),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_870),
.B(n_638),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_893),
.B(n_639),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_848),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_849),
.Y(n_997)
);

BUFx12f_ASAP7_75t_L g998 ( 
.A(n_875),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_896),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_911),
.B(n_912),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_840),
.A2(n_700),
.B1(n_718),
.B2(n_710),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_908),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_909),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_838),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_910),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_914),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_858),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_840),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_901),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_840),
.B(n_399),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_873),
.A2(n_899),
.B1(n_700),
.B2(n_718),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_881),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_L g1013 ( 
.A(n_901),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_881),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_950),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_942),
.A2(n_630),
.B1(n_599),
.B2(n_406),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_982),
.A2(n_858),
.B(n_675),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_922),
.B(n_599),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_956),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_964),
.B(n_405),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_928),
.B(n_411),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_998),
.B(n_630),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_978),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_917),
.B(n_918),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_917),
.B(n_585),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_984),
.A2(n_794),
.B(n_589),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_934),
.B(n_412),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1008),
.A2(n_794),
.B(n_589),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_920),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_920),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_943),
.B(n_585),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_959),
.B(n_417),
.C(n_413),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_936),
.A2(n_710),
.B1(n_718),
.B2(n_700),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_944),
.B(n_598),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_935),
.B(n_418),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_953),
.B(n_419),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_975),
.B(n_598),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_920),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_951),
.B(n_420),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_945),
.A2(n_426),
.B(n_425),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_937),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1008),
.A2(n_794),
.B(n_589),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_925),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_930),
.B(n_428),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_991),
.A2(n_62),
.B(n_61),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_958),
.A2(n_600),
.B(n_587),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_980),
.A2(n_986),
.B(n_970),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_961),
.A2(n_601),
.B(n_600),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_996),
.B(n_429),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_938),
.A2(n_434),
.B1(n_435),
.B2(n_430),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1010),
.A2(n_439),
.B(n_437),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_1006),
.A2(n_710),
.B1(n_723),
.B2(n_722),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1007),
.A2(n_601),
.B(n_600),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_977),
.A2(n_613),
.B(n_601),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_974),
.A2(n_65),
.B(n_64),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_981),
.A2(n_524),
.B(n_443),
.C(n_444),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_923),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_946),
.B(n_440),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_997),
.B(n_446),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_937),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_933),
.B(n_448),
.Y(n_1061)
);

INVx3_ASAP7_75t_SL g1062 ( 
.A(n_988),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_954),
.B(n_1009),
.Y(n_1063)
);

NAND2x1p5_ASAP7_75t_L g1064 ( 
.A(n_921),
.B(n_613),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_924),
.B(n_458),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_1003),
.A2(n_73),
.B(n_68),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_924),
.B(n_459),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_921),
.A2(n_617),
.B(n_613),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_979),
.A2(n_1003),
.B(n_1011),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_993),
.A2(n_530),
.B(n_461),
.C(n_464),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_SL g1071 ( 
.A1(n_1014),
.A2(n_719),
.B(n_722),
.C(n_723),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_974),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_R g1073 ( 
.A(n_1004),
.B(n_751),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_932),
.B(n_460),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_995),
.B(n_465),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_R g1076 ( 
.A(n_972),
.B(n_751),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_921),
.A2(n_619),
.B(n_617),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_941),
.A2(n_619),
.B(n_617),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_967),
.B(n_466),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_962),
.B(n_719),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_941),
.A2(n_968),
.B(n_965),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1006),
.A2(n_528),
.B1(n_479),
.B2(n_481),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_941),
.A2(n_621),
.B(n_619),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_994),
.Y(n_1084)
);

INVx3_ASAP7_75t_SL g1085 ( 
.A(n_952),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1002),
.A2(n_78),
.B(n_74),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_926),
.A2(n_521),
.B(n_482),
.C(n_484),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_929),
.B(n_79),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_948),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_965),
.A2(n_629),
.B(n_621),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_1000),
.B(n_472),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1014),
.A2(n_542),
.B1(n_489),
.B2(n_492),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1006),
.A2(n_722),
.B1(n_719),
.B2(n_723),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_994),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_973),
.B(n_486),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1085),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1017),
.A2(n_1005),
.B(n_949),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_1043),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1030),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1048),
.A2(n_987),
.B(n_985),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1037),
.B(n_992),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1045),
.A2(n_949),
.B(n_927),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_1040),
.A2(n_955),
.B(n_947),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1015),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1019),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1086),
.A2(n_927),
.B(n_989),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1025),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1025),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1062),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_1047),
.A2(n_971),
.B(n_919),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_1051),
.A2(n_983),
.B(n_957),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1034),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1026),
.A2(n_966),
.B(n_990),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1063),
.B(n_999),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1031),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_1055),
.A2(n_976),
.B(n_960),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1030),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1028),
.A2(n_1001),
.B(n_939),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_1094),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1042),
.A2(n_923),
.B(n_965),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1056),
.A2(n_969),
.B(n_1012),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1072),
.Y(n_1122)
);

CKINVDCx11_ASAP7_75t_R g1123 ( 
.A(n_1022),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1081),
.A2(n_923),
.B(n_968),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1035),
.A2(n_1012),
.B(n_968),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_1039),
.A2(n_1013),
.B(n_498),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1030),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1057),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1057),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1018),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1071),
.A2(n_499),
.B(n_497),
.Y(n_1131)
);

NAND2x1p5_ASAP7_75t_L g1132 ( 
.A(n_1029),
.B(n_963),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_1057),
.Y(n_1133)
);

BUFx2_ASAP7_75t_SL g1134 ( 
.A(n_1089),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1018),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1029),
.B(n_621),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1058),
.B(n_501),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1022),
.B(n_940),
.Y(n_1138)
);

AO21x2_ASAP7_75t_L g1139 ( 
.A1(n_1091),
.A2(n_504),
.B(n_503),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_1038),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1046),
.A2(n_84),
.B(n_81),
.Y(n_1141)
);

AOI22x1_ASAP7_75t_L g1142 ( 
.A1(n_1088),
.A2(n_547),
.B1(n_510),
.B2(n_512),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1069),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1060),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1084),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1023),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1073),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1038),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1024),
.Y(n_1149)
);

BUFx5_ASAP7_75t_L g1150 ( 
.A(n_1024),
.Y(n_1150)
);

INVxp67_ASAP7_75t_SL g1151 ( 
.A(n_1069),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1095),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

INVx5_ASAP7_75t_L g1154 ( 
.A(n_1066),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1080),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1032),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_1065),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1061),
.B(n_629),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1074),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1079),
.B(n_508),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1027),
.B(n_514),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1064),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1054),
.A2(n_92),
.B(n_85),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1076),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1049),
.A2(n_520),
.B(n_516),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_SL g1166 ( 
.A1(n_1101),
.A2(n_1016),
.B1(n_1036),
.B2(n_1067),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1143),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1159),
.B(n_1033),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1104),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1115),
.B(n_1075),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1143),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1109),
.A2(n_1020),
.B1(n_931),
.B2(n_1059),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1119),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1122),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1122),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1156),
.A2(n_1157),
.B1(n_1135),
.B2(n_1130),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1105),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1097),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1148),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1151),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1148),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1134),
.Y(n_1182)
);

AOI222xp33_ASAP7_75t_L g1183 ( 
.A1(n_1112),
.A2(n_1021),
.B1(n_1044),
.B2(n_1082),
.C1(n_1050),
.C2(n_526),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1157),
.A2(n_1092),
.B1(n_1093),
.B2(n_1052),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1152),
.B(n_1070),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1151),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1145),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1106),
.A2(n_1053),
.B(n_1068),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1102),
.A2(n_1078),
.B(n_1077),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1114),
.B(n_529),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1131),
.A2(n_1103),
.B(n_1100),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1161),
.A2(n_556),
.B1(n_538),
.B2(n_545),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1146),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1160),
.A2(n_1137),
.B1(n_1114),
.B2(n_1155),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1150),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1153),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1131),
.A2(n_1090),
.B(n_1083),
.Y(n_1197)
);

OA21x2_ASAP7_75t_L g1198 ( 
.A1(n_1100),
.A2(n_554),
.B(n_546),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1150),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1107),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1108),
.A2(n_557),
.B1(n_548),
.B2(n_550),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1160),
.A2(n_1087),
.B1(n_569),
.B2(n_559),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1150),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1155),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1096),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1109),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1137),
.A2(n_660),
.B1(n_655),
.B2(n_629),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1129),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1140),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1110),
.A2(n_211),
.B(n_346),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1141),
.A2(n_660),
.B(n_655),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1150),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1144),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1149),
.A2(n_660),
.B1(n_655),
.B2(n_48),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1138),
.A2(n_1142),
.B1(n_1098),
.B2(n_1111),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1163),
.A2(n_212),
.B(n_338),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1150),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1110),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1150),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1128),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1096),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1120),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1136),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1138),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1118),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1136),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1149),
.A2(n_51),
.B1(n_52),
.B2(n_93),
.Y(n_1227)
);

BUFx2_ASAP7_75t_R g1228 ( 
.A(n_1144),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1128),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1125),
.A2(n_95),
.B(n_96),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1124),
.A2(n_103),
.B(n_106),
.Y(n_1231)
);

NAND2x1p5_ASAP7_75t_L g1232 ( 
.A(n_1154),
.B(n_112),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1133),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1147),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1194),
.A2(n_1154),
.A3(n_1140),
.B1(n_1126),
.B2(n_1165),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1190),
.B(n_1126),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1205),
.B(n_1098),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1166),
.B(n_1147),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1174),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1170),
.B(n_1138),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1174),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1185),
.A2(n_1139),
.B1(n_1165),
.B2(n_1116),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1234),
.A2(n_1192),
.B1(n_1182),
.B2(n_1204),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1206),
.B(n_1123),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1175),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_R g1246 ( 
.A(n_1213),
.B(n_1123),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1175),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1190),
.B(n_1132),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_R g1249 ( 
.A(n_1213),
.B(n_1164),
.Y(n_1249)
);

AO32x2_ASAP7_75t_L g1250 ( 
.A1(n_1214),
.A2(n_1154),
.A3(n_1139),
.B1(n_1116),
.B2(n_1121),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1173),
.B(n_1158),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1185),
.A2(n_1113),
.B1(n_1164),
.B2(n_1158),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1196),
.B(n_1113),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_R g1254 ( 
.A(n_1198),
.B(n_119),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1168),
.A2(n_1154),
.B(n_1162),
.C(n_1133),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_1099),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1206),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_R g1258 ( 
.A(n_1205),
.B(n_1099),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1228),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1183),
.B(n_1121),
.C(n_1133),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1187),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1180),
.A2(n_1133),
.B(n_1127),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1221),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1177),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1208),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1200),
.B(n_1193),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1233),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1209),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1172),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1189),
.A2(n_1127),
.B(n_1117),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1215),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1176),
.B(n_1099),
.Y(n_1273)
);

INVxp33_ASAP7_75t_SL g1274 ( 
.A(n_1224),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_R g1275 ( 
.A(n_1209),
.B(n_1117),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1186),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1167),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1167),
.Y(n_1278)
);

OR2x6_ASAP7_75t_L g1279 ( 
.A(n_1232),
.B(n_1117),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_R g1280 ( 
.A(n_1198),
.B(n_1209),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1184),
.A2(n_1162),
.B1(n_1127),
.B2(n_1117),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1179),
.B(n_1127),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1201),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1220),
.B(n_127),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1186),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1180),
.B(n_129),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1171),
.Y(n_1287)
);

OAI222xp33_ASAP7_75t_L g1288 ( 
.A1(n_1227),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.C1(n_135),
.C2(n_136),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1171),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_R g1290 ( 
.A(n_1179),
.B(n_141),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1229),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_R g1292 ( 
.A(n_1181),
.B(n_1231),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1181),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1171),
.B(n_146),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1181),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1231),
.B(n_147),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1202),
.A2(n_149),
.B(n_152),
.C(n_154),
.Y(n_1297)
);

CKINVDCx16_ASAP7_75t_R g1298 ( 
.A(n_1207),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1195),
.B(n_1199),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1195),
.B(n_1199),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1203),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1276),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1285),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1253),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1236),
.B(n_1191),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1240),
.B(n_1203),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1299),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1256),
.B(n_1191),
.Y(n_1308)
);

OAI221xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1238),
.A2(n_1198),
.B1(n_1225),
.B2(n_1212),
.C(n_1217),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1300),
.B(n_1218),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1266),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1248),
.B(n_1212),
.Y(n_1312)
);

OR2x2_ASAP7_75t_SL g1313 ( 
.A(n_1261),
.B(n_1225),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1262),
.B(n_1191),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1260),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1274),
.A2(n_1217),
.B1(n_1219),
.B2(n_1232),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1265),
.B(n_1219),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1258),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1277),
.B(n_1210),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1278),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1267),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1264),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1267),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1279),
.B(n_1223),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1301),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1257),
.B(n_1232),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_SL g1327 ( 
.A(n_1298),
.B(n_1223),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1251),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1255),
.A2(n_1178),
.A3(n_1222),
.B(n_1226),
.Y(n_1329)
);

NOR2x1_ASAP7_75t_L g1330 ( 
.A(n_1237),
.B(n_1210),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1239),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1271),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1241),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1287),
.B(n_1289),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1243),
.B(n_1226),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1235),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1235),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1247),
.B(n_1210),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1235),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1242),
.B(n_1178),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1291),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1273),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1268),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1295),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1250),
.B(n_1222),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1293),
.B(n_1197),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1250),
.B(n_1230),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1272),
.B(n_157),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1250),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1269),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1279),
.B(n_1230),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1295),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1286),
.Y(n_1354)
);

NAND2x1_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_1211),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1252),
.B(n_1216),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1294),
.B(n_1211),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1269),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1269),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1284),
.B(n_1292),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1281),
.B(n_1211),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1237),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1282),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1259),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1280),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1306),
.B(n_1270),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1366),
.B(n_1297),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1305),
.B(n_1244),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1303),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1303),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1314),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1304),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1308),
.B(n_1296),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1308),
.B(n_1197),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1314),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1310),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1310),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1312),
.B(n_1290),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1307),
.B(n_1283),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1343),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1341),
.B(n_1188),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1328),
.B(n_1246),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1362),
.B(n_1188),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1364),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1335),
.B(n_1288),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1307),
.B(n_159),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1320),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1315),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1321),
.B(n_165),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1311),
.B(n_171),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1320),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1354),
.B(n_1322),
.Y(n_1394)
);

AOI211xp5_ASAP7_75t_L g1395 ( 
.A1(n_1349),
.A2(n_1254),
.B(n_1249),
.C(n_177),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1323),
.B(n_176),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1331),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1331),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1346),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1317),
.B(n_180),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1333),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1346),
.B(n_181),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1362),
.B(n_186),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1319),
.B(n_187),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1319),
.B(n_194),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1333),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1337),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1317),
.B(n_198),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1337),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1339),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1339),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1342),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1348),
.B(n_1336),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1325),
.B(n_203),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1361),
.A2(n_1189),
.B(n_206),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1367),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1378),
.B(n_1336),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1379),
.B(n_1338),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1374),
.B(n_1356),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1386),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1382),
.B(n_1360),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1370),
.B(n_1360),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1367),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1372),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1384),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1368),
.B(n_1380),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1373),
.B(n_1356),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1375),
.B(n_1325),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1326),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1412),
.B(n_1327),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1394),
.B(n_1390),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1373),
.B(n_1338),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1387),
.B(n_1340),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1410),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1413),
.B(n_1344),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1377),
.B(n_1364),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1377),
.B(n_1313),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1411),
.B(n_1313),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1397),
.B(n_1347),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1369),
.B(n_1330),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1371),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1386),
.B(n_1365),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1398),
.B(n_1334),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1411),
.B(n_1353),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1399),
.B(n_1357),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1402),
.B(n_1324),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1416),
.Y(n_1447)
);

INVxp33_ASAP7_75t_L g1448 ( 
.A(n_1442),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1437),
.Y(n_1449)
);

CKINVDCx14_ASAP7_75t_R g1450 ( 
.A(n_1420),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1428),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1425),
.B(n_1376),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1433),
.A2(n_1395),
.B1(n_1425),
.B2(n_1369),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1423),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1424),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1445),
.Y(n_1456)
);

NAND2x2_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1318),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1440),
.B(n_1369),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1438),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1436),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1441),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1435),
.B(n_1376),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1420),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1426),
.A2(n_1316),
.B1(n_1309),
.B2(n_1422),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1429),
.Y(n_1465)
);

XNOR2x2_ASAP7_75t_L g1466 ( 
.A(n_1421),
.B(n_1402),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1461),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1447),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1454),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1455),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1464),
.A2(n_1404),
.B1(n_1405),
.B2(n_1446),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1464),
.A2(n_1404),
.B1(n_1405),
.B2(n_1414),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1449),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1449),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1456),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1456),
.Y(n_1477)
);

OAI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1439),
.B(n_1419),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1450),
.A2(n_1381),
.B(n_1392),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1457),
.A2(n_1318),
.B1(n_1363),
.B2(n_1417),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1457),
.A2(n_1427),
.B1(n_1418),
.B2(n_1432),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1450),
.A2(n_1465),
.B1(n_1448),
.B2(n_1458),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1463),
.A2(n_1385),
.B1(n_1352),
.B2(n_1383),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1472),
.A2(n_1466),
.B1(n_1458),
.B2(n_1451),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1471),
.Y(n_1485)
);

AOI21xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1482),
.A2(n_1458),
.B(n_1460),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1479),
.B(n_1452),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1467),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1478),
.B(n_1462),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1480),
.A2(n_1350),
.B1(n_1396),
.B2(n_1400),
.Y(n_1490)
);

AOI32xp33_ASAP7_75t_L g1491 ( 
.A1(n_1481),
.A2(n_1477),
.A3(n_1475),
.B1(n_1476),
.B2(n_1469),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1483),
.A2(n_1350),
.B1(n_1408),
.B2(n_1403),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1473),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1468),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1474),
.A2(n_1443),
.B(n_1388),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1470),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1485),
.B(n_1434),
.Y(n_1497)
);

NAND2xp33_ASAP7_75t_L g1498 ( 
.A(n_1491),
.B(n_1444),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1493),
.B(n_1358),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1484),
.A2(n_1348),
.B1(n_1383),
.B2(n_1391),
.C(n_1407),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1489),
.B(n_1358),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1495),
.B(n_1359),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_1487),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_SL g1504 ( 
.A(n_1486),
.B(n_1409),
.C(n_1401),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1490),
.B(n_1345),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1499),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1504),
.B(n_1498),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1501),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1503),
.A2(n_1492),
.B1(n_1494),
.B2(n_1496),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1497),
.B(n_1488),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1502),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1505),
.B(n_1500),
.Y(n_1512)
);

OAI211xp5_ASAP7_75t_L g1513 ( 
.A1(n_1507),
.A2(n_1512),
.B(n_1509),
.C(n_1510),
.Y(n_1513)
);

AOI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1511),
.A2(n_1406),
.B1(n_1393),
.B2(n_1389),
.C(n_1324),
.Y(n_1514)
);

AOI222xp33_ASAP7_75t_L g1515 ( 
.A1(n_1511),
.A2(n_1406),
.B1(n_1393),
.B2(n_1389),
.C1(n_1332),
.C2(n_1415),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1506),
.B(n_1355),
.C(n_1332),
.Y(n_1516)
);

NAND4xp25_ASAP7_75t_SL g1517 ( 
.A(n_1508),
.B(n_1357),
.C(n_1415),
.D(n_1351),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1507),
.A2(n_1332),
.B1(n_1355),
.B2(n_1329),
.Y(n_1518)
);

NAND4xp25_ASAP7_75t_L g1519 ( 
.A(n_1507),
.B(n_205),
.C(n_209),
.D(n_213),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1518),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_L g1521 ( 
.A1(n_1513),
.A2(n_215),
.B(n_216),
.C(n_218),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1519),
.A2(n_1329),
.B1(n_232),
.B2(n_237),
.Y(n_1522)
);

NOR2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1517),
.B(n_222),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1514),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1516),
.Y(n_1525)
);

AND3x4_ASAP7_75t_L g1526 ( 
.A(n_1520),
.B(n_1515),
.C(n_1329),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1524),
.Y(n_1527)
);

NOR2x1_ASAP7_75t_L g1528 ( 
.A(n_1521),
.B(n_241),
.Y(n_1528)
);

AOI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1527),
.A2(n_1525),
.B(n_1522),
.C(n_1523),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1528),
.Y(n_1530)
);

CKINVDCx16_ASAP7_75t_R g1531 ( 
.A(n_1526),
.Y(n_1531)
);

XOR2xp5_ASAP7_75t_L g1532 ( 
.A(n_1530),
.B(n_243),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1531),
.A2(n_1329),
.B1(n_247),
.B2(n_249),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1533),
.A2(n_1529),
.B1(n_250),
.B2(n_251),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1532),
.A2(n_246),
.B1(n_256),
.B2(n_260),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1532),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1535),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1534),
.A2(n_266),
.B1(n_269),
.B2(n_272),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1536),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1537),
.A2(n_273),
.B1(n_278),
.B2(n_280),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1539),
.Y(n_1541)
);

NAND3xp33_ASAP7_75t_L g1542 ( 
.A(n_1541),
.B(n_1538),
.C(n_281),
.Y(n_1542)
);

AOI21xp33_ASAP7_75t_L g1543 ( 
.A1(n_1540),
.A2(n_284),
.B(n_287),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1542),
.A2(n_292),
.B1(n_298),
.B2(n_299),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1543),
.A2(n_300),
.B1(n_302),
.B2(n_304),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1545),
.A2(n_342),
.B1(n_328),
.B2(n_329),
.C(n_330),
.Y(n_1546)
);

AOI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1546),
.A2(n_1544),
.B(n_334),
.C(n_336),
.Y(n_1547)
);


endmodule