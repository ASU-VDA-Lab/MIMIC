module fake_jpeg_5541_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_54),
.Y(n_79)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_57),
.Y(n_94)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_26),
.B1(n_34),
.B2(n_33),
.Y(n_99)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_78),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_44),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_0),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_20),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_49),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_43),
.B1(n_42),
.B2(n_48),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_98),
.B1(n_99),
.B2(n_28),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_39),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_52),
.CI(n_49),
.CON(n_104),
.SN(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_92),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_30),
.B1(n_31),
.B2(n_47),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_114),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_107),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_34),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_111),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_115),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_113),
.B1(n_131),
.B2(n_28),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_31),
.B1(n_73),
.B2(n_68),
.Y(n_113)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_39),
.A3(n_36),
.B1(n_67),
.B2(n_53),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_118),
.B1(n_121),
.B2(n_85),
.Y(n_143)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_17),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_53),
.B1(n_66),
.B2(n_64),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_27),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_130),
.Y(n_141)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_39),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_76),
.C(n_29),
.Y(n_139)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_95),
.B(n_0),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_134),
.Y(n_173)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_153),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_22),
.C(n_9),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_120),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_20),
.B1(n_22),
.B2(n_29),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_90),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_70),
.B1(n_93),
.B2(n_76),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_123),
.B1(n_85),
.B2(n_118),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_77),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_92),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_97),
.B1(n_93),
.B2(n_51),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_104),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_184),
.C(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_165),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_124),
.C(n_117),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_156),
.B(n_157),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_163),
.B1(n_157),
.B2(n_144),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_19),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_126),
.B1(n_105),
.B2(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_153),
.B(n_147),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_175),
.B(n_19),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_90),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_180),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_106),
.B(n_112),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_95),
.B1(n_81),
.B2(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_132),
.B1(n_81),
.B2(n_145),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx10_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_91),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_203),
.B(n_184),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_212),
.B(n_21),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_175),
.C(n_170),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_190),
.B(n_192),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_145),
.B1(n_154),
.B2(n_134),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_17),
.Y(n_238)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_207),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_97),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_178),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_171),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_17),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_127),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_213),
.B(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_233),
.B1(n_211),
.B2(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_163),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_180),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_161),
.B(n_167),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_238),
.C(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_177),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_182),
.B(n_178),
.Y(n_225)
);

XNOR2x2_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_237),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_195),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_236),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_19),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_188),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_200),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_240),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_245),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_185),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_254),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_193),
.C(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_187),
.C(n_196),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_187),
.B1(n_207),
.B2(n_103),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_257),
.B1(n_213),
.B2(n_218),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_137),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_17),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_103),
.B1(n_137),
.B2(n_21),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_97),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_214),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_19),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_234),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_216),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_264),
.B(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_215),
.B(n_223),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_8),
.B(n_16),
.Y(n_290)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_216),
.B1(n_224),
.B2(n_220),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_279),
.B1(n_251),
.B2(n_247),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_249),
.C(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_220),
.B1(n_230),
.B2(n_222),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_241),
.A2(n_219),
.B1(n_23),
.B2(n_47),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_247),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_290),
.B(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

A2O1A1O1Ixp25_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_239),
.B(n_246),
.C(n_256),
.D(n_219),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_268),
.B(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_23),
.C(n_1),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.C(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_23),
.C(n_1),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_300),
.B(n_301),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_279),
.B1(n_273),
.B2(n_274),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_310),
.B1(n_292),
.B2(n_293),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_265),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_0),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_305),
.B(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_1),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_9),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_300),
.B1(n_8),
.B2(n_11),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_23),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_298),
.C(n_308),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_317),
.B(n_319),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_297),
.A2(n_284),
.B1(n_296),
.B2(n_291),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_313),
.B(n_318),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_294),
.Y(n_314)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_11),
.B(n_15),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_283),
.C(n_289),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_1),
.C(n_2),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_324),
.A2(n_320),
.B(n_311),
.C(n_317),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_7),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_7),
.Y(n_328)
);

OAI21x1_ASAP7_75t_SL g329 ( 
.A1(n_314),
.A2(n_7),
.B(n_13),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_334),
.B(n_322),
.C(n_12),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_4),
.B(n_6),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_330),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.A3(n_332),
.B1(n_4),
.B2(n_6),
.C1(n_12),
.C2(n_13),
.Y(n_339)
);

OAI21x1_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_13),
.B(n_16),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_16),
.C(n_2),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_3),
.B(n_328),
.Y(n_342)
);


endmodule