module fake_ariane_1344_n_167 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_167);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_167;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_94;
wire n_101;
wire n_48;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_121;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_0),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_2),
.C(n_3),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_3),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_4),
.C(n_5),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_32),
.B(n_6),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_47),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_47),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_54),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_50),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_62),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_R g91 ( 
.A(n_85),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_81),
.B(n_76),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_66),
.B(n_61),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_73),
.B(n_72),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_56),
.B(n_66),
.C(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_68),
.B(n_64),
.Y(n_100)
);

OA21x2_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_88),
.B(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_85),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_60),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_86),
.C(n_57),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_83),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_95),
.B(n_104),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_108),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_109),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_41),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_107),
.C(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_107),
.B1(n_110),
.B2(n_63),
.Y(n_134)
);

NAND4xp75_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_134),
.C(n_133),
.D(n_129),
.Y(n_135)
);

AOI211xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_57),
.B(n_63),
.C(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_118),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_122),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_92),
.B1(n_48),
.B2(n_111),
.Y(n_139)
);

AOI311xp33_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_45),
.A3(n_49),
.B(n_73),
.C(n_7),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_122),
.Y(n_141)
);

AOI222xp33_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_64),
.B1(n_83),
.B2(n_119),
.C1(n_126),
.C2(n_72),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_111),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_72),
.C(n_66),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_59),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

AOI211xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_66),
.B(n_103),
.C(n_59),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_10),
.C(n_11),
.Y(n_152)
);

NAND4xp75_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_96),
.C(n_103),
.D(n_101),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_10),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND4xp75_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_101),
.C(n_96),
.D(n_109),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_150),
.A3(n_146),
.B1(n_145),
.B2(n_147),
.C1(n_59),
.C2(n_66),
.Y(n_157)
);

BUFx4f_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_59),
.A3(n_151),
.B1(n_93),
.B2(n_71),
.C1(n_60),
.C2(n_106),
.Y(n_159)
);

OAI31xp33_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_155),
.A3(n_153),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_156),
.B1(n_105),
.B2(n_101),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_71),
.B(n_17),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_163),
.B(n_160),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_165),
.B1(n_162),
.B2(n_160),
.C(n_164),
.Y(n_167)
);


endmodule