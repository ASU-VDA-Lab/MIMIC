module fake_ariane_3235_n_1940 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1940);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1940;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_206;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_261;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_1524;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1759;
wire n_1557;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_82),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_31),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_47),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_65),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_75),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_115),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_28),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_71),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_48),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_59),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_123),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

BUFx8_ASAP7_75t_SL g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_141),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_68),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_12),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_54),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_33),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_128),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_20),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_44),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_96),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_76),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_50),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_30),
.Y(n_215)
);

CKINVDCx12_ASAP7_75t_R g216 ( 
.A(n_62),
.Y(n_216)
);

INVx4_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_25),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_36),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_57),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_130),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_131),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_19),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_66),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_24),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_114),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_38),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_51),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_36),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_107),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_20),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_26),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_83),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_21),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_149),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_22),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_3),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_64),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_135),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_153),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_106),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_45),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_13),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_63),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_103),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_92),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_108),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_91),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_146),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_26),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_119),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_8),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_80),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_0),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_89),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_46),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_35),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_10),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_105),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_117),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_10),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_35),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_2),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_39),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_25),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_40),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_22),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

BUFx2_ASAP7_75t_SL g303 ( 
.A(n_11),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_142),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_49),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_4),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_38),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_31),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_15),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_74),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_53),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_188),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_229),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_164),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_307),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_174),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_211),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_221),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_228),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_237),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_297),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_249),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_219),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_219),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_179),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_275),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_288),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_162),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_190),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_167),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_204),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_193),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_197),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_159),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_199),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_172),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_184),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_184),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_212),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_240),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_247),
.Y(n_363)
);

BUFx2_ASAP7_75t_SL g364 ( 
.A(n_194),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_216),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_260),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_262),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_179),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_264),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_215),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_223),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_285),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_194),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_198),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_226),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_161),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_168),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_198),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_257),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_173),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_257),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_322),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

NAND2x1p5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_195),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_195),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_325),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_324),
.A2(n_189),
.B(n_183),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_194),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_389),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_234),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_329),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_196),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

NAND2x1_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_217),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_200),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_357),
.B(n_279),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_337),
.B(n_369),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_330),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_368),
.B(n_279),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_340),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_337),
.B(n_205),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_360),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_335),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_314),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_377),
.B(n_207),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_385),
.B(n_386),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_347),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_336),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_317),
.B(n_279),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_338),
.A2(n_210),
.B(n_218),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_341),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_169),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_319),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_441),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_426),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_444),
.A2(n_364),
.B1(n_352),
.B2(n_234),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_392),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_407),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_406),
.B(n_351),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_396),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_406),
.B(n_399),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_391),
.Y(n_478)
);

HB1xp67_ASAP7_75t_SL g479 ( 
.A(n_401),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_353),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_358),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

BUFx6f_ASAP7_75t_SL g486 ( 
.A(n_444),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_441),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_426),
.A2(n_376),
.B1(n_332),
.B2(n_339),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_449),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_427),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_420),
.B(n_303),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_398),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_395),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

INVx11_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

BUFx6f_ASAP7_75t_SL g512 ( 
.A(n_444),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_398),
.Y(n_514)
);

BUFx6f_ASAP7_75t_SL g515 ( 
.A(n_411),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_449),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_400),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_399),
.A2(n_222),
.B1(n_159),
.B2(n_287),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_407),
.B(n_323),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_398),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_457),
.B(n_230),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_400),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_371),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_403),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_408),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_410),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_398),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_409),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_417),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_456),
.B(n_331),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_452),
.A2(n_363),
.B1(n_378),
.B2(n_348),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_409),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_452),
.B(n_232),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_345),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_373),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_457),
.B(n_380),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_419),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_445),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_445),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_445),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_412),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_421),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_415),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_423),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_404),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_425),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_456),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_425),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_437),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_429),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_404),
.B(n_239),
.C(n_235),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_433),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_450),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_442),
.B(n_366),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_458),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_451),
.B(n_158),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_450),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_435),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_451),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_442),
.B(n_432),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_428),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_430),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_439),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_451),
.B(n_346),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_432),
.B(n_349),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_411),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_430),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_404),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_424),
.Y(n_601)
);

OA22x2_ASAP7_75t_L g602 ( 
.A1(n_422),
.A2(n_370),
.B1(n_372),
.B2(n_374),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_431),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_450),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_422),
.B(n_361),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_435),
.B(n_320),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_448),
.B(n_361),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_450),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_499),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_460),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_460),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_500),
.B(n_448),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_447),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_463),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_472),
.B(n_411),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_573),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_472),
.B(n_411),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_463),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_461),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_326),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_526),
.B(n_527),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_498),
.B(n_343),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_527),
.B(n_404),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_473),
.B(n_344),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_411),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_589),
.B(n_158),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_485),
.B(n_362),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_563),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_578),
.A2(n_418),
.B(n_431),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_464),
.B(n_362),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_597),
.B(n_365),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_529),
.B(n_404),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_517),
.B(n_171),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_477),
.B(n_447),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_511),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_590),
.B(n_434),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_461),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_576),
.B(n_418),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_483),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_365),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_521),
.B(n_367),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_493),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_530),
.B(n_452),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_493),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_497),
.B(n_434),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_531),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_453),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_539),
.B(n_438),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_531),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_533),
.B(n_452),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_462),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_452),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_589),
.B(n_438),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_543),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_534),
.B(n_447),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_534),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_536),
.Y(n_667)
);

NAND3x1_ASAP7_75t_L g668 ( 
.A(n_519),
.B(n_375),
.C(n_367),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_466),
.Y(n_669)
);

NAND3x1_ASAP7_75t_L g670 ( 
.A(n_519),
.B(n_379),
.C(n_375),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_496),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_536),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_502),
.A2(n_185),
.B1(n_236),
.B2(n_238),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_588),
.B(n_160),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_466),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_381),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_552),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_539),
.B(n_453),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_596),
.A2(n_579),
.B1(n_523),
.B2(n_287),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_468),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_606),
.B(n_439),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_605),
.B(n_447),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_479),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_539),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_544),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_515),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_595),
.A2(n_309),
.B1(n_293),
.B2(n_308),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_502),
.A2(n_522),
.B1(n_535),
.B2(n_514),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_598),
.B(n_455),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_598),
.B(n_455),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_515),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_480),
.B(n_440),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_552),
.B(n_439),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_566),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_517),
.B(n_382),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_556),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_595),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_556),
.B(n_415),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_583),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

NAND2x1p5_ASAP7_75t_L g705 ( 
.A(n_525),
.B(n_440),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_525),
.B(n_549),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_171),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_515),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_486),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_481),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_557),
.B(n_415),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_486),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_588),
.B(n_160),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_468),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_559),
.B(n_415),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_584),
.B(n_454),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_470),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_559),
.B(n_436),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_523),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_564),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_588),
.B(n_163),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_470),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_564),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_478),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_585),
.B(n_293),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_588),
.B(n_295),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_584),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_486),
.B(n_295),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_514),
.B(n_163),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_478),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_481),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_602),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_549),
.B(n_440),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_549),
.B(n_446),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_488),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_522),
.B(n_165),
.Y(n_736)
);

INVx8_ASAP7_75t_L g737 ( 
.A(n_512),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_565),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_565),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_575),
.Y(n_740)
);

AO21x2_ASAP7_75t_L g741 ( 
.A1(n_578),
.A2(n_281),
.B(n_251),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_488),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_501),
.B(n_446),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_SL g744 ( 
.A1(n_465),
.A2(n_308),
.B1(n_309),
.B2(n_241),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_567),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_607),
.B(n_446),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_567),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_584),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_584),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_602),
.A2(n_263),
.B1(n_231),
.B2(n_244),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_501),
.B(n_454),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_513),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_568),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_512),
.B(n_246),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_575),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_575),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_568),
.B(n_436),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_571),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_490),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_501),
.B(n_454),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_501),
.B(n_436),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_490),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_575),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_491),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_571),
.B(n_574),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_574),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_491),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_523),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_501),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_592),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_494),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_513),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_512),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_592),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_494),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_503),
.Y(n_778)
);

INVx4_ASAP7_75t_SL g779 ( 
.A(n_523),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_513),
.B(n_248),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_513),
.B(n_258),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_631),
.Y(n_782)
);

BUFx6f_ASAP7_75t_SL g783 ( 
.A(n_669),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_710),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_618),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_621),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_752),
.B(n_535),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_641),
.B(n_593),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_654),
.B(n_593),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_687),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_645),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_640),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_690),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_656),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_710),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_726),
.A2(n_523),
.B1(n_482),
.B2(n_602),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_690),
.B(n_599),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_731),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_659),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_742),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_666),
.B(n_667),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_672),
.B(n_599),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_678),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_706),
.B(n_603),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_R g806 ( 
.A(n_676),
.B(n_523),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_703),
.A2(n_523),
.B1(n_553),
.B2(n_603),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_693),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_699),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_742),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_618),
.B(n_278),
.C(n_274),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_615),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_706),
.B(n_545),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_623),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_704),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_752),
.B(n_551),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_759),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_748),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_640),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_694),
.B(n_541),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_680),
.A2(n_476),
.B(n_459),
.C(n_489),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_625),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_687),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_720),
.B(n_459),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_723),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_671),
.A2(n_548),
.B1(n_283),
.B2(n_284),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_SL g827 ( 
.A(n_688),
.B(n_286),
.C(n_166),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_638),
.B(n_601),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_759),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_773),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_698),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_774),
.B(n_551),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_738),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_739),
.B(n_469),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_778),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_630),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_650),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_774),
.B(n_551),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_687),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_745),
.B(n_747),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_680),
.B(n_572),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_663),
.B(n_469),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_753),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_684),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_612),
.B(n_471),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_758),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_778),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_766),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_671),
.A2(n_548),
.B1(n_600),
.B2(n_570),
.Y(n_850)
);

AND2x4_ASAP7_75t_SL g851 ( 
.A(n_694),
.B(n_570),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_780),
.A2(n_475),
.B(n_505),
.C(n_504),
.Y(n_852)
);

BUFx4f_ASAP7_75t_L g853 ( 
.A(n_737),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_769),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_708),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_781),
.A2(n_548),
.B1(n_600),
.B2(n_570),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_617),
.B(n_471),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_771),
.B(n_475),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_772),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_749),
.B(n_716),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_776),
.B(n_476),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_650),
.Y(n_862)
);

NAND2x1_ASAP7_75t_L g863 ( 
.A(n_658),
.B(n_489),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_624),
.B(n_495),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_744),
.A2(n_570),
.B1(n_600),
.B2(n_541),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_677),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_610),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_624),
.B(n_495),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_611),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_622),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_643),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_749),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_644),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_614),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_708),
.B(n_638),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_SL g876 ( 
.A(n_627),
.B(n_166),
.C(n_165),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_634),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_744),
.A2(n_600),
.B1(n_547),
.B2(n_550),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_646),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_732),
.A2(n_550),
.B1(n_547),
.B2(n_503),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_765),
.B(n_504),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_646),
.B(n_467),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_661),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_655),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_638),
.B(n_572),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_677),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_765),
.B(n_505),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_617),
.B(n_487),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_619),
.B(n_487),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_657),
.A2(n_572),
.B1(n_594),
.B2(n_538),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_646),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_705),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_700),
.B(n_664),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_675),
.B(n_594),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_675),
.B(n_594),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_750),
.A2(n_608),
.B1(n_604),
.B2(n_555),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_675),
.B(n_467),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_700),
.B(n_728),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_754),
.B(n_467),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_647),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_619),
.B(n_487),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_633),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_709),
.B(n_555),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_737),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_685),
.B(n_467),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_743),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_639),
.B(n_608),
.C(n_604),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_709),
.B(n_558),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_634),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_685),
.B(n_484),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_628),
.B(n_484),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_649),
.Y(n_912)
);

AND2x6_ASAP7_75t_SL g913 ( 
.A(n_725),
.B(n_252),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_SL g914 ( 
.A(n_673),
.B(n_291),
.C(n_182),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_727),
.B(n_484),
.Y(n_915)
);

INVx5_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_642),
.B(n_492),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_647),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_649),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_712),
.B(n_558),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_642),
.B(n_492),
.Y(n_921)
);

NOR2x2_ASAP7_75t_L g922 ( 
.A(n_743),
.B(n_560),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_707),
.B(n_484),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_642),
.B(n_492),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_665),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_668),
.A2(n_516),
.B1(n_518),
.B2(n_528),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_642),
.B(n_633),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_750),
.A2(n_628),
.B1(n_760),
.B2(n_751),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_681),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_673),
.B(n_516),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_614),
.B(n_620),
.Y(n_931)
);

BUFx4f_ASAP7_75t_L g932 ( 
.A(n_737),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_629),
.B(n_516),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_691),
.B(n_518),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_712),
.B(n_560),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_692),
.B(n_518),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_609),
.B(n_616),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_626),
.A2(n_528),
.B(n_538),
.C(n_546),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_733),
.B(n_561),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_746),
.B(n_528),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_683),
.B(n_538),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_636),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_658),
.B(n_546),
.Y(n_943)
);

CKINVDCx11_ASAP7_75t_R g944 ( 
.A(n_775),
.Y(n_944)
);

AO22x1_ASAP7_75t_L g945 ( 
.A1(n_770),
.A2(n_170),
.B1(n_182),
.B2(n_313),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_682),
.B(n_436),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_665),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_751),
.A2(n_561),
.B1(n_591),
.B2(n_587),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_658),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_614),
.B(n_546),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_761),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_620),
.B(n_506),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_620),
.B(n_506),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_637),
.B(n_507),
.Y(n_954)
);

AND3x1_ASAP7_75t_L g955 ( 
.A(n_696),
.B(n_540),
.C(n_507),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_658),
.B(n_508),
.Y(n_956)
);

CKINVDCx11_ASAP7_75t_R g957 ( 
.A(n_637),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_729),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_733),
.B(n_562),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_734),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_637),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_679),
.B(n_508),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_714),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_651),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_670),
.B(n_562),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_679),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_679),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_717),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_734),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_760),
.A2(n_569),
.B1(n_591),
.B2(n_587),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_679),
.B(n_509),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_651),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_722),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_701),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_898),
.B(n_674),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_786),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_785),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_867),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_902),
.Y(n_979)
);

BUFx8_ASAP7_75t_L g980 ( 
.A(n_783),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_869),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_794),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_840),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_925),
.B(n_695),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_785),
.B(n_651),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_949),
.B(n_761),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_805),
.B(n_779),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_884),
.B(n_713),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_800),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_804),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_902),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_949),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_812),
.B(n_721),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_870),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_809),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_837),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_871),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_852),
.A2(n_701),
.B(n_757),
.C(n_718),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_768),
.B(n_757),
.C(n_718),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_923),
.A2(n_711),
.B(n_715),
.C(n_736),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_947),
.B(n_735),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_864),
.A2(n_635),
.B(n_626),
.Y(n_1003)
);

INVx3_ASAP7_75t_SL g1004 ( 
.A(n_782),
.Y(n_1004)
);

AOI22x1_ASAP7_75t_L g1005 ( 
.A1(n_974),
.A2(n_825),
.B1(n_834),
.B2(n_815),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_793),
.B(n_762),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_872),
.B(n_697),
.Y(n_1007)
);

AOI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_914),
.A2(n_289),
.B1(n_255),
.B2(n_256),
.C(n_269),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_883),
.Y(n_1009)
);

BUFx5_ASAP7_75t_L g1010 ( 
.A(n_939),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_844),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_826),
.A2(n_813),
.B1(n_814),
.B2(n_831),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_929),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_963),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_821),
.A2(n_715),
.B(n_711),
.C(n_696),
.Y(n_1015)
);

CKINVDCx16_ASAP7_75t_R g1016 ( 
.A(n_783),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_893),
.B(n_613),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_847),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_894),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_864),
.B(n_764),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_805),
.B(n_779),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_966),
.B(n_697),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_813),
.A2(n_719),
.B1(n_777),
.B2(n_767),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_808),
.B(n_697),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_849),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_868),
.B(n_635),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_894),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_854),
.Y(n_1028)
);

INVxp33_ASAP7_75t_L g1029 ( 
.A(n_791),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_868),
.B(n_724),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_968),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_827),
.A2(n_300),
.B1(n_652),
.B2(n_660),
.C(n_662),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_912),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_838),
.B(n_702),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_966),
.B(n_702),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_859),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_802),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_862),
.B(n_702),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_802),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_790),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_866),
.B(n_648),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_841),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_840),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_790),
.B(n_648),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_L g1045 ( 
.A(n_944),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_886),
.A2(n_653),
.B1(n_686),
.B2(n_689),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_841),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_957),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_973),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_881),
.B(n_730),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_790),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_845),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_822),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_966),
.B(n_653),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_784),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_879),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_881),
.B(n_652),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_919),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_967),
.B(n_686),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_937),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_887),
.B(n_660),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_876),
.A2(n_686),
.B1(n_689),
.B2(n_662),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_877),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_909),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_887),
.A2(n_843),
.B(n_938),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_824),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_967),
.B(n_689),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_788),
.A2(n_763),
.B1(n_756),
.B2(n_755),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_824),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_818),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_840),
.Y(n_1071)
);

AND2x6_ASAP7_75t_L g1072 ( 
.A(n_875),
.B(n_740),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_895),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_835),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_961),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_835),
.Y(n_1076)
);

INVxp67_ASAP7_75t_SL g1077 ( 
.A(n_969),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_788),
.A2(n_789),
.B1(n_803),
.B2(n_858),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_895),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_960),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_964),
.Y(n_1081)
);

AND3x2_ASAP7_75t_SL g1082 ( 
.A(n_913),
.B(n_586),
.C(n_582),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_823),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_904),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_899),
.A2(n_582),
.B(n_569),
.C(n_577),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_951),
.B(n_632),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_789),
.B(n_632),
.Y(n_1087)
);

AO22x1_ASAP7_75t_L g1088 ( 
.A1(n_875),
.A2(n_181),
.B1(n_180),
.B2(n_170),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_967),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_823),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_823),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_858),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_891),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_803),
.B(n_740),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_853),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_969),
.B(n_741),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_846),
.B(n_740),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_861),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_939),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_861),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_951),
.B(n_755),
.Y(n_1101)
);

CKINVDCx11_ASAP7_75t_R g1102 ( 
.A(n_874),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_795),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_853),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_797),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_906),
.B(n_763),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_SL g1107 ( 
.A1(n_798),
.A2(n_741),
.B1(n_224),
.B2(n_181),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_799),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_906),
.B(n_755),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_906),
.B(n_763),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_939),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_801),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_960),
.B(n_756),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_810),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_927),
.A2(n_175),
.B1(n_180),
.B2(n_291),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_927),
.B(n_756),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_932),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_817),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_807),
.B(n_577),
.C(n_586),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_939),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_959),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_828),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_928),
.A2(n_580),
.B1(n_537),
.B2(n_532),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_811),
.A2(n_178),
.B1(n_176),
.B2(n_175),
.C(n_294),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_922),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_959),
.Y(n_1126)
);

AND2x6_ASAP7_75t_L g1127 ( 
.A(n_792),
.B(n_580),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_798),
.B(n_509),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_798),
.B(n_510),
.Y(n_1129)
);

AND2x4_ASAP7_75t_SL g1130 ( 
.A(n_1117),
.B(n_972),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_977),
.B(n_945),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_975),
.B(n_874),
.Y(n_1132)
);

AO22x1_ASAP7_75t_L g1133 ( 
.A1(n_980),
.A2(n_855),
.B1(n_916),
.B2(n_942),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1111),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_978),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_981),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1045),
.Y(n_1137)
);

INVx5_ASAP7_75t_L g1138 ( 
.A(n_1113),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1102),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1111),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1117),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1008),
.A2(n_798),
.B1(n_965),
.B2(n_860),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_987),
.B(n_916),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_1113),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1078),
.A2(n_941),
.B(n_890),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1052),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1037),
.B(n_850),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1078),
.A2(n_856),
.B1(n_857),
.B2(n_878),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1039),
.B(n_940),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_1017),
.Y(n_1151)
);

OAI33xp33_ASAP7_75t_L g1152 ( 
.A1(n_1060),
.A2(n_958),
.A3(n_930),
.B1(n_890),
.B2(n_888),
.B3(n_889),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1111),
.B(n_916),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1033),
.B(n_892),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1008),
.A2(n_842),
.B1(n_955),
.B2(n_940),
.C(n_880),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1042),
.B(n_874),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1111),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_994),
.Y(n_1158)
);

NAND2x1p5_ASAP7_75t_L g1159 ( 
.A(n_1099),
.B(n_1120),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1012),
.A2(n_965),
.B1(n_806),
.B2(n_820),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_976),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1058),
.B(n_888),
.Y(n_1162)
);

BUFx8_ASAP7_75t_SL g1163 ( 
.A(n_1070),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_997),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1075),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_999),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_982),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1107),
.A2(n_965),
.B1(n_820),
.B2(n_848),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1032),
.A2(n_865),
.B1(n_882),
.B2(n_955),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_996),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1026),
.A2(n_941),
.B(n_921),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1026),
.A2(n_921),
.B(n_917),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_988),
.B(n_972),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1004),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1009),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1013),
.Y(n_1176)
);

AOI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_946),
.B(n_907),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_980),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1014),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1057),
.A2(n_924),
.B(n_917),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_987),
.B(n_855),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1081),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1029),
.B(n_972),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_989),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_L g1185 ( 
.A(n_1127),
.B(n_792),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1031),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1047),
.B(n_934),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1077),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_986),
.B(n_903),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1126),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_990),
.Y(n_1191)
);

CKINVDCx11_ASAP7_75t_R g1192 ( 
.A(n_1016),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1117),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1021),
.B(n_855),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1053),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1056),
.B(n_1024),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1083),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_L g1198 ( 
.A(n_1104),
.B(n_931),
.Y(n_1198)
);

CKINVDCx8_ASAP7_75t_R g1199 ( 
.A(n_979),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1084),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1049),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_986),
.B(n_903),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1083),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1066),
.B(n_936),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_995),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_926),
.B1(n_889),
.B2(n_901),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1011),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1018),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1074),
.A2(n_787),
.B1(n_911),
.B2(n_933),
.Y(n_1209)
);

AND2x2_ASAP7_75t_SL g1210 ( 
.A(n_991),
.B(n_932),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1113),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1025),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1007),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1082),
.A2(n_935),
.B1(n_908),
.B2(n_920),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1028),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1036),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1063),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1126),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1099),
.B(n_1120),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1095),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1021),
.B(n_908),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1083),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1071),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_983),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1064),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1112),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1077),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1114),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1034),
.B(n_920),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_983),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1055),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1113),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1076),
.B(n_829),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1057),
.A2(n_1061),
.B(n_1065),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1038),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_983),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1103),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1072),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_986),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1105),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1106),
.B(n_935),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1108),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1118),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1090),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1106),
.B(n_828),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1092),
.A2(n_915),
.B1(n_839),
.B2(n_816),
.Y(n_1246)
);

AO22x1_ASAP7_75t_L g1247 ( 
.A1(n_1125),
.A2(n_832),
.B1(n_830),
.B2(n_836),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1006),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1043),
.Y(n_1249)
);

AOI222xp33_ASAP7_75t_L g1250 ( 
.A1(n_1124),
.A2(n_176),
.B1(n_306),
.B2(n_305),
.C1(n_304),
.C2(n_178),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1098),
.B(n_924),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1006),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1100),
.B(n_833),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1090),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_984),
.B(n_956),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1072),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1002),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1072),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1002),
.Y(n_1259)
);

AO22x1_ASAP7_75t_L g1260 ( 
.A1(n_1125),
.A2(n_993),
.B1(n_1082),
.B2(n_1044),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1121),
.B(n_896),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_984),
.B(n_956),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1090),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1019),
.B(n_851),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1093),
.B(n_2),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1005),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1094),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1072),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1043),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1107),
.A2(n_1124),
.B1(n_1094),
.B2(n_1086),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1043),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1080),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1061),
.B(n_962),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1088),
.A2(n_294),
.B1(n_305),
.B2(n_306),
.C(n_313),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1020),
.B(n_962),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1080),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1020),
.B(n_948),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1019),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1096),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1109),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1041),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1001),
.A2(n_950),
.B(n_885),
.C(n_943),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1027),
.B(n_819),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1027),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1250),
.A2(n_1023),
.B1(n_1087),
.B2(n_1030),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1149),
.A2(n_1000),
.B(n_1068),
.C(n_1015),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1260),
.B(n_1128),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1205),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1266),
.A2(n_1065),
.B(n_1068),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1234),
.A2(n_1003),
.B(n_1087),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1149),
.A2(n_1010),
.B1(n_1050),
.B2(n_1030),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1180),
.A2(n_1003),
.B(n_1128),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1216),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_1188),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1177),
.A2(n_907),
.B(n_1119),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1138),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1129),
.B(n_998),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1138),
.B(n_1109),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1171),
.A2(n_1129),
.B(n_998),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1146),
.A2(n_1119),
.B(n_1085),
.Y(n_1300)
);

BUFx12f_ASAP7_75t_L g1301 ( 
.A(n_1192),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1171),
.A2(n_1097),
.B(n_1050),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1177),
.A2(n_1097),
.B(n_1062),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1248),
.A2(n_971),
.A3(n_943),
.B(n_540),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1151),
.B(n_1131),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1238),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1169),
.A2(n_1116),
.B(n_952),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1252),
.B(n_1073),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1189),
.B(n_1110),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1169),
.A2(n_1115),
.B(n_1123),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1200),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1161),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1167),
.Y(n_1313)
);

BUFx5_ASAP7_75t_L g1314 ( 
.A(n_1267),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1238),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1241),
.B(n_1110),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1213),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1172),
.A2(n_953),
.B(n_954),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1184),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1148),
.A2(n_905),
.B(n_910),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1282),
.A2(n_1275),
.B(n_1141),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1138),
.B(n_1089),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1196),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1145),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1191),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1275),
.A2(n_863),
.B(n_1089),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1270),
.A2(n_985),
.B(n_1059),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1268),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1134),
.A2(n_1122),
.B(n_992),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1207),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1227),
.Y(n_1331)
);

BUFx8_ASAP7_75t_L g1332 ( 
.A(n_1139),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1250),
.A2(n_1079),
.B1(n_1073),
.B2(n_1010),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1201),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1268),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1270),
.A2(n_1067),
.B(n_1035),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1134),
.A2(n_1122),
.B(n_992),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1163),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1257),
.B(n_1079),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1143),
.A2(n_1155),
.B1(n_1145),
.B2(n_1209),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1259),
.B(n_1010),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1206),
.A2(n_1046),
.B(n_897),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1272),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1185),
.A2(n_1022),
.B(n_1054),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1274),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.C(n_270),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1151),
.B(n_1051),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1145),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1208),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1212),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1215),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1235),
.B(n_1101),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_SL g1352 ( 
.A1(n_1204),
.A2(n_1091),
.B(n_1040),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1143),
.A2(n_542),
.B(n_537),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1141),
.A2(n_510),
.B(n_520),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1237),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1217),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1211),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1148),
.A2(n_542),
.B(n_532),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_524),
.B(n_520),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1274),
.B(n_301),
.C(n_302),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1187),
.A2(n_524),
.B(n_918),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1225),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1226),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1155),
.A2(n_1277),
.B(n_1273),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1157),
.A2(n_918),
.B(n_819),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_L g1366 ( 
.A(n_1173),
.B(n_1040),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1206),
.A2(n_1127),
.B(n_970),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1147),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1228),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1277),
.A2(n_1010),
.B(n_1044),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1223),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1157),
.A2(n_900),
.B(n_1010),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1273),
.A2(n_250),
.B(n_191),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1240),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1220),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1187),
.A2(n_254),
.B(n_192),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1231),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1255),
.A2(n_1091),
.A3(n_1127),
.B(n_424),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1255),
.A2(n_1127),
.A3(n_424),
.B(n_437),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_1154),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1150),
.B(n_575),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1251),
.A2(n_214),
.B(n_225),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1135),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1136),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1150),
.A2(n_253),
.B(n_201),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1251),
.A2(n_900),
.B(n_437),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_SL g1387 ( 
.A(n_1140),
.Y(n_1387)
);

BUFx2_ASAP7_75t_R g1388 ( 
.A(n_1178),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1132),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1137),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1189),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1195),
.B(n_6),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1276),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1262),
.A2(n_437),
.B(n_424),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1242),
.Y(n_1395)
);

INVx8_ASAP7_75t_L g1396 ( 
.A(n_1222),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1243),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1158),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1164),
.Y(n_1399)
);

CKINVDCx14_ASAP7_75t_R g1400 ( 
.A(n_1139),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1211),
.B(n_601),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1262),
.A2(n_1159),
.B(n_1219),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1159),
.A2(n_437),
.B(n_424),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1166),
.Y(n_1404)
);

OAI222xp33_ASAP7_75t_L g1405 ( 
.A1(n_1261),
.A2(n_273),
.B1(n_203),
.B2(n_186),
.C1(n_208),
.C2(n_209),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1170),
.B(n_437),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1263),
.Y(n_1407)
);

OAI221xp5_ASAP7_75t_L g1408 ( 
.A1(n_1209),
.A2(n_206),
.B1(n_213),
.B2(n_227),
.C(n_233),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1246),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1175),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1279),
.A2(n_424),
.A3(n_437),
.B(n_601),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1232),
.Y(n_1412)
);

AO21x1_ASAP7_75t_L g1413 ( 
.A1(n_1156),
.A2(n_424),
.B(n_15),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1199),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1176),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1219),
.A2(n_1239),
.B(n_1253),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1239),
.A2(n_424),
.B(n_601),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1253),
.A2(n_601),
.B(n_282),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1233),
.A2(n_601),
.B(n_102),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1179),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1246),
.A2(n_277),
.B(n_272),
.Y(n_1421)
);

AOI22x1_ASAP7_75t_SL g1422 ( 
.A1(n_1271),
.A2(n_271),
.B1(n_267),
.B2(n_266),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1186),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1233),
.A2(n_70),
.B(n_156),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1139),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1152),
.A2(n_265),
.B(n_261),
.Y(n_1426)
);

BUFx8_ASAP7_75t_L g1427 ( 
.A(n_1165),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1142),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1162),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1210),
.B(n_7),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1232),
.A2(n_69),
.B(n_155),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1153),
.A2(n_67),
.B(n_152),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1390),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1340),
.A2(n_1281),
.B1(n_1160),
.B2(n_1214),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1393),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1368),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1391),
.B(n_1202),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1340),
.A2(n_1229),
.B1(n_1168),
.B2(n_1190),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_SL g1439 ( 
.A(n_1345),
.B(n_1265),
.C(n_1182),
.Y(n_1439)
);

AO22x2_ASAP7_75t_L g1440 ( 
.A1(n_1288),
.A2(n_1190),
.B1(n_1218),
.B2(n_1174),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1334),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1373),
.A2(n_1218),
.B1(n_1258),
.B2(n_1256),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1310),
.A2(n_1221),
.B1(n_1241),
.B2(n_1202),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1311),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1311),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1409),
.A2(n_1183),
.B1(n_1247),
.B2(n_1133),
.C(n_1278),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1323),
.B(n_1284),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1373),
.A2(n_1258),
.B1(n_1256),
.B2(n_1189),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1293),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1409),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.C(n_1142),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1333),
.A2(n_1202),
.B1(n_1221),
.B2(n_1194),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1310),
.A2(n_1241),
.B1(n_1144),
.B2(n_1280),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

AND2x6_ASAP7_75t_L g1454 ( 
.A(n_1296),
.B(n_1264),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1333),
.A2(n_1144),
.B1(n_1280),
.B2(n_1198),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1287),
.B(n_1153),
.Y(n_1456)
);

NAND2xp33_ASAP7_75t_L g1457 ( 
.A(n_1314),
.B(n_1193),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1429),
.B(n_1203),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1396),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1312),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1355),
.Y(n_1461)
);

AND2x2_ASAP7_75t_SL g1462 ( 
.A(n_1296),
.B(n_1181),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1408),
.A2(n_1193),
.B1(n_1142),
.B2(n_1245),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1391),
.B(n_1280),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1313),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1305),
.B(n_1230),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1374),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1408),
.A2(n_1283),
.B1(n_1264),
.B2(n_1193),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1400),
.A2(n_1430),
.B1(n_1392),
.B2(n_1291),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1345),
.A2(n_1181),
.B1(n_1194),
.B2(n_1283),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1405),
.A2(n_1269),
.B1(n_1236),
.B2(n_1249),
.C(n_1224),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1376),
.A2(n_1245),
.B1(n_1254),
.B2(n_1244),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1301),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1380),
.B(n_1317),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1332),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1357),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1319),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1373),
.A2(n_1245),
.B1(n_1254),
.B2(n_1244),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1380),
.B(n_1346),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1376),
.A2(n_1254),
.B1(n_1244),
.B2(n_1203),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_SL g1481 ( 
.A1(n_1421),
.A2(n_1203),
.B(n_1197),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1430),
.A2(n_1130),
.B1(n_1197),
.B2(n_19),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1357),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1343),
.B(n_1325),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1383),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1421),
.A2(n_1197),
.B1(n_18),
.B2(n_23),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1343),
.B(n_17),
.Y(n_1487)
);

NAND2xp33_ASAP7_75t_SL g1488 ( 
.A(n_1371),
.B(n_1390),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1330),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1382),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1385),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1348),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1349),
.B(n_27),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1360),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.C(n_40),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1385),
.A2(n_37),
.B1(n_52),
.B2(n_60),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1332),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1389),
.B(n_78),
.C(n_94),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1294),
.B(n_98),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1382),
.A2(n_1364),
.B1(n_1285),
.B2(n_1287),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1350),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1391),
.B(n_116),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1294),
.B(n_1331),
.Y(n_1502)
);

AO21x1_ASAP7_75t_L g1503 ( 
.A1(n_1389),
.A2(n_122),
.B(n_129),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1291),
.A2(n_133),
.B1(n_145),
.B2(n_1285),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1331),
.B(n_1356),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1396),
.B(n_1425),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1391),
.B(n_1309),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1382),
.A2(n_1364),
.B1(n_1287),
.B2(n_1367),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1289),
.A2(n_1386),
.B(n_1290),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1384),
.Y(n_1511)
);

AO31x2_ASAP7_75t_L g1512 ( 
.A1(n_1341),
.A2(n_1361),
.A3(n_1377),
.B(n_1397),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1363),
.B(n_1369),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1412),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1339),
.B(n_1308),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1286),
.B(n_1392),
.C(n_1300),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1405),
.A2(n_1286),
.B(n_1321),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1396),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1367),
.A2(n_1420),
.B1(n_1410),
.B2(n_1415),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1339),
.B(n_1308),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1395),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1400),
.A2(n_1300),
.B1(n_1328),
.B2(n_1306),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1338),
.Y(n_1523)
);

AOI22x1_ASAP7_75t_L g1524 ( 
.A1(n_1352),
.A2(n_1328),
.B1(n_1315),
.B2(n_1335),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1414),
.B(n_1422),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1398),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1399),
.A2(n_1423),
.B1(n_1404),
.B2(n_1327),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1336),
.A2(n_1327),
.B1(n_1316),
.B2(n_1309),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1309),
.B(n_1296),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1358),
.A2(n_1418),
.B(n_1353),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1299),
.A2(n_1297),
.B(n_1292),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1341),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1306),
.A2(n_1335),
.B1(n_1315),
.B2(n_1407),
.Y(n_1533)
);

INVx6_ASAP7_75t_L g1534 ( 
.A(n_1427),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1407),
.A2(n_1351),
.B1(n_1342),
.B2(n_1366),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1314),
.Y(n_1536)
);

AND2x6_ASAP7_75t_L g1537 ( 
.A(n_1296),
.B(n_1347),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1381),
.B(n_1427),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1314),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1314),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1314),
.Y(n_1541)
);

BUFx4f_ASAP7_75t_SL g1542 ( 
.A(n_1428),
.Y(n_1542)
);

AND2x6_ASAP7_75t_L g1543 ( 
.A(n_1324),
.B(n_1347),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1412),
.Y(n_1544)
);

BUFx10_ASAP7_75t_L g1545 ( 
.A(n_1388),
.Y(n_1545)
);

AO21x1_ASAP7_75t_SL g1546 ( 
.A1(n_1342),
.A2(n_1381),
.B(n_1406),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_SL g1547 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1344),
.C(n_1426),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1336),
.A2(n_1418),
.B1(n_1370),
.B2(n_1307),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1370),
.A2(n_1307),
.B1(n_1314),
.B2(n_1303),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1316),
.B(n_1402),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1387),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1324),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1324),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1320),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1324),
.B(n_1347),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1502),
.B(n_1302),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1436),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1516),
.A2(n_1426),
.B(n_1361),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1516),
.A2(n_1320),
.B1(n_1303),
.B2(n_1344),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1456),
.B(n_1347),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1504),
.A2(n_1416),
.B(n_1424),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1435),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1453),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_R g1564 ( 
.A(n_1506),
.B(n_1302),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1523),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1486),
.A2(n_1359),
.B1(n_1322),
.B2(n_1298),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1486),
.A2(n_1359),
.B1(n_1322),
.B2(n_1298),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_SL g1568 ( 
.A(n_1546),
.B(n_1353),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1474),
.B(n_1378),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1532),
.B(n_1304),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_1433),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1479),
.B(n_1378),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1515),
.B(n_1520),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1456),
.B(n_1326),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1545),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1449),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1456),
.B(n_1432),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1484),
.B(n_1304),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1513),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1508),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1526),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1466),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1447),
.B(n_1378),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1444),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1445),
.B(n_1550),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1441),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1552),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_R g1588 ( 
.A(n_1506),
.B(n_1431),
.Y(n_1588)
);

NAND2xp33_ASAP7_75t_R g1589 ( 
.A(n_1501),
.B(n_1329),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1444),
.B(n_1378),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1501),
.B(n_1337),
.Y(n_1591)
);

CKINVDCx14_ASAP7_75t_R g1592 ( 
.A(n_1545),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_SL g1593 ( 
.A(n_1482),
.B(n_1413),
.C(n_1401),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1505),
.B(n_1304),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1473),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_R g1596 ( 
.A(n_1488),
.B(n_1379),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1475),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1512),
.B(n_1304),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1512),
.B(n_1295),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1469),
.A2(n_1295),
.B1(n_1358),
.B2(n_1318),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1512),
.B(n_1379),
.Y(n_1601)
);

NOR3xp33_ASAP7_75t_SL g1602 ( 
.A(n_1533),
.B(n_1365),
.C(n_1419),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1528),
.B(n_1507),
.Y(n_1603)
);

CKINVDCx8_ASAP7_75t_R g1604 ( 
.A(n_1525),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1528),
.B(n_1379),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1460),
.B(n_1379),
.Y(n_1606)
);

CKINVDCx11_ASAP7_75t_R g1607 ( 
.A(n_1496),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1439),
.A2(n_1372),
.B(n_1403),
.C(n_1394),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1465),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1521),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1538),
.B(n_1318),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1476),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1477),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1507),
.B(n_1354),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1489),
.B(n_1411),
.Y(n_1615)
);

AO31x2_ASAP7_75t_L g1616 ( 
.A1(n_1503),
.A2(n_1411),
.A3(n_1417),
.B(n_1401),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_SL g1617 ( 
.A(n_1522),
.B(n_1411),
.C(n_1487),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_R g1618 ( 
.A(n_1493),
.B(n_1411),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1492),
.B(n_1500),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1461),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1544),
.B(n_1440),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1458),
.B(n_1554),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1440),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1476),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1483),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1467),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1483),
.B(n_1514),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1485),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1475),
.Y(n_1629)
);

OR2x6_ASAP7_75t_L g1630 ( 
.A(n_1529),
.B(n_1437),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1509),
.B(n_1499),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1511),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1621),
.B(n_1539),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1624),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1563),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1611),
.A2(n_1469),
.B1(n_1494),
.B2(n_1517),
.C(n_1450),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1599),
.A2(n_1549),
.B(n_1548),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1585),
.B(n_1536),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1562),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1583),
.B(n_1540),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1576),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1625),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1622),
.B(n_1541),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1609),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1573),
.B(n_1514),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1556),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1593),
.A2(n_1482),
.B1(n_1470),
.B2(n_1451),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1586),
.Y(n_1648)
);

NAND2x1_ASAP7_75t_L g1649 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1569),
.B(n_1572),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1556),
.B(n_1518),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1579),
.B(n_1531),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1617),
.B(n_1490),
.C(n_1491),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1571),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1619),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1620),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1632),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1580),
.B(n_1510),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1590),
.B(n_1510),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1603),
.B(n_1574),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1626),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1613),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1610),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1628),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1573),
.Y(n_1667)
);

BUFx4f_ASAP7_75t_SL g1668 ( 
.A(n_1597),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1582),
.B(n_1535),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1581),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1623),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1577),
.B(n_1529),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1570),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1570),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1675)
);

INVx8_ASAP7_75t_L g1676 ( 
.A(n_1577),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1594),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1627),
.B(n_1442),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1605),
.B(n_1530),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1612),
.B(n_1594),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1633),
.B(n_1612),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1647),
.A2(n_1592),
.B(n_1497),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1667),
.B(n_1559),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1646),
.B(n_1559),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1606),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1635),
.B(n_1615),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1681),
.B(n_1558),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1568),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1558),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1678),
.B(n_1599),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1659),
.B(n_1600),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1659),
.B(n_1596),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1636),
.A2(n_1591),
.B1(n_1589),
.B2(n_1564),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1651),
.B(n_1575),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1634),
.B(n_1602),
.C(n_1561),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1653),
.A2(n_1470),
.B(n_1587),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1671),
.A2(n_1631),
.B1(n_1478),
.B2(n_1448),
.C(n_1495),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1669),
.A2(n_1593),
.B(n_1561),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1642),
.B(n_1480),
.C(n_1601),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1640),
.B(n_1605),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1656),
.B(n_1631),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1639),
.B(n_1598),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1673),
.A2(n_1598),
.B(n_1608),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1633),
.A2(n_1587),
.B(n_1629),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1644),
.Y(n_1708)
);

OAI221xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1675),
.A2(n_1446),
.B1(n_1498),
.B2(n_1434),
.C(n_1463),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1639),
.B(n_1574),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1654),
.B(n_1534),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1652),
.B(n_1588),
.C(n_1618),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1652),
.B(n_1567),
.C(n_1566),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1654),
.A2(n_1451),
.B1(n_1577),
.B2(n_1472),
.Y(n_1714)
);

AND2x2_ASAP7_75t_SL g1715 ( 
.A(n_1662),
.B(n_1462),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1661),
.B(n_1519),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1675),
.A2(n_1438),
.B1(n_1455),
.B2(n_1471),
.C(n_1452),
.Y(n_1717)
);

AND4x1_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1534),
.C(n_1604),
.D(n_1595),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1661),
.B(n_1566),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1673),
.B(n_1567),
.C(n_1547),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1643),
.A2(n_1459),
.B(n_1551),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1674),
.A2(n_1680),
.B(n_1662),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1644),
.B(n_1553),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1641),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1664),
.B(n_1553),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1685),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1708),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1682),
.B(n_1679),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1682),
.B(n_1643),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1713),
.B(n_1662),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1705),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1684),
.B(n_1700),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1687),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1691),
.B(n_1664),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1692),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.B(n_1650),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1689),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1674),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1701),
.B(n_1650),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1670),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1693),
.B(n_1665),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1688),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1720),
.B(n_1696),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1702),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1697),
.B(n_1680),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1696),
.B(n_1677),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1710),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1677),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1716),
.B(n_1649),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1715),
.B(n_1677),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1637),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1707),
.B(n_1655),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1695),
.B(n_1637),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1712),
.A2(n_1676),
.B1(n_1637),
.B2(n_1672),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1722),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1655),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1722),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1721),
.B(n_1660),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1756),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1756),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1760),
.B(n_1711),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1729),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1759),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1760),
.B(n_1711),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1759),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1729),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1761),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1734),
.B(n_1683),
.C(n_1565),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1742),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1730),
.B(n_1738),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1703),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1727),
.B(n_1706),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1739),
.B(n_1698),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1738),
.B(n_1706),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1736),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1730),
.B(n_1718),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1745),
.B(n_1668),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1733),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1735),
.B(n_1706),
.Y(n_1783)
);

INVxp67_ASAP7_75t_SL g1784 ( 
.A(n_1745),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1761),
.B(n_1660),
.Y(n_1785)
);

AND2x4_ASAP7_75t_L g1786 ( 
.A(n_1748),
.B(n_1660),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1748),
.B(n_1587),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1748),
.B(n_1672),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1733),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1745),
.B(n_1557),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1745),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1759),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1735),
.B(n_1637),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1744),
.B(n_1724),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1748),
.B(n_1672),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1746),
.B(n_1714),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1753),
.B(n_1672),
.Y(n_1797)
);

NAND2x1_ASAP7_75t_L g1798 ( 
.A(n_1732),
.B(n_1724),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1743),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1737),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1743),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1518),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1737),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1726),
.B(n_1676),
.Y(n_1804)
);

OAI211xp5_ASAP7_75t_L g1805 ( 
.A1(n_1784),
.A2(n_1747),
.B(n_1746),
.C(n_1757),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1766),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1774),
.B(n_1755),
.Y(n_1807)
);

NAND2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1787),
.B(n_1732),
.Y(n_1808)
);

OAI211xp5_ASAP7_75t_L g1809 ( 
.A1(n_1791),
.A2(n_1751),
.B(n_1755),
.C(n_1754),
.Y(n_1809)
);

NOR2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1780),
.B(n_1751),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1766),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1812)
);

OR2x6_ASAP7_75t_L g1813 ( 
.A(n_1763),
.B(n_1752),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1765),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1787),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1770),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1773),
.B(n_1741),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1765),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1780),
.B(n_1732),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1781),
.B(n_1732),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1770),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1801),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1801),
.Y(n_1823)
);

AOI32xp33_ASAP7_75t_L g1824 ( 
.A1(n_1796),
.A2(n_1768),
.A3(n_1778),
.B1(n_1777),
.B2(n_1771),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1798),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1799),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1798),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1799),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1772),
.A2(n_1750),
.B1(n_1752),
.B2(n_1758),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1799),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1763),
.A2(n_1750),
.B1(n_1752),
.B2(n_1762),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1764),
.B(n_1750),
.Y(n_1832)
);

NOR2x1p5_ASAP7_75t_SL g1833 ( 
.A(n_1771),
.B(n_1749),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1773),
.B(n_1740),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1776),
.A2(n_1699),
.B1(n_1749),
.B2(n_1676),
.Y(n_1835)
);

O2A1O1Ixp5_ASAP7_75t_R g1836 ( 
.A1(n_1764),
.A2(n_1728),
.B(n_1726),
.C(n_1731),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1776),
.A2(n_1676),
.B1(n_1762),
.B2(n_1614),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1785),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1782),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1806),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1820),
.B(n_1805),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1814),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1815),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1818),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1819),
.B(n_1768),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1811),
.Y(n_1846)
);

INVxp67_ASAP7_75t_SL g1847 ( 
.A(n_1820),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1819),
.B(n_1802),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1810),
.B(n_1802),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1817),
.B(n_1779),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1816),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1808),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1838),
.B(n_1790),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1824),
.B(n_1779),
.Y(n_1854)
);

OR4x1_ASAP7_75t_L g1855 ( 
.A(n_1836),
.B(n_1800),
.C(n_1789),
.D(n_1782),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1807),
.B(n_1786),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1813),
.Y(n_1857)
);

OAI21xp33_ASAP7_75t_SL g1858 ( 
.A1(n_1824),
.A2(n_1771),
.B(n_1797),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1821),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1834),
.B(n_1812),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1813),
.B(n_1804),
.Y(n_1861)
);

NOR2xp67_ASAP7_75t_L g1862 ( 
.A(n_1829),
.B(n_1786),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1809),
.B(n_1786),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.Y(n_1864)
);

AOI21xp33_ASAP7_75t_L g1865 ( 
.A1(n_1841),
.A2(n_1826),
.B(n_1830),
.Y(n_1865)
);

NAND4xp25_ASAP7_75t_SL g1866 ( 
.A(n_1858),
.B(n_1827),
.C(n_1825),
.D(n_1833),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1845),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1854),
.A2(n_1847),
.B1(n_1862),
.B2(n_1863),
.Y(n_1868)
);

NAND2x1_ASAP7_75t_L g1869 ( 
.A(n_1845),
.B(n_1832),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1857),
.A2(n_1823),
.B(n_1822),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1842),
.Y(n_1871)
);

OAI32xp33_ASAP7_75t_L g1872 ( 
.A1(n_1860),
.A2(n_1831),
.A3(n_1783),
.B1(n_1828),
.B2(n_1793),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1842),
.Y(n_1873)
);

AOI31xp33_ASAP7_75t_L g1874 ( 
.A1(n_1843),
.A2(n_1800),
.A3(n_1789),
.B(n_1803),
.Y(n_1874)
);

OAI22x1_ASAP7_75t_L g1875 ( 
.A1(n_1844),
.A2(n_1786),
.B1(n_1785),
.B2(n_1795),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1860),
.B(n_1832),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1848),
.Y(n_1877)
);

AND2x2_ASAP7_75t_SL g1878 ( 
.A(n_1844),
.B(n_1795),
.Y(n_1878)
);

OAI31xp33_ASAP7_75t_SL g1879 ( 
.A1(n_1849),
.A2(n_1835),
.A3(n_1837),
.B(n_1767),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1840),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1855),
.A2(n_1767),
.B1(n_1792),
.B2(n_1769),
.C(n_1783),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1852),
.A2(n_1832),
.B1(n_1813),
.B2(n_1775),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1840),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1867),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1871),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1877),
.B(n_1848),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_L g1887 ( 
.A(n_1865),
.B(n_1852),
.C(n_1846),
.Y(n_1887)
);

INVx4_ASAP7_75t_L g1888 ( 
.A(n_1873),
.Y(n_1888)
);

O2A1O1Ixp33_ASAP7_75t_SL g1889 ( 
.A1(n_1869),
.A2(n_1864),
.B(n_1846),
.C(n_1859),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1878),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1874),
.B(n_1850),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1850),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1868),
.A2(n_1856),
.B1(n_1861),
.B2(n_1849),
.Y(n_1893)
);

OAI221xp5_ASAP7_75t_L g1894 ( 
.A1(n_1879),
.A2(n_1793),
.B1(n_1861),
.B2(n_1769),
.C(n_1792),
.Y(n_1894)
);

NOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1888),
.B(n_1866),
.Y(n_1895)
);

AOI221x1_ASAP7_75t_SL g1896 ( 
.A1(n_1892),
.A2(n_1876),
.B1(n_1880),
.B2(n_1883),
.C(n_1882),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1891),
.A2(n_1881),
.B1(n_1853),
.B2(n_1870),
.Y(n_1897)
);

AOI321xp33_ASAP7_75t_L g1898 ( 
.A1(n_1894),
.A2(n_1872),
.A3(n_1879),
.B1(n_1859),
.B2(n_1851),
.C(n_1864),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1890),
.A2(n_1853),
.B1(n_1875),
.B2(n_1785),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1888),
.B(n_1851),
.Y(n_1900)
);

NOR3xp33_ASAP7_75t_L g1901 ( 
.A(n_1887),
.B(n_1885),
.C(n_1893),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1884),
.A2(n_1855),
.B1(n_1803),
.B2(n_1785),
.C1(n_1788),
.C2(n_1797),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1886),
.A2(n_1788),
.B1(n_1775),
.B2(n_1794),
.Y(n_1903)
);

AOI21xp33_ASAP7_75t_L g1904 ( 
.A1(n_1889),
.A2(n_1794),
.B(n_1481),
.Y(n_1904)
);

NOR2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1900),
.B(n_1804),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1895),
.B(n_1728),
.Y(n_1906)
);

OA22x2_ASAP7_75t_L g1907 ( 
.A1(n_1899),
.A2(n_1731),
.B1(n_1468),
.B2(n_1555),
.Y(n_1907)
);

OA22x2_ASAP7_75t_L g1908 ( 
.A1(n_1897),
.A2(n_1560),
.B1(n_1630),
.B2(n_1529),
.Y(n_1908)
);

AOI211x1_ASAP7_75t_L g1909 ( 
.A1(n_1896),
.A2(n_1709),
.B(n_1542),
.C(n_1524),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1898),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1901),
.Y(n_1911)
);

NOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1902),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_L g1913 ( 
.A(n_1910),
.B(n_1904),
.C(n_1903),
.Y(n_1913)
);

NAND3xp33_ASAP7_75t_L g1914 ( 
.A(n_1909),
.B(n_1717),
.C(n_1457),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1905),
.B(n_1641),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1906),
.B(n_1666),
.C(n_1663),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1443),
.C(n_1560),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1912),
.B(n_1908),
.Y(n_1918)
);

OA22x2_ASAP7_75t_L g1919 ( 
.A1(n_1915),
.A2(n_1560),
.B1(n_1630),
.B2(n_1666),
.Y(n_1919)
);

NOR3x2_ASAP7_75t_L g1920 ( 
.A(n_1913),
.B(n_1914),
.C(n_1917),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1916),
.A2(n_1630),
.B(n_1530),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1912),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1922),
.B(n_1454),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1918),
.A2(n_1454),
.B1(n_1543),
.B2(n_1537),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1920),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1925),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1926),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1924),
.B1(n_1923),
.B2(n_1919),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1927),
.B(n_1921),
.Y(n_1929)
);

OR4x2_ASAP7_75t_L g1930 ( 
.A(n_1928),
.B(n_1537),
.C(n_1543),
.D(n_1454),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1929),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1931),
.B(n_1663),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_SL g1933 ( 
.A1(n_1930),
.A2(n_1543),
.B1(n_1537),
.B2(n_1454),
.Y(n_1933)
);

AOI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1932),
.A2(n_1464),
.B(n_1437),
.C(n_1658),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1934),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1935),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1936),
.B(n_1933),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1937),
.A2(n_1537),
.B1(n_1543),
.B2(n_1648),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1938),
.A2(n_1648),
.B1(n_1657),
.B2(n_1658),
.Y(n_1939)
);

AOI211xp5_ASAP7_75t_L g1940 ( 
.A1(n_1939),
.A2(n_1464),
.B(n_1657),
.C(n_1616),
.Y(n_1940)
);


endmodule