module fake_jpeg_31961_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_63),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_64),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_48),
.B1(n_52),
.B2(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_46),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_49),
.Y(n_72)
);

AO21x2_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_43),
.B(n_48),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_56),
.B(n_54),
.Y(n_79)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_48),
.B1(n_47),
.B2(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_82),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_87),
.B(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_45),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_0),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_86),
.C(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_21),
.B1(n_35),
.B2(n_34),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_18),
.C(n_33),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_71),
.B(n_69),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_90),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_19),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_1),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_22),
.B(n_32),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_101),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_3),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_4),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_24),
.C(n_31),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_5),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_114),
.B(n_91),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_25),
.B(n_27),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_93),
.Y(n_119)
);

FAx1_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_124),
.CI(n_109),
.CON(n_126),
.SN(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_117),
.C(n_112),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_122),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_120),
.B(n_119),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_129),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_113),
.C(n_118),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_115),
.B(n_116),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_111),
.Y(n_135)
);


endmodule