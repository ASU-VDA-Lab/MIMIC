module fake_jpeg_9330_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_28),
.B1(n_16),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_55),
.B1(n_68),
.B2(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_28),
.B1(n_16),
.B2(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_37),
.B1(n_19),
.B2(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_67),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_25),
.B1(n_35),
.B2(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_37),
.B1(n_19),
.B2(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_40),
.B1(n_18),
.B2(n_20),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_80),
.B(n_71),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_17),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_37),
.B1(n_34),
.B2(n_20),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_60),
.B1(n_90),
.B2(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_89),
.Y(n_104)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

OAI22x1_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_87),
.B1(n_80),
.B2(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_69),
.B1(n_70),
.B2(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_77),
.B1(n_67),
.B2(n_84),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_63),
.C(n_65),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_105),
.C(n_119),
.Y(n_120)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_116),
.B1(n_77),
.B2(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_46),
.B1(n_50),
.B2(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_89),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_93),
.B1(n_82),
.B2(n_50),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_56),
.Y(n_137)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_94),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_65),
.C(n_62),
.Y(n_119)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_122),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_17),
.B(n_33),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_74),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_123),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_130),
.B1(n_134),
.B2(n_119),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_96),
.B1(n_118),
.B2(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_137),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_82),
.C(n_65),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_111),
.C(n_114),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_139),
.B1(n_143),
.B2(n_46),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_113),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_113),
.B1(n_110),
.B2(n_47),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_115),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_46),
.B1(n_50),
.B2(n_47),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_100),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_155),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_154),
.B1(n_139),
.B2(n_141),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_106),
.B1(n_111),
.B2(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_120),
.C(n_133),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_108),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_12),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_1),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_166),
.B(n_169),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_14),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_52),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_66),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_172),
.B(n_17),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_121),
.B1(n_140),
.B2(n_66),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_1),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_130),
.B1(n_128),
.B2(n_135),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_173),
.A2(n_180),
.B1(n_186),
.B2(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_183),
.B1(n_184),
.B2(n_152),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_188),
.C(n_191),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_140),
.B1(n_138),
.B2(n_125),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_140),
.B1(n_121),
.B2(n_32),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_22),
.B1(n_122),
.B2(n_33),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_192),
.B(n_169),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_122),
.C(n_41),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_41),
.C(n_17),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_170),
.B(n_147),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_41),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_161),
.C(n_155),
.Y(n_214)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_202),
.B1(n_206),
.B2(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_208),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_195),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_214),
.C(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_180),
.B1(n_185),
.B2(n_182),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_166),
.C(n_146),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_146),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_213),
.B(n_215),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_167),
.C(n_159),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

XNOR2x2_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_165),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_194),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_172),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_188),
.C(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_185),
.A2(n_172),
.B1(n_33),
.B2(n_32),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_201),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_229),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_178),
.B1(n_174),
.B2(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_220),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_8),
.B(n_14),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_195),
.C(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_233),
.C(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_33),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_32),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_203),
.C(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_237),
.C(n_240),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_198),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_22),
.C(n_31),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_239),
.A2(n_207),
.B1(n_210),
.B2(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_256),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_252),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_255),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_10),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_10),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_253),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_22),
.CI(n_31),
.CON(n_252),
.SN(n_252)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_31),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_19),
.C(n_2),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_256),
.C(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_9),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_243),
.A2(n_238),
.B1(n_237),
.B2(n_224),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_7),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_233),
.B1(n_223),
.B2(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_265),
.B1(n_254),
.B2(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_249),
.B1(n_242),
.B2(n_245),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_268),
.C(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_223),
.C(n_10),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_265),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_252),
.B(n_8),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_271),
.A3(n_277),
.B1(n_272),
.B2(n_280),
.C1(n_275),
.C2(n_270),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_269),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_1),
.C(n_2),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_259),
.B1(n_261),
.B2(n_268),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_6),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_279),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

AOI211xp5_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_260),
.B(n_5),
.C(n_11),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_288),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_5),
.B1(n_12),
.B2(n_15),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_12),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.C(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_15),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_15),
.B(n_2),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_287),
.B(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_3),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_290),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_297),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_300),
.Y(n_304)
);


endmodule