module real_jpeg_6402_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_1),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_1),
.Y(n_401)
);

BUFx5_ASAP7_75t_L g443 ( 
.A(n_1),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_2),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_2),
.A2(n_103),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_2),
.A2(n_103),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_2),
.A2(n_103),
.B1(n_147),
.B2(n_330),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_230),
.B1(n_234),
.B2(n_236),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_248),
.C(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_3),
.B(n_134),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_3),
.B(n_175),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_79),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_3),
.B(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_4),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_5),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_5),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_49),
.B1(n_148),
.B2(n_178),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_5),
.A2(n_113),
.B1(n_114),
.B2(n_148),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_5),
.A2(n_148),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_7),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_8),
.A2(n_45),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_8),
.A2(n_45),
.B1(n_269),
.B2(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_9),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_9),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_72),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_72),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_37),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_13),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_13),
.A2(n_85),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_13),
.A2(n_85),
.B1(n_335),
.B2(n_339),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_13),
.A2(n_55),
.B1(n_76),
.B2(n_85),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_14),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_14),
.A2(n_191),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_14),
.A2(n_191),
.B1(n_230),
.B2(n_317),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_14),
.A2(n_151),
.B1(n_191),
.B2(n_419),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_15),
.A2(n_49),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_15),
.A2(n_277),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_15),
.A2(n_277),
.B1(n_364),
.B2(n_365),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_15),
.A2(n_277),
.B1(n_442),
.B2(n_444),
.Y(n_441)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_220),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_218),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_194),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_20),
.B(n_194),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_121),
.C(n_163),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_21),
.A2(n_22),
.B1(n_121),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_23),
.A2(n_24),
.B(n_82),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_24),
.A2(n_81),
.B1(n_82),
.B2(n_120),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_24),
.A2(n_43),
.B1(n_120),
.B2(n_430),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_36),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_25),
.A2(n_36),
.B1(n_166),
.B2(n_173),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_25),
.A2(n_258),
.B(n_265),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_25),
.A2(n_236),
.B(n_265),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_25),
.A2(n_174),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_26),
.B(n_268),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_26),
.A2(n_266),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_26),
.A2(n_334),
.B1(n_371),
.B2(n_377),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_26),
.A2(n_406),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_29),
.Y(n_378)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_29),
.Y(n_438)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_33),
.Y(n_172)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_41),
.Y(n_264)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_43),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_52),
.B1(n_71),
.B2(n_79),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_44),
.A2(n_52),
.B1(n_79),
.B2(n_177),
.Y(n_176)
);

AO22x2_ASAP7_75t_L g134 ( 
.A1(n_46),
.A2(n_135),
.B1(n_138),
.B2(n_141),
.Y(n_134)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_48),
.Y(n_140)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_48),
.Y(n_346)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_51),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_52),
.A2(n_71),
.B1(n_79),
.B2(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_52),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_52),
.B(n_238),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_62),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_57),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_62),
.A2(n_276),
.B(n_280),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_67),
.Y(n_255)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_67),
.Y(n_338)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_78),
.Y(n_235)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_79),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_101),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_84),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g414 ( 
.A1(n_86),
.A2(n_236),
.B(n_397),
.Y(n_414)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_90),
.B(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_91),
.B(n_236),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_91),
.A2(n_187),
.B1(n_188),
.B2(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_91)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_92),
.Y(n_391)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g330 ( 
.A(n_94),
.Y(n_330)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_96),
.Y(n_365)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_97),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_97),
.Y(n_396)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_101),
.A2(n_200),
.B(n_441),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_108),
.Y(n_101)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_108),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_108),
.A2(n_414),
.B(n_415),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_119),
.Y(n_393)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_121),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_155),
.B(n_162),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_134),
.B1(n_143),
.B2(n_149),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_124),
.A2(n_322),
.B(n_328),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_124),
.B(n_367),
.Y(n_366)
);

AOI22x1_ASAP7_75t_L g447 ( 
.A1(n_124),
.A2(n_134),
.B1(n_367),
.B2(n_448),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_124),
.A2(n_328),
.B(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_125),
.A2(n_144),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_125),
.A2(n_185),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_125),
.A2(n_185),
.B1(n_363),
.B2(n_418),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_128),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_131),
.Y(n_352)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_140),
.Y(n_319)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g345 ( 
.A1(n_146),
.A2(n_325),
.A3(n_346),
.B1(n_347),
.B2(n_350),
.Y(n_345)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_153),
.Y(n_419)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_195),
.CI(n_196),
.CON(n_194),
.SN(n_194)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_163),
.B(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_180),
.C(n_186),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_164),
.B(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_176),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_165),
.B(n_176),
.Y(n_458)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_166),
.Y(n_436)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_171),
.Y(n_295)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_177),
.Y(n_434)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_180),
.B(n_186),
.Y(n_428)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_181),
.Y(n_448)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_185),
.B(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_185),
.A2(n_363),
.B(n_366),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B(n_193),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_193),
.Y(n_415)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_194),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_217),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_216),
.Y(n_202)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_229),
.B(n_237),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_204),
.A2(n_205),
.B1(n_276),
.B2(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_204),
.A2(n_237),
.B(n_316),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_204),
.A2(n_205),
.B1(n_421),
.B2(n_434),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_205),
.A2(n_280),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI311xp33_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_424),
.A3(n_466),
.B1(n_484),
.C1(n_485),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_381),
.B(n_423),
.Y(n_222)
);

AO21x1_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_354),
.B(n_380),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_310),
.B(n_353),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_283),
.B(n_309),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_256),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_227),
.B(n_256),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_242),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_228),
.A2(n_242),
.B1(n_243),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

INVx5_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_236),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_236),
.B(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_273),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_274),
.C(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_258),
.Y(n_305)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_271),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_281),
.B2(n_282),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g350 ( 
.A(n_278),
.B(n_351),
.Y(n_350)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_302),
.B(n_308),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_292),
.B(n_301),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_289),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_300),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_298),
.B(n_299),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_333),
.B(n_342),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_306),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_312),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_331),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_320),
.B2(n_321),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_320),
.C(n_331),
.Y(n_355)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_345),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_345),
.Y(n_360)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx4_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_355),
.B(n_356),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_361),
.B2(n_379),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_360),
.C(n_379),
.Y(n_382)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_368),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_362),
.B(n_369),
.C(n_370),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g387 ( 
.A1(n_365),
.A2(n_388),
.A3(n_390),
.B1(n_392),
.B2(n_397),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_382),
.B(n_383),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_411),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.Y(n_384)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_402),
.B2(n_403),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_402),
.Y(n_462)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

INVx6_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_408),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_408),
.B(n_409),
.C(n_411),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_416),
.B2(n_422),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_412),
.B(n_417),
.C(n_420),
.Y(n_475)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_416),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_452),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_SL g485 ( 
.A1(n_425),
.A2(n_452),
.B(n_486),
.C(n_489),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_449),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_449),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.C(n_431),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g465 ( 
.A(n_427),
.B(n_429),
.CI(n_431),
.CON(n_465),
.SN(n_465)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_447),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_435),
.Y(n_474)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_439),
.A2(n_440),
.B1(n_447),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_465),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_465),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.C(n_459),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.C(n_463),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_460),
.A2(n_461),
.B1(n_463),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_463),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g491 ( 
.A(n_465),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_479),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_468),
.A2(n_487),
.B(n_488),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_476),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_476),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.C(n_475),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_482),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_474),
.B1(n_475),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_481),
.Y(n_487)
);


endmodule