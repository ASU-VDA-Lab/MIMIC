module real_aes_7431_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g480 ( .A1(n_0), .A2(n_163), .B(n_481), .C(n_484), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_1), .B(n_475), .Y(n_486) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_2), .B(n_91), .C(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
INVx1_ASAP7_75t_L g201 ( .A(n_3), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_4), .B(n_164), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g141 ( .A1(n_5), .A2(n_142), .B1(n_143), .B2(n_449), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_5), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_5), .A2(n_98), .B1(n_449), .B2(n_749), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_6), .A2(n_460), .B(n_507), .Y(n_506) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_7), .A2(n_170), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_8), .A2(n_39), .B1(n_167), .B2(n_219), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_9), .B(n_170), .Y(n_187) );
AND2x6_ASAP7_75t_L g172 ( .A(n_10), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_11), .A2(n_172), .B(n_463), .C(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_12), .B(n_40), .Y(n_109) );
INVx1_ASAP7_75t_L g154 ( .A(n_13), .Y(n_154) );
INVx1_ASAP7_75t_L g193 ( .A(n_14), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_15), .B(n_160), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_16), .A2(n_42), .B1(n_535), .B2(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_16), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_17), .B(n_164), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_18), .B(n_150), .Y(n_149) );
AO32x2_ASAP7_75t_L g230 ( .A1(n_19), .A2(n_170), .A3(n_171), .B1(n_190), .B2(n_231), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_20), .A2(n_106), .B1(n_115), .B2(n_756), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_21), .B(n_167), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_22), .B(n_150), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_23), .A2(n_55), .B1(n_167), .B2(n_219), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g227 ( .A1(n_24), .A2(n_83), .B1(n_160), .B2(n_167), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_25), .B(n_167), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_26), .A2(n_171), .B(n_463), .C(n_465), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_27), .A2(n_171), .B(n_463), .C(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_28), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_29), .A2(n_99), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_29), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_30), .B(n_209), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_31), .A2(n_460), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_32), .B(n_209), .Y(n_246) );
INVx2_ASAP7_75t_L g162 ( .A(n_33), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_34), .A2(n_495), .B(n_496), .C(n_500), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_35), .B(n_167), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_36), .B(n_209), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_37), .A2(n_134), .B1(n_137), .B2(n_138), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_37), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_38), .B(n_215), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_41), .B(n_459), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_42), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_43), .B(n_164), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_44), .B(n_460), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_45), .A2(n_495), .B(n_500), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_46), .B(n_167), .Y(n_180) );
INVx1_ASAP7_75t_L g482 ( .A(n_47), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_48), .A2(n_751), .B1(n_752), .B2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g754 ( .A(n_48), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_49), .A2(n_92), .B1(n_219), .B2(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g521 ( .A(n_50), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_51), .B(n_167), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_52), .B(n_167), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_53), .B(n_460), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_54), .B(n_185), .Y(n_184) );
AOI22xp33_ASAP7_75t_SL g166 ( .A1(n_56), .A2(n_61), .B1(n_160), .B2(n_167), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_57), .A2(n_131), .B1(n_132), .B2(n_133), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_57), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_58), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_59), .B(n_167), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_60), .B(n_167), .Y(n_266) );
INVx1_ASAP7_75t_L g173 ( .A(n_62), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_63), .B(n_460), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_64), .B(n_475), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_65), .A2(n_185), .B(n_196), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_66), .B(n_167), .Y(n_202) );
INVx1_ASAP7_75t_L g153 ( .A(n_67), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_69), .B(n_164), .Y(n_498) );
AO32x2_ASAP7_75t_L g223 ( .A1(n_70), .A2(n_170), .A3(n_171), .B1(n_224), .B2(n_228), .Y(n_223) );
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_71), .A2(n_129), .B1(n_130), .B2(n_139), .C1(n_734), .C2(n_740), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_72), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_73), .B(n_165), .Y(n_532) );
INVx1_ASAP7_75t_L g265 ( .A(n_74), .Y(n_265) );
INVx1_ASAP7_75t_L g241 ( .A(n_75), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_76), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_77), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_78), .A2(n_463), .B(n_500), .C(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_79), .B(n_160), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g508 ( .A(n_80), .Y(n_508) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_82), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_84), .B(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_85), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_86), .B(n_160), .Y(n_245) );
INVx2_ASAP7_75t_L g151 ( .A(n_87), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_88), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_89), .B(n_157), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_90), .B(n_160), .Y(n_181) );
OR2x2_ASAP7_75t_L g123 ( .A(n_91), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g450 ( .A(n_91), .B(n_125), .Y(n_450) );
INVx2_ASAP7_75t_L g733 ( .A(n_91), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_93), .A2(n_104), .B1(n_160), .B2(n_161), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_94), .B(n_460), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_95), .Y(n_497) );
INVxp67_ASAP7_75t_L g511 ( .A(n_96), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_97), .B(n_160), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_98), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_99), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g528 ( .A(n_101), .Y(n_528) );
INVx1_ASAP7_75t_L g557 ( .A(n_102), .Y(n_557) );
AND2x2_ASAP7_75t_L g523 ( .A(n_103), .B(n_209), .Y(n_523) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_108), .Y(n_756) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g125 ( .A(n_109), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_128), .B1(n_743), .B2(n_744), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g743 ( .A(n_118), .Y(n_743) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_120), .A2(n_745), .B(n_755), .Y(n_744) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_127), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_123), .Y(n_755) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_124), .B(n_733), .Y(n_742) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g732 ( .A(n_125), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_134), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_450), .B1(n_451), .B2(n_732), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_141), .A2(n_735), .B1(n_737), .B2(n_738), .Y(n_734) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
XNOR2xp5_ASAP7_75t_L g747 ( .A(n_143), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_383), .Y(n_143) );
NOR5xp2_ASAP7_75t_L g144 ( .A(n_145), .B(n_296), .C(n_342), .D(n_355), .E(n_367), .Y(n_144) );
OAI211xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_204), .B(n_250), .C(n_277), .Y(n_145) );
INVx1_ASAP7_75t_SL g378 ( .A(n_146), .Y(n_378) );
OR2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_174), .Y(n_146) );
AND2x2_ASAP7_75t_L g302 ( .A(n_147), .B(n_175), .Y(n_302) );
AND2x2_ASAP7_75t_L g330 ( .A(n_147), .B(n_276), .Y(n_330) );
AND2x2_ASAP7_75t_L g338 ( .A(n_147), .B(n_281), .Y(n_338) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g268 ( .A(n_148), .B(n_176), .Y(n_268) );
INVx2_ASAP7_75t_L g280 ( .A(n_148), .Y(n_280) );
AND2x2_ASAP7_75t_L g405 ( .A(n_148), .B(n_347), .Y(n_405) );
OR2x2_ASAP7_75t_L g407 ( .A(n_148), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_155), .Y(n_148) );
INVx1_ASAP7_75t_L g274 ( .A(n_149), .Y(n_274) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx1_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_151), .B(n_152), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NAND3xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_169), .C(n_171), .Y(n_155) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_156), .A2(n_169), .B(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B1(n_163), .B2(n_166), .Y(n_156) );
INVx2_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
OAI22xp5_ASAP7_75t_SL g224 ( .A1(n_157), .A2(n_165), .B1(n_225), .B2(n_227), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_157), .A2(n_163), .B1(n_232), .B2(n_233), .Y(n_231) );
INVx4_ASAP7_75t_L g483 ( .A(n_157), .Y(n_483) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
INVx1_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
AND2x2_ASAP7_75t_L g461 ( .A(n_158), .B(n_186), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_158), .Y(n_464) );
INVx2_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g168 ( .A(n_162), .Y(n_168) );
INVx1_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_163), .A2(n_183), .B(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_164), .A2(n_180), .B(n_181), .Y(n_179) );
O2A1O1Ixp5_ASAP7_75t_SL g239 ( .A1(n_164), .A2(n_240), .B(n_241), .C(n_242), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_164), .A2(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_164), .B(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_167), .Y(n_559) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
BUFx3_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
AND2x6_ASAP7_75t_L g463 ( .A(n_168), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g475 ( .A(n_169), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_169), .B(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_169), .A2(n_527), .B(n_534), .Y(n_526) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_169), .A2(n_554), .B(n_561), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_169), .B(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_170), .A2(n_178), .B(n_187), .Y(n_177) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_170), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_170), .A2(n_539), .B(n_540), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_171), .A2(n_261), .B(n_264), .Y(n_260) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_179), .B(n_182), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_192), .B(n_199), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_172), .A2(n_211), .B(n_216), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_172), .A2(n_239), .B(n_243), .Y(n_238) );
AND2x4_ASAP7_75t_L g460 ( .A(n_172), .B(n_461), .Y(n_460) );
INVx4_ASAP7_75t_SL g485 ( .A(n_172), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_172), .B(n_461), .Y(n_529) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g318 ( .A(n_175), .B(n_290), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_175), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g432 ( .A(n_175), .B(n_272), .Y(n_432) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_188), .Y(n_175) );
AND2x2_ASAP7_75t_L g275 ( .A(n_176), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g322 ( .A(n_176), .Y(n_322) );
AND2x2_ASAP7_75t_L g347 ( .A(n_176), .B(n_259), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_176), .B(n_380), .Y(n_417) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g281 ( .A(n_177), .B(n_259), .Y(n_281) );
AND2x2_ASAP7_75t_L g295 ( .A(n_177), .B(n_258), .Y(n_295) );
AND2x2_ASAP7_75t_L g312 ( .A(n_177), .B(n_188), .Y(n_312) );
AND2x2_ASAP7_75t_L g369 ( .A(n_177), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_177), .B(n_276), .Y(n_382) );
AND2x2_ASAP7_75t_L g434 ( .A(n_177), .B(n_359), .Y(n_434) );
INVx2_ASAP7_75t_L g200 ( .A(n_185), .Y(n_200) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g257 ( .A(n_188), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g276 ( .A(n_188), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_188), .B(n_259), .Y(n_353) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_191), .B(n_203), .Y(n_188) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_189), .A2(n_260), .B(n_267), .Y(n_259) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_190), .B(n_535), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_196), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_194), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_194), .A2(n_542), .B(n_543), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_196), .A2(n_557), .B(n_558), .C(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_197), .A2(n_244), .B(n_245), .Y(n_243) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g467 ( .A(n_198), .Y(n_467) );
O2A1O1Ixp5_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_220), .B(n_265), .C(n_266), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_200), .A2(n_466), .B(n_468), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_234), .B(n_247), .Y(n_204) );
INVx1_ASAP7_75t_SL g366 ( .A(n_205), .Y(n_366) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_222), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_207), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g249 ( .A(n_208), .Y(n_249) );
INVx1_ASAP7_75t_L g286 ( .A(n_208), .Y(n_286) );
AND2x2_ASAP7_75t_L g307 ( .A(n_208), .B(n_229), .Y(n_307) );
AND2x2_ASAP7_75t_L g341 ( .A(n_208), .B(n_230), .Y(n_341) );
OR2x2_ASAP7_75t_L g360 ( .A(n_208), .B(n_236), .Y(n_360) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_208), .Y(n_374) );
AND2x2_ASAP7_75t_L g387 ( .A(n_208), .B(n_388), .Y(n_387) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_221), .Y(n_208) );
INVx2_ASAP7_75t_L g228 ( .A(n_209), .Y(n_228) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_209), .A2(n_238), .B(n_246), .Y(n_237) );
INVx1_ASAP7_75t_L g473 ( .A(n_209), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_209), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_209), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_220), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_222), .A2(n_309), .B1(n_310), .B2(n_319), .Y(n_308) );
AND2x2_ASAP7_75t_L g392 ( .A(n_222), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
INVx1_ASAP7_75t_L g253 ( .A(n_223), .Y(n_253) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_223), .Y(n_290) );
INVx1_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
AND2x2_ASAP7_75t_L g316 ( .A(n_223), .B(n_230), .Y(n_316) );
INVx2_ASAP7_75t_L g484 ( .A(n_226), .Y(n_484) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_226), .Y(n_499) );
INVx1_ASAP7_75t_L g470 ( .A(n_228), .Y(n_470) );
OR2x2_ASAP7_75t_L g270 ( .A(n_229), .B(n_255), .Y(n_270) );
AND2x2_ASAP7_75t_L g300 ( .A(n_229), .B(n_301), .Y(n_300) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_229), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g248 ( .A(n_230), .B(n_249), .Y(n_248) );
BUFx2_ASAP7_75t_L g357 ( .A(n_230), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_234), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g335 ( .A(n_235), .B(n_301), .Y(n_335) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g247 ( .A(n_236), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g255 ( .A(n_237), .Y(n_255) );
OR2x2_ASAP7_75t_L g285 ( .A(n_237), .B(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_237), .Y(n_340) );
AOI32xp33_ASAP7_75t_L g377 ( .A1(n_247), .A2(n_307), .A3(n_378), .B1(n_379), .B2(n_381), .Y(n_377) );
AND2x2_ASAP7_75t_L g303 ( .A(n_248), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_248), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_248), .B(n_335), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_248), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_256), .B1(n_269), .B2(n_271), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g356 ( .A(n_252), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_253), .B(n_255), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_254), .A2(n_278), .B1(n_282), .B2(n_292), .Y(n_277) );
AND2x2_ASAP7_75t_L g299 ( .A(n_254), .B(n_300), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_254), .A2(n_268), .B(n_316), .C(n_351), .Y(n_350) );
OAI332xp33_ASAP7_75t_L g355 ( .A1(n_254), .A2(n_356), .A3(n_358), .B1(n_360), .B2(n_361), .B3(n_363), .C1(n_364), .C2(n_366), .Y(n_355) );
INVx2_ASAP7_75t_L g396 ( .A(n_254), .Y(n_396) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_255), .Y(n_314) );
INVx1_ASAP7_75t_L g389 ( .A(n_255), .Y(n_389) );
AND2x2_ASAP7_75t_L g443 ( .A(n_255), .B(n_307), .Y(n_443) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_268), .Y(n_256) );
AND2x2_ASAP7_75t_L g323 ( .A(n_258), .B(n_273), .Y(n_323) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g371 ( .A(n_259), .B(n_273), .Y(n_371) );
INVx1_ASAP7_75t_L g380 ( .A(n_259), .Y(n_380) );
INVx1_ASAP7_75t_L g354 ( .A(n_268), .Y(n_354) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g438 ( .A(n_270), .B(n_290), .Y(n_438) );
INVx1_ASAP7_75t_SL g349 ( .A(n_271), .Y(n_349) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
AND2x2_ASAP7_75t_L g376 ( .A(n_272), .B(n_334), .Y(n_376) );
INVx1_ASAP7_75t_L g395 ( .A(n_272), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_272), .B(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
AND2x2_ASAP7_75t_L g298 ( .A(n_275), .B(n_279), .Y(n_298) );
AND2x2_ASAP7_75t_L g365 ( .A(n_275), .B(n_323), .Y(n_365) );
INVx2_ASAP7_75t_L g408 ( .A(n_275), .Y(n_408) );
INVx2_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_276), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g309 ( .A(n_279), .Y(n_309) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_280), .B(n_353), .Y(n_359) );
OR2x2_ASAP7_75t_L g423 ( .A(n_280), .B(n_382), .Y(n_423) );
INVx1_ASAP7_75t_L g447 ( .A(n_280), .Y(n_447) );
INVx1_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
AND2x2_ASAP7_75t_L g448 ( .A(n_281), .B(n_291), .Y(n_448) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_285), .A2(n_311), .B1(n_313), .B2(n_317), .Y(n_310) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI322xp33_ASAP7_75t_SL g394 ( .A1(n_288), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_398), .C1(n_401), .C2(n_403), .Y(n_394) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g391 ( .A(n_289), .B(n_307), .Y(n_391) );
OR2x2_ASAP7_75t_L g425 ( .A(n_289), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g428 ( .A(n_289), .B(n_360), .Y(n_428) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g373 ( .A(n_290), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g429 ( .A(n_290), .B(n_360), .Y(n_429) );
INVx3_ASAP7_75t_L g362 ( .A(n_291), .Y(n_362) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g418 ( .A(n_293), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g297 ( .A1(n_295), .A2(n_298), .B1(n_299), .B2(n_302), .C1(n_303), .C2(n_305), .Y(n_297) );
INVx1_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
NAND3xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_308), .C(n_325), .Y(n_296) );
AND2x2_ASAP7_75t_L g413 ( .A(n_300), .B(n_314), .Y(n_413) );
BUFx2_ASAP7_75t_L g304 ( .A(n_301), .Y(n_304) );
INVx1_ASAP7_75t_L g345 ( .A(n_301), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_302), .A2(n_338), .B1(n_391), .B2(n_392), .C(n_394), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_304), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_307), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_307), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_312), .B(n_323), .Y(n_324) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_314), .A2(n_320), .B(n_324), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_314), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g411 ( .A(n_316), .B(n_393), .Y(n_411) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g334 ( .A(n_322), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_323), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_331), .B1(n_332), .B2(n_335), .C(n_336), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_327), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g436 ( .A(n_335), .B(n_341), .Y(n_436) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
OAI31xp33_ASAP7_75t_SL g404 ( .A1(n_339), .A2(n_378), .A3(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g393 ( .A(n_340), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_341), .B(n_345), .Y(n_444) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_346), .B1(n_348), .B2(n_349), .C(n_350), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_344), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_347), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g363 ( .A(n_356), .Y(n_363) );
INVx2_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g385 ( .A(n_362), .B(n_371), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_362), .A2(n_379), .B(n_436), .C(n_437), .Y(n_435) );
OAI221xp5_ASAP7_75t_SL g367 ( .A1(n_363), .A2(n_368), .B1(n_372), .B2(n_375), .C(n_377), .Y(n_367) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_366), .A2(n_431), .B(n_433), .C(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_369), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_427), .Y(n_419) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NOR4xp25_ASAP7_75t_L g383 ( .A(n_384), .B(n_409), .C(n_430), .D(n_441), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .B(n_390), .C(n_404), .Y(n_384) );
INVx1_ASAP7_75t_SL g439 ( .A(n_391), .Y(n_439) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_SL g402 ( .A(n_400), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_407), .A2(n_416), .B1(n_428), .B2(n_429), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_414), .C(n_419), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI31xp33_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_442), .A3(n_444), .B(n_445), .Y(n_441) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g736 ( .A(n_450), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_451), .Y(n_737) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_668), .Y(n_451) );
NOR5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_599), .C(n_628), .D(n_648), .E(n_655), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_487), .B(n_544), .C(n_586), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_455), .A2(n_671), .B1(n_673), .B2(n_674), .Y(n_670) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_474), .Y(n_455) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_456), .Y(n_547) );
AND2x4_ASAP7_75t_L g579 ( .A(n_456), .B(n_580), .Y(n_579) );
INVx5_ASAP7_75t_L g597 ( .A(n_456), .Y(n_597) );
AND2x2_ASAP7_75t_L g606 ( .A(n_456), .B(n_598), .Y(n_606) );
AND2x2_ASAP7_75t_L g618 ( .A(n_456), .B(n_491), .Y(n_618) );
AND2x2_ASAP7_75t_L g714 ( .A(n_456), .B(n_582), .Y(n_714) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_471), .Y(n_456) );
AOI21xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_462), .B(n_470), .Y(n_457) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
INVx2_ASAP7_75t_L g469 ( .A(n_467), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_469), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_469), .A2(n_499), .B(n_521), .C(n_522), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g580 ( .A(n_474), .Y(n_580) );
AND2x2_ASAP7_75t_L g598 ( .A(n_474), .B(n_553), .Y(n_598) );
AND2x2_ASAP7_75t_L g617 ( .A(n_474), .B(n_552), .Y(n_617) );
AND2x2_ASAP7_75t_L g657 ( .A(n_474), .B(n_597), .Y(n_657) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_486), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_479), .B(n_480), .C(n_485), .Y(n_477) );
INVx2_ASAP7_75t_L g495 ( .A(n_479), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_479), .A2(n_485), .B(n_508), .C(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g500 ( .A(n_485), .Y(n_500) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_513), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI322xp5_ASAP7_75t_L g716 ( .A1(n_490), .A2(n_524), .A3(n_571), .B1(n_579), .B2(n_633), .C1(n_717), .C2(n_720), .Y(n_716) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_503), .Y(n_490) );
INVx5_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
AND2x2_ASAP7_75t_L g565 ( .A(n_491), .B(n_551), .Y(n_565) );
BUFx2_ASAP7_75t_L g643 ( .A(n_491), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_491), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g720 ( .A(n_491), .B(n_627), .Y(n_720) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_503), .B(n_515), .Y(n_574) );
INVx1_ASAP7_75t_L g601 ( .A(n_503), .Y(n_601) );
AND2x2_ASAP7_75t_L g614 ( .A(n_503), .B(n_536), .Y(n_614) );
AND2x2_ASAP7_75t_L g715 ( .A(n_503), .B(n_633), .Y(n_715) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g569 ( .A(n_504), .B(n_515), .Y(n_569) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_504), .Y(n_577) );
OR2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_536), .Y(n_584) );
AND2x2_ASAP7_75t_L g594 ( .A(n_504), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_504), .B(n_526), .Y(n_623) );
INVxp67_ASAP7_75t_L g647 ( .A(n_504), .Y(n_647) );
AND2x2_ASAP7_75t_L g654 ( .A(n_504), .B(n_524), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_504), .B(n_536), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_504), .B(n_525), .Y(n_680) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_515), .B(n_537), .Y(n_624) );
OR2x2_ASAP7_75t_L g646 ( .A(n_515), .B(n_525), .Y(n_646) );
AND2x2_ASAP7_75t_L g659 ( .A(n_515), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_515), .B(n_614), .Y(n_665) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_515), .A2(n_670), .B(n_675), .C(n_684), .Y(n_669) );
AND2x2_ASAP7_75t_L g730 ( .A(n_515), .B(n_536), .Y(n_730) );
INVx5_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g583 ( .A(n_516), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_516), .B(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_516), .B(n_578), .Y(n_590) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_516), .Y(n_592) );
OR2x2_ASAP7_75t_L g603 ( .A(n_516), .B(n_525), .Y(n_603) );
AND2x2_ASAP7_75t_SL g608 ( .A(n_516), .B(n_594), .Y(n_608) );
AND2x2_ASAP7_75t_L g633 ( .A(n_516), .B(n_525), .Y(n_633) );
AND2x2_ASAP7_75t_L g653 ( .A(n_516), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g691 ( .A(n_516), .B(n_524), .Y(n_691) );
OR2x2_ASAP7_75t_L g694 ( .A(n_516), .B(n_680), .Y(n_694) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_525), .A2(n_638), .B(n_641), .C(n_647), .Y(n_637) );
INVx5_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_526), .B(n_536), .Y(n_568) );
AND2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_537), .Y(n_572) );
OR2x2_ASAP7_75t_L g578 ( .A(n_526), .B(n_536), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_SL g595 ( .A(n_536), .Y(n_595) );
OR2x2_ASAP7_75t_L g723 ( .A(n_536), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_563), .B(n_566), .C(n_575), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI31xp33_ASAP7_75t_L g648 ( .A1(n_546), .A2(n_649), .A3(n_651), .B(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_547), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_548), .B(n_579), .Y(n_585) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_549), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g605 ( .A(n_549), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_549), .B(n_580), .Y(n_610) );
AND2x2_ASAP7_75t_L g620 ( .A(n_549), .B(n_579), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_549), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g640 ( .A(n_549), .B(n_597), .Y(n_640) );
AND2x2_ASAP7_75t_L g645 ( .A(n_549), .B(n_617), .Y(n_645) );
OR2x2_ASAP7_75t_L g664 ( .A(n_549), .B(n_551), .Y(n_664) );
OR2x2_ASAP7_75t_L g666 ( .A(n_549), .B(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_549), .Y(n_713) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g613 ( .A(n_551), .B(n_580), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_551), .B(n_597), .Y(n_636) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g582 ( .A(n_553), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g673 ( .A(n_565), .B(n_597), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_565), .A2(n_579), .A3(n_617), .B1(n_676), .B2(n_677), .C1(n_678), .C2(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g683 ( .A(n_565), .Y(n_683) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx1_ASAP7_75t_SL g677 ( .A(n_567), .Y(n_677) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g629 ( .A(n_568), .B(n_574), .Y(n_629) );
INVx1_ASAP7_75t_L g660 ( .A(n_568), .Y(n_660) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .A3(n_581), .B1(n_583), .B2(n_585), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_578), .A2(n_593), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g630 ( .A(n_579), .Y(n_630) );
AND2x4_ASAP7_75t_L g627 ( .A(n_580), .B(n_597), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_580), .B(n_663), .Y(n_662) );
AOI322xp5_ASAP7_75t_L g692 ( .A1(n_581), .A2(n_608), .A3(n_627), .B1(n_660), .B2(n_693), .C1(n_695), .C2(n_696), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_581), .A2(n_658), .B1(n_722), .B2(n_723), .C(n_725), .Y(n_721) );
AND2x2_ASAP7_75t_L g609 ( .A(n_582), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g589 ( .A(n_584), .Y(n_589) );
OR2x2_ASAP7_75t_L g661 ( .A(n_584), .B(n_646), .Y(n_661) );
OAI31xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .A3(n_591), .B(n_596), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_587), .A2(n_620), .B1(n_621), .B2(n_625), .Y(n_619) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g632 ( .A(n_589), .B(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_591), .A2(n_632), .B1(n_685), .B2(n_688), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g674 ( .A(n_594), .B(n_643), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_594), .B(n_633), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_595), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g708 ( .A(n_595), .B(n_646), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_596), .A2(n_691), .B1(n_704), .B2(n_707), .Y(n_703) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_L g612 ( .A(n_597), .Y(n_612) );
AND2x2_ASAP7_75t_L g695 ( .A(n_597), .B(n_617), .Y(n_695) );
OR2x2_ASAP7_75t_L g697 ( .A(n_597), .B(n_664), .Y(n_697) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_597), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_598), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_598), .B(n_643), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_604), .B(n_607), .C(n_619), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_611), .B2(n_614), .C(n_615), .Y(n_607) );
INVxp67_ASAP7_75t_L g719 ( .A(n_610), .Y(n_719) );
INVx1_ASAP7_75t_L g686 ( .A(n_611), .Y(n_686) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g650 ( .A(n_612), .B(n_617), .Y(n_650) );
INVx1_ASAP7_75t_L g667 ( .A(n_613), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_613), .B(n_640), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g682 ( .A(n_617), .Y(n_682) );
AND2x2_ASAP7_75t_L g688 ( .A(n_617), .B(n_643), .Y(n_688) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_SL g676 ( .A(n_624), .Y(n_676) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_627), .B(n_663), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_634), .C(n_637), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g724 ( .A(n_633), .Y(n_724) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g642 ( .A(n_636), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_640), .B(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B(n_646), .Y(n_641) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_644), .A2(n_690), .B(n_692), .C(n_698), .Y(n_689) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g701 ( .A(n_646), .Y(n_701) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI222xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B1(n_661), .B2(n_662), .C1(n_665), .C2(n_666), .Y(n_655) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g731 ( .A(n_662), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_663), .B(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_663), .A2(n_710), .B1(n_712), .B2(n_715), .Y(n_709) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g668 ( .A(n_669), .B(n_689), .C(n_702), .D(n_721), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_671), .B(n_701), .Y(n_711) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g678 ( .A(n_676), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_679), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_709), .C(n_716), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_L g718 ( .A(n_714), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_728), .B(n_731), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g739 ( .A(n_732), .Y(n_739) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XOR2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_750), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
endmodule