module real_aes_8439_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_0), .B(n_83), .C(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g452 ( .A(n_1), .Y(n_452) );
INVx1_ASAP7_75t_L g255 ( .A(n_2), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_3), .A2(n_37), .B1(n_205), .B2(n_491), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g216 ( .A1(n_4), .A2(n_138), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_5), .B(n_160), .Y(n_477) );
AND2x6_ASAP7_75t_L g143 ( .A(n_6), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_7), .A2(n_137), .B(n_145), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_8), .B(n_38), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_9), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g222 ( .A(n_10), .Y(n_222) );
INVx1_ASAP7_75t_L g135 ( .A(n_11), .Y(n_135) );
INVx1_ASAP7_75t_L g446 ( .A(n_12), .Y(n_446) );
INVx1_ASAP7_75t_L g155 ( .A(n_13), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_14), .B(n_229), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_15), .A2(n_100), .B1(n_109), .B2(n_726), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_16), .B(n_161), .Y(n_479) );
AO32x2_ASAP7_75t_L g525 ( .A1(n_17), .A2(n_160), .A3(n_176), .B1(n_465), .B2(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_18), .B(n_205), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_19), .B(n_172), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_20), .B(n_161), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_21), .A2(n_49), .B1(n_205), .B2(n_491), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_22), .B(n_138), .Y(n_165) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_23), .A2(n_74), .B1(n_205), .B2(n_229), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_24), .B(n_205), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_25), .B(n_215), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_26), .A2(n_152), .B(n_154), .C(n_156), .Y(n_151) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_27), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_28), .B(n_131), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_29), .B(n_187), .Y(n_256) );
AOI222xp33_ASAP7_75t_SL g121 ( .A1(n_30), .A2(n_88), .B1(n_122), .B2(n_711), .C1(n_712), .C2(n_715), .Y(n_121) );
INVx1_ASAP7_75t_L g711 ( .A(n_30), .Y(n_711) );
INVx1_ASAP7_75t_L g234 ( .A(n_31), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_32), .B(n_131), .Y(n_503) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_34), .B(n_205), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_35), .B(n_131), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_36), .A2(n_143), .B(n_148), .C(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g232 ( .A(n_39), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_40), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_41), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_42), .B(n_205), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_43), .A2(n_84), .B1(n_157), .B2(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_44), .B(n_205), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_45), .B(n_205), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_46), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_47), .B(n_451), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_48), .B(n_138), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_50), .A2(n_59), .B1(n_205), .B2(n_229), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_51), .A2(n_148), .B1(n_229), .B2(n_231), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_52), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_53), .B(n_205), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_54), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_55), .B(n_205), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_56), .A2(n_220), .B(n_221), .C(n_223), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_57), .Y(n_191) );
INVx1_ASAP7_75t_L g218 ( .A(n_58), .Y(n_218) );
INVx1_ASAP7_75t_L g144 ( .A(n_60), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_61), .B(n_205), .Y(n_453) );
INVx1_ASAP7_75t_L g134 ( .A(n_62), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_63), .Y(n_113) );
AO32x2_ASAP7_75t_L g488 ( .A1(n_64), .A2(n_160), .A3(n_197), .B1(n_465), .B2(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g463 ( .A(n_65), .Y(n_463) );
INVx1_ASAP7_75t_L g498 ( .A(n_66), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_SL g242 ( .A1(n_67), .A2(n_172), .B(n_223), .C(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g244 ( .A(n_68), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_69), .B(n_229), .Y(n_499) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_71), .Y(n_237) );
INVx1_ASAP7_75t_L g182 ( .A(n_72), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_73), .A2(n_124), .B1(n_713), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_73), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_75), .A2(n_143), .B(n_148), .C(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_76), .B(n_491), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_77), .B(n_229), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_78), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_80), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_81), .B(n_229), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_82), .A2(n_143), .B(n_148), .C(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g116 ( .A(n_83), .B(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g123 ( .A(n_83), .B(n_118), .Y(n_123) );
INVx2_ASAP7_75t_L g435 ( .A(n_83), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_85), .A2(n_98), .B1(n_229), .B2(n_230), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_86), .B(n_131), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_87), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_89), .A2(n_143), .B(n_148), .C(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_90), .Y(n_208) );
INVx1_ASAP7_75t_L g241 ( .A(n_91), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_92), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_93), .B(n_169), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_94), .B(n_229), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_95), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_97), .A2(n_138), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g726 ( .A(n_102), .Y(n_726) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
AND2x2_ASAP7_75t_L g118 ( .A(n_103), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AOI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_121), .B1(n_718), .B2(n_721), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g720 ( .A(n_113), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_114), .A2(n_722), .B(n_724), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g114 ( .A(n_115), .B(n_120), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g725 ( .A(n_116), .Y(n_725) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_117), .B(n_435), .Y(n_717) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g434 ( .A(n_118), .B(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_432), .B2(n_436), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_123), .A2(n_434), .B1(n_713), .B2(n_714), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_124), .Y(n_713) );
OR4x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_328), .C(n_387), .D(n_414), .Y(n_124) );
NAND3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_270), .C(n_295), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_193), .B(n_213), .C(n_246), .Y(n_126) );
AOI211xp5_ASAP7_75t_SL g418 ( .A1(n_127), .A2(n_419), .B(n_421), .C(n_424), .Y(n_418) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
INVx1_ASAP7_75t_L g293 ( .A(n_128), .Y(n_293) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g268 ( .A(n_129), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g300 ( .A(n_129), .Y(n_300) );
AND2x2_ASAP7_75t_L g355 ( .A(n_129), .B(n_324), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_129), .B(n_211), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_129), .B(n_212), .Y(n_413) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g274 ( .A(n_130), .Y(n_274) );
AND2x2_ASAP7_75t_L g317 ( .A(n_130), .B(n_180), .Y(n_317) );
AND2x2_ASAP7_75t_L g335 ( .A(n_130), .B(n_212), .Y(n_335) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .B(n_159), .Y(n_130) );
INVx1_ASAP7_75t_L g192 ( .A(n_131), .Y(n_192) );
INVx2_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_131), .A2(n_496), .B(n_503), .Y(n_495) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_131), .A2(n_505), .B(n_513), .Y(n_504) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_L g161 ( .A(n_132), .B(n_133), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_139), .B(n_143), .Y(n_183) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g451 ( .A(n_140), .Y(n_451) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
INVx1_ASAP7_75t_L g230 ( .A(n_141), .Y(n_230) );
INVx1_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
INVx3_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
INVx4_ASAP7_75t_SL g158 ( .A(n_143), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g444 ( .A1(n_143), .A2(n_445), .B(n_449), .Y(n_444) );
BUFx3_ASAP7_75t_L g465 ( .A(n_143), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_143), .A2(n_471), .B(n_474), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_143), .A2(n_497), .B(n_500), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_143), .A2(n_506), .B(n_510), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_151), .C(n_158), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_147), .A2(n_158), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_147), .A2(n_158), .B(n_241), .C(n_242), .Y(n_240) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
INVx1_ASAP7_75t_L g491 ( .A(n_149), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_152), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g448 ( .A(n_152), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_152), .A2(n_501), .B(n_502), .Y(n_500) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g231 ( .A1(n_153), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_231) );
INVx2_ASAP7_75t_L g233 ( .A(n_153), .Y(n_233) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g174 ( .A(n_157), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g227 ( .A1(n_158), .A2(n_183), .B1(n_228), .B2(n_235), .Y(n_227) );
INVx4_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_160), .A2(n_239), .B(n_245), .Y(n_238) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_160), .A2(n_470), .B(n_477), .Y(n_469) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g176 ( .A(n_161), .Y(n_176) );
INVx4_ASAP7_75t_L g267 ( .A(n_162), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_162), .A2(n_323), .B(n_325), .Y(n_322) );
AND2x2_ASAP7_75t_L g403 ( .A(n_162), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_180), .Y(n_162) );
INVx1_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
AND2x2_ASAP7_75t_L g272 ( .A(n_163), .B(n_212), .Y(n_272) );
OR2x2_ASAP7_75t_L g301 ( .A(n_163), .B(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g315 ( .A(n_163), .Y(n_315) );
INVx3_ASAP7_75t_L g324 ( .A(n_163), .Y(n_324) );
AND2x2_ASAP7_75t_L g334 ( .A(n_163), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g367 ( .A(n_163), .B(n_273), .Y(n_367) );
AND2x2_ASAP7_75t_L g391 ( .A(n_163), .B(n_347), .Y(n_391) );
OR2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_177), .Y(n_163) );
AOI21xp5_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_175), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_173), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_169), .A2(n_255), .B(n_256), .C(n_257), .Y(n_254) );
INVx2_ASAP7_75t_L g454 ( .A(n_169), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_169), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_169), .A2(n_472), .B(n_473), .Y(n_471) );
O2A1O1Ixp5_ASAP7_75t_SL g497 ( .A1(n_169), .A2(n_223), .B(n_498), .C(n_499), .Y(n_497) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_170), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_170), .B(n_244), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_170), .A2(n_187), .B1(n_490), .B2(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g509 ( .A(n_172), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_173), .A2(n_186), .B(n_188), .Y(n_185) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_175), .A2(n_444), .B(n_455), .Y(n_443) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_175), .A2(n_458), .B(n_466), .Y(n_457) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_176), .A2(n_227), .B(n_236), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_176), .B(n_237), .Y(n_236) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_176), .A2(n_251), .B(n_258), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx3_ASAP7_75t_L g215 ( .A(n_179), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_179), .B(n_465), .C(n_481), .Y(n_480) );
AO21x1_ASAP7_75t_L g559 ( .A1(n_179), .A2(n_481), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g212 ( .A(n_180), .Y(n_212) );
AND2x2_ASAP7_75t_L g427 ( .A(n_180), .B(n_269), .Y(n_427) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_189), .B(n_190), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_183), .A2(n_252), .B(n_253), .Y(n_251) );
INVx4_ASAP7_75t_L g203 ( .A(n_187), .Y(n_203) );
INVx2_ASAP7_75t_L g220 ( .A(n_187), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_187), .A2(n_454), .B1(n_482), .B2(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_187), .A2(n_454), .B1(n_527), .B2(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_192), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_192), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_209), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_195), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g347 ( .A(n_195), .B(n_335), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_195), .B(n_324), .Y(n_409) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g269 ( .A(n_196), .Y(n_269) );
AND2x2_ASAP7_75t_L g273 ( .A(n_196), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g314 ( .A(n_196), .B(n_315), .Y(n_314) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_207), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_206), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_204), .Y(n_200) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g223 ( .A(n_205), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_209), .B(n_310), .Y(n_332) );
INVx1_ASAP7_75t_L g371 ( .A(n_209), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_209), .B(n_298), .Y(n_415) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AND2x2_ASAP7_75t_L g278 ( .A(n_210), .B(n_273), .Y(n_278) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_212), .B(n_269), .Y(n_302) );
INVx1_ASAP7_75t_L g381 ( .A(n_212), .Y(n_381) );
AOI322xp5_ASAP7_75t_L g405 ( .A1(n_213), .A2(n_320), .A3(n_380), .B1(n_406), .B2(n_408), .C1(n_410), .C2(n_412), .Y(n_405) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_214), .B(n_225), .Y(n_213) );
AND2x2_ASAP7_75t_L g260 ( .A(n_214), .B(n_238), .Y(n_260) );
INVx1_ASAP7_75t_SL g263 ( .A(n_214), .Y(n_263) );
AND2x2_ASAP7_75t_L g265 ( .A(n_214), .B(n_226), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_214), .B(n_282), .Y(n_288) );
INVx2_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
AND2x2_ASAP7_75t_L g320 ( .A(n_214), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g358 ( .A(n_214), .B(n_282), .Y(n_358) );
BUFx2_ASAP7_75t_L g375 ( .A(n_214), .Y(n_375) );
AND2x2_ASAP7_75t_L g389 ( .A(n_214), .B(n_249), .Y(n_389) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_224), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_L g462 ( .A1(n_220), .A2(n_450), .B(n_463), .C(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_220), .A2(n_511), .B(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_225), .B(n_277), .Y(n_304) );
AND2x2_ASAP7_75t_L g431 ( .A(n_225), .B(n_307), .Y(n_431) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_238), .Y(n_225) );
OR2x2_ASAP7_75t_L g276 ( .A(n_226), .B(n_277), .Y(n_276) );
INVx3_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
AND2x2_ASAP7_75t_L g327 ( .A(n_226), .B(n_250), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_226), .B(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_226), .Y(n_411) );
INVx2_ASAP7_75t_L g257 ( .A(n_229), .Y(n_257) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g262 ( .A(n_238), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g284 ( .A(n_238), .Y(n_284) );
BUFx2_ASAP7_75t_L g290 ( .A(n_238), .Y(n_290) );
AND2x2_ASAP7_75t_L g309 ( .A(n_238), .B(n_282), .Y(n_309) );
INVx3_ASAP7_75t_L g321 ( .A(n_238), .Y(n_321) );
OR2x2_ASAP7_75t_L g331 ( .A(n_238), .B(n_282), .Y(n_331) );
AOI31xp33_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_261), .A3(n_264), .B(n_266), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_260), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_248), .B(n_283), .Y(n_294) );
OR2x2_ASAP7_75t_L g318 ( .A(n_248), .B(n_288), .Y(n_318) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_249), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g339 ( .A(n_249), .B(n_331), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_249), .B(n_321), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_249), .B(n_357), .Y(n_356) );
NAND2x1_ASAP7_75t_L g384 ( .A(n_249), .B(n_320), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_249), .B(n_375), .Y(n_385) );
AND2x2_ASAP7_75t_L g397 ( .A(n_249), .B(n_282), .Y(n_397) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_257), .A2(n_446), .B(n_447), .C(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_260), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_262), .B(n_338), .Y(n_372) );
AND2x4_ASAP7_75t_L g283 ( .A(n_263), .B(n_284), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g362 ( .A(n_268), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_268), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g310 ( .A(n_269), .B(n_300), .Y(n_310) );
AND2x2_ASAP7_75t_L g404 ( .A(n_269), .B(n_274), .Y(n_404) );
INVx1_ASAP7_75t_L g429 ( .A(n_269), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B1(n_278), .B2(n_279), .C(n_285), .Y(n_270) );
CKINVDCx14_ASAP7_75t_R g291 ( .A(n_271), .Y(n_291) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_272), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_275), .B(n_326), .Y(n_345) );
INVx3_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g394 ( .A(n_276), .B(n_290), .Y(n_394) );
AND2x2_ASAP7_75t_L g308 ( .A(n_277), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g338 ( .A(n_277), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_277), .B(n_321), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g408 ( .A(n_277), .B(n_378), .C(n_409), .Y(n_408) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_278), .A2(n_342), .B(n_344), .C(n_352), .Y(n_341) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_280), .A2(n_331), .B1(n_332), .B2(n_333), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_281), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_281), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g423 ( .A(n_283), .B(n_397), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_291), .B1(n_292), .B2(n_294), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_289), .B(n_338), .Y(n_369) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_292), .A2(n_384), .B1(n_415), .B2(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_303), .B1(n_305), .B2(n_310), .C(n_311), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_301), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_301), .A2(n_312), .B1(n_318), .B2(n_319), .C(n_322), .Y(n_311) );
INVx1_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_SL g326 ( .A(n_307), .Y(n_326) );
OR2x2_ASAP7_75t_L g399 ( .A(n_307), .B(n_331), .Y(n_399) );
AND2x2_ASAP7_75t_L g401 ( .A(n_307), .B(n_309), .Y(n_401) );
INVx1_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_313), .A2(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g377 ( .A(n_313), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_335), .Y(n_351) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp33_ASAP7_75t_SL g368 ( .A(n_319), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_320), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_321), .B(n_357), .Y(n_420) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_324), .A2(n_337), .B(n_339), .C(n_340), .Y(n_336) );
NAND2x1_ASAP7_75t_SL g361 ( .A(n_324), .B(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_325), .A2(n_374), .B1(n_376), .B2(n_379), .Y(n_373) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_327), .B(n_417), .Y(n_416) );
NAND5xp2_ASAP7_75t_L g328 ( .A(n_329), .B(n_341), .C(n_359), .D(n_373), .E(n_382), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_336), .Y(n_329) );
INVx1_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_334), .A2(n_353), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_335), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_338), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_338), .B(n_404), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_348), .B2(n_350), .Y(n_344) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g426 ( .A(n_355), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_363), .B1(n_367), .B2(n_368), .C(n_370), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g410 ( .A(n_365), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g417 ( .A(n_375), .Y(n_417) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B(n_392), .C(n_405), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_390), .A2(n_415), .B(n_416), .C(n_418), .Y(n_414) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_394), .B(n_396), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_428), .B(n_430), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g714 ( .A(n_436), .Y(n_714) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR5x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_602), .C(n_660), .D(n_696), .E(n_703), .Y(n_438) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_548), .C(n_572), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_484), .B1(n_514), .B2(n_519), .C(n_529), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_441), .A2(n_683), .B(n_685), .Y(n_682) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_467), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_442), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_456), .Y(n_442) );
INVx2_ASAP7_75t_L g518 ( .A(n_443), .Y(n_518) );
AND2x2_ASAP7_75t_L g531 ( .A(n_443), .B(n_469), .Y(n_531) );
AND2x2_ASAP7_75t_L g585 ( .A(n_443), .B(n_468), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_443), .B(n_457), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B(n_453), .C(n_454), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_454), .A2(n_475), .B(n_476), .Y(n_474) );
AND2x2_ASAP7_75t_L g618 ( .A(n_456), .B(n_559), .Y(n_618) );
AND2x2_ASAP7_75t_L g651 ( .A(n_456), .B(n_469), .Y(n_651) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g558 ( .A(n_457), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g571 ( .A(n_457), .B(n_469), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_457), .B(n_559), .Y(n_578) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_457), .Y(n_587) );
AND2x2_ASAP7_75t_L g594 ( .A(n_457), .B(n_468), .Y(n_594) );
INVx1_ASAP7_75t_L g625 ( .A(n_457), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_465), .Y(n_458) );
INVx1_ASAP7_75t_L g601 ( .A(n_467), .Y(n_601) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
INVx2_ASAP7_75t_L g557 ( .A(n_468), .Y(n_557) );
AND2x2_ASAP7_75t_L g579 ( .A(n_468), .B(n_518), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_468), .B(n_625), .Y(n_630) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_469), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g702 ( .A(n_469), .B(n_666), .Y(n_702) );
INVx2_ASAP7_75t_L g516 ( .A(n_478), .Y(n_516) );
INVx3_ASAP7_75t_L g617 ( .A(n_478), .Y(n_617) );
OR2x2_ASAP7_75t_L g647 ( .A(n_478), .B(n_648), .Y(n_647) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_478), .B(n_557), .Y(n_673) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g560 ( .A(n_479), .Y(n_560) );
AOI33xp33_ASAP7_75t_L g693 ( .A1(n_484), .A2(n_531), .A3(n_545), .B1(n_617), .B2(n_694), .B3(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
OR2x2_ASAP7_75t_L g546 ( .A(n_486), .B(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_486), .B(n_543), .Y(n_605) );
OR2x2_ASAP7_75t_L g658 ( .A(n_486), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g584 ( .A(n_487), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g609 ( .A(n_487), .B(n_493), .Y(n_609) );
AND2x2_ASAP7_75t_L g676 ( .A(n_487), .B(n_521), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_487), .A2(n_576), .B(n_702), .Y(n_701) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
AND2x2_ASAP7_75t_L g555 ( .A(n_488), .B(n_525), .Y(n_555) );
AND2x2_ASAP7_75t_L g604 ( .A(n_488), .B(n_524), .Y(n_604) );
INVx2_ASAP7_75t_SL g646 ( .A(n_493), .Y(n_646) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
INVx2_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
INVx1_ASAP7_75t_L g697 ( .A(n_494), .Y(n_697) );
AND2x2_ASAP7_75t_L g710 ( .A(n_494), .B(n_591), .Y(n_710) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g537 ( .A(n_495), .Y(n_537) );
OR2x2_ASAP7_75t_L g543 ( .A(n_495), .B(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_504), .Y(n_521) );
AND2x2_ASAP7_75t_L g538 ( .A(n_504), .B(n_524), .Y(n_538) );
INVx1_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
INVx1_ASAP7_75t_L g551 ( .A(n_504), .Y(n_551) );
AND2x2_ASAP7_75t_L g576 ( .A(n_504), .B(n_525), .Y(n_576) );
INVx2_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
AND2x2_ASAP7_75t_L g685 ( .A(n_504), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_504), .B(n_566), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g540 ( .A(n_516), .Y(n_540) );
INVx1_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_516), .B(n_600), .Y(n_666) );
INVx1_ASAP7_75t_SL g626 ( .A(n_517), .Y(n_626) );
INVx2_ASAP7_75t_L g547 ( .A(n_518), .Y(n_547) );
AND2x2_ASAP7_75t_L g616 ( .A(n_518), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g632 ( .A(n_518), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g694 ( .A(n_520), .Y(n_694) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g549 ( .A(n_522), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g652 ( .A(n_522), .B(n_642), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_522), .A2(n_663), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g565 ( .A(n_523), .B(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g590 ( .A(n_523), .Y(n_590) );
INVx1_ASAP7_75t_L g614 ( .A(n_523), .Y(n_614) );
OR2x2_ASAP7_75t_L g678 ( .A(n_524), .B(n_537), .Y(n_678) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_524), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g591 ( .A(n_525), .B(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_532), .B1(n_539), .B2(n_541), .Y(n_529) );
OR2x2_ASAP7_75t_L g608 ( .A(n_530), .B(n_558), .Y(n_608) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_531), .A2(n_650), .B1(n_652), .B2(n_653), .C1(n_654), .C2(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g596 ( .A(n_535), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x2_ASAP7_75t_SL g550 ( .A(n_537), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
AND2x2_ASAP7_75t_L g669 ( .A(n_537), .B(n_538), .Y(n_669) );
INVx1_ASAP7_75t_L g687 ( .A(n_537), .Y(n_687) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g653 ( .A(n_540), .B(n_579), .Y(n_653) );
AND2x2_ASAP7_75t_L g695 ( .A(n_540), .B(n_571), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_542), .B(n_590), .Y(n_677) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_543), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g570 ( .A(n_547), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g638 ( .A(n_547), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_552), .B(n_556), .C(n_561), .Y(n_548) );
INVxp67_ASAP7_75t_L g562 ( .A(n_549), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_550), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_550), .B(n_597), .Y(n_692) );
BUFx3_ASAP7_75t_L g656 ( .A(n_551), .Y(n_656) );
INVx1_ASAP7_75t_L g563 ( .A(n_552), .Y(n_563) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g582 ( .A(n_554), .B(n_576), .Y(n_582) );
INVx1_ASAP7_75t_SL g622 ( .A(n_555), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g612 ( .A(n_557), .Y(n_612) );
AND2x2_ASAP7_75t_L g635 ( .A(n_557), .B(n_618), .Y(n_635) );
INVx1_ASAP7_75t_SL g606 ( .A(n_558), .Y(n_606) );
INVx1_ASAP7_75t_L g633 ( .A(n_559), .Y(n_633) );
AOI31xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .A3(n_564), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g654 ( .A(n_565), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
BUFx2_ASAP7_75t_L g642 ( .A(n_566), .Y(n_642) );
AND2x2_ASAP7_75t_L g670 ( .A(n_566), .B(n_591), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g643 ( .A(n_570), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_571), .B(n_638), .Y(n_684) );
AND2x2_ASAP7_75t_L g691 ( .A(n_571), .B(n_617), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_580), .C(n_595), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_577), .A2(n_604), .B1(n_605), .B2(n_606), .C(n_607), .Y(n_603) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_L g611 ( .A(n_578), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g648 ( .A(n_579), .Y(n_648) );
OAI32xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .A3(n_586), .B1(n_588), .B2(n_593), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_582), .A2(n_635), .B(n_636), .C(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI21xp5_ASAP7_75t_SL g698 ( .A1(n_590), .A2(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g659 ( .A(n_591), .Y(n_659) );
INVxp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_597), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g645 ( .A(n_597), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND4xp25_ASAP7_75t_SL g602 ( .A(n_603), .B(n_615), .C(n_634), .D(n_649), .Y(n_602) );
AND2x2_ASAP7_75t_L g641 ( .A(n_604), .B(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g663 ( .A(n_604), .B(n_656), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_606), .B(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_610), .B2(n_613), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_608), .A2(n_659), .B1(n_690), .B2(n_692), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_608), .A2(n_697), .B(n_698), .C(n_701), .Y(n_696) );
INVx2_ASAP7_75t_L g667 ( .A(n_609), .Y(n_667) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_611), .A2(n_645), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_667), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_619), .C(n_623), .Y(n_615) );
INVx1_ASAP7_75t_L g681 ( .A(n_616), .Y(n_681) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_620), .A2(n_624), .B1(n_627), .B2(n_629), .Y(n_623) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g650 ( .A(n_632), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g708 ( .A(n_635), .Y(n_708) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B1(n_644), .B2(n_647), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_642), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g699 ( .A(n_647), .Y(n_699) );
INVx1_ASAP7_75t_L g680 ( .A(n_651), .Y(n_680) );
CKINVDCx16_ASAP7_75t_R g707 ( .A(n_653), .Y(n_707) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_661), .B(n_668), .C(n_682), .D(n_688), .E(n_693), .Y(n_660) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_671), .C(n_674), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI31xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .A3(n_678), .B(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g700 ( .A(n_676), .Y(n_700) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_690), .A2(n_692), .B1(n_704), .B2(n_707), .C1(n_708), .C2(n_709), .Y(n_703) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
endmodule