module fake_jpeg_19993_n_311 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_26),
.Y(n_43)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_5),
.Y(n_28)
);

BUFx2_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_31),
.B1(n_41),
.B2(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_27),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_60),
.B(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_27),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_45),
.B1(n_51),
.B2(n_39),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_33),
.B1(n_60),
.B2(n_26),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_40),
.A3(n_29),
.B1(n_41),
.B2(n_31),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_65),
.B(n_67),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_29),
.A3(n_41),
.B1(n_31),
.B2(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_28),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_36),
.B1(n_34),
.B2(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_60),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_46),
.B(n_23),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_30),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_23),
.B(n_33),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_90),
.B1(n_91),
.B2(n_71),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_97),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_34),
.B1(n_36),
.B2(n_42),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_71),
.B(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_78),
.Y(n_91)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_64),
.B1(n_52),
.B2(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_57),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_104),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_90),
.B1(n_96),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_105),
.B1(n_49),
.B2(n_52),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_118),
.B(n_82),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_25),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_124),
.C(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_111),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_75),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_75),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_96),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_74),
.C(n_56),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_88),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_28),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_89),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_103),
.B1(n_122),
.B2(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_138),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_95),
.B(n_85),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_110),
.B(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_83),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_152),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_149),
.B(n_153),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_95),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_102),
.B(n_93),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_154),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_119),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_80),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_100),
.B1(n_88),
.B2(n_15),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_100),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_100),
.B1(n_49),
.B2(n_88),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_142),
.Y(n_181)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_105),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_181),
.Y(n_209)
);

NOR4xp25_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_108),
.C(n_118),
.D(n_122),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_165),
.A2(n_144),
.B(n_81),
.C(n_47),
.D(n_30),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_125),
.C(n_123),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_173),
.B1(n_145),
.B2(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_172),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_176),
.B(n_179),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_70),
.B1(n_62),
.B2(n_56),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_62),
.B1(n_15),
.B2(n_52),
.Y(n_179)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_23),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_182),
.B(n_81),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_21),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_93),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_81),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_77),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_184),
.A2(n_154),
.B1(n_148),
.B2(n_147),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_195),
.B1(n_173),
.B2(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_201),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_147),
.B1(n_150),
.B2(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_152),
.C(n_131),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.C(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_130),
.C(n_141),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_128),
.B(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_47),
.B1(n_16),
.B2(n_13),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_207),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_135),
.C(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_176),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_212),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_44),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_229),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_168),
.C(n_160),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_167),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_175),
.C(n_178),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_164),
.C(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_185),
.B(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_182),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_179),
.B1(n_159),
.B2(n_49),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_58),
.B1(n_15),
.B2(n_22),
.Y(n_227)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_14),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_14),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_21),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_206),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_8),
.B(n_9),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_217),
.B(n_189),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_194),
.C(n_200),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_218),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_202),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_232),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_201),
.C(n_200),
.Y(n_248)
);

AOI221xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_192),
.B1(n_195),
.B2(n_210),
.C(n_22),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_17),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_21),
.C(n_11),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_32),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_32),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_215),
.C(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_220),
.C(n_219),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_249),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_234),
.CI(n_17),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_264),
.Y(n_274)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_16),
.B(n_13),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_238),
.B(n_13),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_32),
.C(n_21),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_245),
.C(n_243),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_250),
.B1(n_239),
.B2(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_8),
.B(n_9),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_258),
.B1(n_16),
.B2(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_273),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_236),
.C(n_11),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_11),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_277),
.B(n_6),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_8),
.B(n_9),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_6),
.B(n_7),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_7),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_275),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_286),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_267),
.B(n_263),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_283),
.B(n_288),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_277),
.A2(n_253),
.B(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_11),
.C(n_32),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_19),
.B(n_4),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_280),
.B(n_19),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_300),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_19),
.B(n_1),
.C(n_2),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_19),
.C(n_7),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_19),
.C(n_291),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_281),
.A2(n_19),
.B(n_1),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_302),
.B(n_0),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_294),
.B1(n_299),
.B2(n_298),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_305),
.A2(n_306),
.B(n_303),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_302),
.C2(n_295),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_308),
.A2(n_0),
.B(n_1),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_3),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_311)
);


endmodule