module fake_jpeg_23265_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_26),
.B(n_27),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_41),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_20),
.B(n_16),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_50),
.B(n_38),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_25),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_12),
.B1(n_31),
.B2(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_44),
.B(n_36),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_23),
.C(n_15),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_58),
.C(n_12),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.C(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_18),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_46),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_41),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_43),
.B(n_37),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_72),
.B1(n_75),
.B2(n_63),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_65),
.B1(n_70),
.B2(n_59),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_58),
.C(n_37),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.C(n_67),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_54),
.C(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_76),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_90),
.B(n_80),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_69),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.C(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_93),
.C(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_87),
.C(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_86),
.C(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_10),
.B(n_6),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.C(n_98),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_102)
);


endmodule