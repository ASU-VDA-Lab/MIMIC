module real_jpeg_15518_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_641, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_641;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_578;
wire n_149;
wire n_328;
wire n_366;
wire n_620;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_638),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_0),
.B(n_639),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_62),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_62),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_1),
.A2(n_62),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_2),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_2),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_2),
.Y(n_496)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_3),
.B(n_56),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_3),
.B(n_96),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_3),
.A2(n_229),
.B1(n_538),
.B2(n_544),
.Y(n_537)
);

OAI32xp33_ASAP7_75t_L g555 ( 
.A1(n_3),
.A2(n_76),
.A3(n_479),
.B1(n_556),
.B2(n_560),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_3),
.A2(n_219),
.B1(n_570),
.B2(n_574),
.Y(n_569)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_5),
.A2(n_220),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_5),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_5),
.A2(n_261),
.B1(n_379),
.B2(n_383),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_5),
.A2(n_261),
.B1(n_482),
.B2(n_485),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_5),
.A2(n_261),
.B1(n_539),
.B2(n_543),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_136),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_6),
.A2(n_136),
.B1(n_300),
.B2(n_304),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_6),
.A2(n_136),
.B1(n_418),
.B2(n_423),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_54),
.B1(n_118),
.B2(n_123),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_7),
.A2(n_54),
.B1(n_243),
.B2(n_276),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_7),
.A2(n_54),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g465 ( 
.A(n_8),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_9),
.Y(n_248)
);

BUFx4f_ASAP7_75t_L g475 ( 
.A(n_9),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_10),
.A2(n_51),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_10),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_10),
.A2(n_226),
.B1(n_267),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_10),
.A2(n_267),
.B1(n_293),
.B2(n_510),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g516 ( 
.A1(n_10),
.A2(n_267),
.B1(n_517),
.B2(n_520),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_11),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_11),
.A2(n_209),
.B1(n_326),
.B2(n_329),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_11),
.A2(n_209),
.B1(n_490),
.B2(n_492),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_11),
.A2(n_209),
.B1(n_579),
.B2(n_581),
.Y(n_578)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_13),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_111),
.B1(n_189),
.B2(n_193),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_13),
.A2(n_111),
.B1(n_253),
.B2(n_257),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_13),
.A2(n_111),
.B1(n_289),
.B2(n_293),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_14),
.A2(n_131),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_14),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_14),
.A2(n_183),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_14),
.A2(n_183),
.B1(n_333),
.B2(n_337),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_14),
.A2(n_183),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_15),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_16),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_17),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_17),
.A2(n_214),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_17),
.A2(n_214),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_17),
.A2(n_214),
.B1(n_499),
.B2(n_501),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g135 ( 
.A(n_19),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_19),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_171),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_169),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_63),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_25),
.A2(n_48),
.B1(n_55),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_25),
.A2(n_55),
.B1(n_129),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_25),
.A2(n_55),
.B1(n_266),
.B2(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_25),
.A2(n_39),
.B1(n_325),
.B2(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_25),
.A2(n_39),
.B1(n_180),
.B2(n_411),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_26),
.A2(n_56),
.B1(n_107),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_26),
.A2(n_56),
.B1(n_260),
.B2(n_265),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_26),
.A2(n_56),
.B1(n_260),
.B2(n_352),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_34),
.B(n_39),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_32),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_35),
.Y(n_132)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_36),
.Y(n_328)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_37),
.Y(n_225)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22x1_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_43),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_44),
.Y(n_384)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_46),
.Y(n_195)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_53),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_63),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_63),
.B(n_174),
.Y(n_637)
);

FAx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_105),
.CI(n_114),
.CON(n_63),
.SN(n_63)
);

OAI21xp33_ASAP7_75t_R g64 ( 
.A1(n_65),
.A2(n_96),
.B(n_99),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_65),
.A2(n_96),
.B1(n_205),
.B2(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_65),
.A2(n_96),
.B1(n_348),
.B2(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_65),
.A2(n_96),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_97),
.B1(n_100),
.B2(n_117),
.Y(n_116)
);

OAI22x1_ASAP7_75t_L g187 ( 
.A1(n_66),
.A2(n_97),
.B1(n_117),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_66),
.A2(n_97),
.B1(n_204),
.B2(n_212),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_66),
.A2(n_97),
.B1(n_212),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_66),
.A2(n_97),
.B1(n_332),
.B2(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_66),
.A2(n_97),
.B1(n_378),
.B2(n_569),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_76),
.B(n_85),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_75),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_84),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_84),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g573 ( 
.A(n_84),
.Y(n_573)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_93),
.Y(n_584)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_94),
.Y(n_317)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_94),
.Y(n_470)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_108),
.Y(n_264)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_112),
.Y(n_353)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_113),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_127),
.C(n_137),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_115),
.A2(n_116),
.B1(n_137),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_123),
.A2(n_218),
.B1(n_223),
.B2(n_227),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_126),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_135),
.Y(n_412)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_186),
.C(n_187),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_137),
.B(n_187),
.Y(n_618)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_150),
.B(n_162),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_138),
.B(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_138),
.A2(n_150),
.B1(n_355),
.B2(n_359),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_138),
.A2(n_150),
.B1(n_162),
.B2(n_437),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_138),
.A2(n_150),
.B1(n_478),
.B2(n_481),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_138),
.A2(n_150),
.B1(n_481),
.B2(n_509),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_138),
.A2(n_150),
.B1(n_509),
.B2(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_139),
.A2(n_299),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_139),
.A2(n_288),
.B1(n_309),
.B2(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_139),
.B(n_219),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_139),
.A2(n_309),
.B1(n_595),
.B2(n_596),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_140)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_142),
.Y(n_284)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_143),
.Y(n_373)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_144),
.Y(n_493)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_145),
.Y(n_283)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_150),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_150),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_155),
.B1(n_157),
.B2(n_159),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_160),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_164),
.Y(n_397)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g358 ( 
.A(n_165),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_165),
.Y(n_580)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_196),
.B(n_636),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_184),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_176),
.A2(n_179),
.B1(n_186),
.B2(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_176),
.Y(n_625)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_179),
.A2(n_186),
.B1(n_618),
.B2(n_619),
.Y(n_617)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_185),
.B(n_624),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_188),
.Y(n_435)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_192),
.Y(n_339)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_611),
.B(n_633),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_448),
.B(n_606),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_389),
.C(n_428),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_340),
.B(n_360),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_200),
.B(n_340),
.C(n_608),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_271),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_201),
.B(n_272),
.C(n_306),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_216),
.C(n_259),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_203),
.B(n_259),
.Y(n_343)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_216),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_217),
.B(n_228),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_218),
.A2(n_219),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_219),
.B(n_467),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_SL g478 ( 
.A1(n_219),
.A2(n_466),
.B(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_219),
.B(n_534),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_219),
.B(n_305),
.Y(n_560)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_222),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_237),
.B1(n_249),
.B2(n_252),
.Y(n_228)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_229),
.A2(n_252),
.B1(n_275),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_229),
.A2(n_281),
.B(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_229),
.A2(n_489),
.B1(n_494),
.B2(n_497),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_229),
.A2(n_249),
.B1(n_516),
.B2(n_538),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_230),
.Y(n_536)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_230),
.Y(n_544)
);

INVx4_ASAP7_75t_SL g563 ( 
.A(n_230),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_231),
.Y(n_322)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_236),
.Y(n_461)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_238),
.A2(n_277),
.B1(n_367),
.B2(n_374),
.Y(n_366)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_241),
.Y(n_491)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_241),
.Y(n_500)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_247),
.Y(n_504)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_247),
.Y(n_542)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_256),
.Y(n_521)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_258),
.Y(n_370)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_306),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_285),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_273),
.A2(n_286),
.B(n_297),
.Y(n_424)
);

AOI22x1_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_277),
.A2(n_515),
.B1(n_522),
.B2(n_523),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_277),
.A2(n_367),
.B1(n_498),
.B2(n_562),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_279),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_297),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_292),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_292),
.Y(n_486)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_296),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_323),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_318),
.Y(n_307)
);

XOR2x2_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_313),
.Y(n_457)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_315),
.Y(n_510)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_331),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_324),
.B(n_331),
.C(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_345),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_342),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_346),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.C(n_354),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_354),
.Y(n_363)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_363),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_355),
.Y(n_596)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_386),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_361),
.B(n_386),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.C(n_365),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_362),
.B(n_603),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_364),
.B(n_365),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_376),
.C(n_385),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_366),
.B(n_385),
.Y(n_590)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_376),
.B(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_384),
.Y(n_575)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);

A2O1A1O1Ixp25_ASAP7_75t_L g606 ( 
.A1(n_389),
.A2(n_428),
.B(n_607),
.C(n_609),
.D(n_610),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_427),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_390),
.B(n_427),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_408),
.B1(n_425),
.B2(n_426),
.Y(n_393)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_426),
.C(n_447),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_395),
.A2(n_402),
.B1(n_403),
.B2(n_407),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_403),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_402),
.A2(n_403),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_402),
.A2(n_445),
.B1(n_622),
.B2(n_641),
.Y(n_621)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_424),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_416),
.C(n_424),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_446),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_429),
.B(n_446),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_430),
.B(n_628),
.C(n_629),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.Y(n_431)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_432),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_436),
.B(n_438),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_433),
.B(n_436),
.Y(n_438)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_438),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_438),
.A2(n_617),
.B1(n_620),
.B2(n_632),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_439),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_442),
.B2(n_445),
.Y(n_439)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_444),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_601),
.B(n_605),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_586),
.B(n_600),
.Y(n_449)
);

AOI21x1_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_551),
.B(n_585),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_512),
.B(n_550),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_487),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_453),
.B(n_487),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_476),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_454),
.A2(n_476),
.B1(n_477),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

OAI32xp33_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_458),
.A3(n_462),
.B1(n_466),
.B2(n_471),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_461),
.Y(n_519)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_472),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_505),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_488),
.B(n_507),
.C(n_511),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_508),
.B2(n_511),
.Y(n_505)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_506),
.Y(n_511)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_526),
.B(n_549),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_524),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_524),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_517),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_545),
.B(n_548),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_537),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_533),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_553),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_552),
.B(n_553),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_566),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_567),
.C(n_577),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_555),
.A2(n_561),
.B1(n_564),
.B2(n_565),
.Y(n_554)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_555),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_565),
.Y(n_593)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_561),
.Y(n_565)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_567),
.A2(n_568),
.B1(n_576),
.B2(n_577),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_573),
.Y(n_572)
);

INVx6_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_587),
.B(n_599),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_587),
.B(n_599),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_588),
.A2(n_589),
.B1(n_591),
.B2(n_592),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_594),
.C(n_597),
.Y(n_604)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_593),
.A2(n_594),
.B1(n_597),
.B2(n_598),
.Y(n_592)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_593),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_594),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_602),
.B(n_604),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_602),
.B(n_604),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_626),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_614),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_614),
.A2(n_634),
.B(n_635),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_623),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_615),
.B(n_623),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_616),
.B(n_620),
.C(n_621),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_617),
.Y(n_632)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_618),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_621),
.B(n_631),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_627),
.B(n_630),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_630),
.Y(n_634)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);


endmodule