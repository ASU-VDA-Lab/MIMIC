module fake_jpeg_29098_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_16),
.C(n_10),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_21),
.B(n_18),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_26),
.B1(n_17),
.B2(n_20),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_35),
.C(n_22),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_20),
.B1(n_11),
.B2(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_28),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_22),
.C(n_17),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_29),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_33),
.C(n_7),
.Y(n_44)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_46),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_32),
.B(n_35),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_0),
.C(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_47),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_36),
.B(n_5),
.C(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_54),
.Y(n_55)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_51),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_53),
.C(n_42),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_3),
.B(n_4),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);


endmodule