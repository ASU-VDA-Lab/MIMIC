module fake_netlist_6_4165_n_1863 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1863);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1863;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx2_ASAP7_75t_SL g186 ( 
.A(n_17),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_63),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_41),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_18),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_39),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_164),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_48),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_123),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_14),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_73),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_13),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_105),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_50),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_8),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_27),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_77),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_101),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_48),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_38),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_80),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_22),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_126),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_111),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_13),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_89),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_176),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_153),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_160),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_16),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_177),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_4),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_138),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_15),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_41),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_135),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_79),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_120),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_145),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_45),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_51),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_6),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_14),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_128),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_62),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_116),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_20),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_139),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_54),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_165),
.Y(n_273)
);

CKINVDCx11_ASAP7_75t_R g274 ( 
.A(n_88),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_106),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_29),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_7),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_86),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_68),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_42),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_141),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_109),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_148),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_108),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_60),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_26),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_157),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_32),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_24),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_81),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_64),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_72),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_57),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_27),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_85),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_98),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_11),
.Y(n_307)
);

BUFx2_ASAP7_75t_SL g308 ( 
.A(n_19),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_21),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_119),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_103),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_152),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_83),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_47),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_59),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_122),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_33),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_76),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_29),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_174),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_169),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_74),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_127),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_49),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_30),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_30),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_118),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_121),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_115),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_34),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_69),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_47),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_155),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_114),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_131),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_156),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_71),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_8),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_84),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_154),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_39),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_134),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_136),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_56),
.Y(n_350)
);

INVxp33_ASAP7_75t_R g351 ( 
.A(n_33),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_162),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_49),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_166),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_28),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_2),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_43),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_263),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_263),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_R g362 ( 
.A(n_182),
.B(n_172),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_232),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_263),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_263),
.Y(n_366)
);

BUFx6f_ASAP7_75t_SL g367 ( 
.A(n_220),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_320),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_263),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_263),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_219),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_219),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_264),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_200),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_182),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_200),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_216),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_195),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_267),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_194),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_262),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_188),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_203),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_216),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_204),
.B(n_0),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_225),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_192),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_267),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_198),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_211),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_227),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_225),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_237),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_262),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_250),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_213),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_253),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_271),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_288),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_289),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_195),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_215),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_206),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_294),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_325),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_237),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_222),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_239),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_206),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_180),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_183),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_184),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_185),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_239),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_187),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_312),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_286),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_189),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_223),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_304),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_190),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_286),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_193),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_295),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_315),
.B(n_1),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_259),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_295),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_259),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_214),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_302),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_302),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_226),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_228),
.Y(n_446)
);

NAND2x1p5_ASAP7_75t_L g447 ( 
.A(n_393),
.B(n_202),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_202),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_360),
.B(n_209),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_370),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_360),
.B(n_212),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_349),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_370),
.B(n_214),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_372),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_365),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_373),
.B(n_349),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_424),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_442),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_376),
.A2(n_217),
.B1(n_287),
.B2(n_303),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_387),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_378),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_235),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_409),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_409),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_385),
.A2(n_217),
.B1(n_287),
.B2(n_303),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_179),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_179),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_197),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_374),
.A2(n_331),
.B(n_272),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_374),
.B(n_272),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_375),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_382),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_375),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_331),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_436),
.B(n_196),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_386),
.B(n_210),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_384),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_384),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_439),
.B(n_336),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_390),
.B(n_191),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_197),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_399),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_403),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_393),
.A2(n_230),
.B(n_229),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_439),
.B(n_242),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_406),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_414),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_457),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_441),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_441),
.Y(n_527)
);

BUFx8_ASAP7_75t_SL g528 ( 
.A(n_512),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_476),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_397),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_389),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_469),
.B(n_443),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_447),
.B(n_389),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_447),
.B(n_395),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_448),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_447),
.B(n_281),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_476),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_447),
.B(n_186),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_474),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_458),
.B(n_385),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_455),
.B(n_395),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_443),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_508),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_455),
.B(n_404),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_517),
.A2(n_336),
.B1(n_308),
.B2(n_438),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_460),
.B(n_404),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_477),
.A2(n_221),
.B1(n_326),
.B2(n_309),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_477),
.B(n_412),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_456),
.B(n_412),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_478),
.B(n_419),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_448),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx8_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

CKINVDCx6p67_ASAP7_75t_R g563 ( 
.A(n_459),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_474),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_469),
.B(n_496),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_419),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_515),
.Y(n_568)
);

BUFx4f_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_505),
.B(n_270),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_517),
.A2(n_505),
.B1(n_518),
.B2(n_451),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_467),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_422),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_474),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_486),
.B(n_432),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_486),
.B(n_445),
.C(n_432),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_465),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_465),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_489),
.B(n_445),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_191),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_496),
.B(n_444),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_450),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_489),
.B(n_446),
.C(n_402),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_491),
.B(n_446),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_491),
.B(n_363),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_472),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_517),
.A2(n_417),
.B1(n_420),
.B2(n_418),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_506),
.B(n_362),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_506),
.B(n_364),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_479),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_457),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_453),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_453),
.Y(n_603)
);

INVxp33_ASAP7_75t_SL g604 ( 
.A(n_472),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_468),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_468),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_521),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_521),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_521),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_505),
.A2(n_319),
.B1(n_191),
.B2(n_205),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_471),
.B(n_181),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_480),
.Y(n_615)
);

OAI21xp33_ASAP7_75t_SL g616 ( 
.A1(n_495),
.A2(n_444),
.B(n_283),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_471),
.B(n_273),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_521),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_513),
.B(n_364),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_479),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_471),
.B(n_224),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_479),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_480),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_518),
.B(n_369),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_483),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_479),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_483),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_483),
.Y(n_631)
);

CKINVDCx6p67_ASAP7_75t_R g632 ( 
.A(n_518),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_504),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_451),
.A2(n_324),
.B1(n_276),
.B2(n_284),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_504),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_515),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_470),
.B(n_369),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_479),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_479),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_451),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_451),
.B(n_359),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_496),
.B(n_388),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_470),
.B(n_300),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_510),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_482),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_457),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_482),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_482),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_514),
.B(n_367),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_515),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_484),
.B(n_356),
.C(n_274),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_515),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_482),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_510),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_519),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_519),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_482),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_502),
.B(n_359),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_367),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_457),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_516),
.B(n_359),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_519),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_484),
.A2(n_340),
.B1(n_346),
.B2(n_357),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_519),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_519),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_464),
.B(n_231),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_502),
.A2(n_510),
.B1(n_523),
.B2(n_522),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_502),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_522),
.A2(n_205),
.B1(n_321),
.B2(n_319),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_541),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_541),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_584),
.B(n_205),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_556),
.B(n_530),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_639),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_647),
.A2(n_340),
.B1(n_394),
.B2(n_380),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_663),
.B(n_391),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_523),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_578),
.B(n_199),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_532),
.B(n_519),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_543),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_642),
.B(n_482),
.Y(n_687)
);

NOR2x1_ASAP7_75t_L g688 ( 
.A(n_579),
.B(n_454),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_638),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_543),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_638),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_554),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_584),
.B(n_205),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_584),
.B(n_256),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_529),
.B(n_473),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_565),
.B(n_485),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_565),
.B(n_485),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_551),
.A2(n_495),
.B1(n_310),
.B2(n_318),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_648),
.B(n_199),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_566),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_485),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_567),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_663),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_644),
.Y(n_705)
);

NOR2xp67_ASAP7_75t_L g706 ( 
.A(n_588),
.B(n_473),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_673),
.B(n_485),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_549),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_574),
.B(n_256),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_561),
.B(n_485),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_575),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_648),
.B(n_256),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_561),
.B(n_485),
.Y(n_714)
);

BUFx8_ASAP7_75t_L g715 ( 
.A(n_566),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_590),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_659),
.B(n_256),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_570),
.B(n_575),
.Y(n_719)
);

BUFx12f_ASAP7_75t_L g720 ( 
.A(n_530),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_646),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_534),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_534),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_582),
.B(n_485),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_537),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_576),
.B(n_475),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_582),
.B(n_520),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_659),
.B(n_520),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_614),
.B(n_520),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_646),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_617),
.B(n_520),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_549),
.B(n_520),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_475),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_604),
.A2(n_495),
.B1(n_327),
.B2(n_306),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_609),
.B(n_498),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_609),
.B(n_498),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_610),
.B(n_498),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_620),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_540),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_537),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_526),
.B(n_400),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_610),
.B(n_498),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_546),
.B(n_201),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_531),
.A2(n_401),
.B1(n_416),
.B2(n_421),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_535),
.B(n_201),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_559),
.Y(n_746)
);

CKINVDCx11_ASAP7_75t_R g747 ( 
.A(n_563),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_647),
.A2(n_338),
.B1(n_332),
.B2(n_311),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_558),
.B(n_539),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_620),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_611),
.B(n_498),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_L g753 ( 
.A1(n_591),
.A2(n_346),
.B1(n_350),
.B2(n_353),
.C(n_357),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_542),
.B(n_351),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_550),
.B(n_207),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_672),
.A2(n_592),
.B1(n_647),
.B2(n_552),
.C(n_668),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_585),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_611),
.B(n_498),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_618),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_559),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_656),
.B(n_319),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_618),
.B(n_498),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_572),
.B(n_501),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_545),
.B(n_555),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_616),
.A2(n_524),
.B(n_509),
.C(n_507),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_557),
.B(n_350),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_572),
.B(n_501),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_572),
.B(n_501),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_536),
.B(n_319),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_526),
.B(n_527),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_612),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_612),
.B(n_321),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_572),
.B(n_321),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_583),
.B(n_207),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_591),
.A2(n_553),
.B1(n_668),
.B2(n_353),
.C(n_343),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_527),
.B(n_501),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_528),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_533),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_589),
.B(n_208),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_539),
.B(n_524),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_586),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_533),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_626),
.B(n_208),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_547),
.B(n_524),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_616),
.B(n_321),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_547),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_647),
.A2(n_492),
.B(n_509),
.C(n_507),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_540),
.B(n_427),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_619),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_580),
.B(n_501),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_619),
.Y(n_791)
);

NOR2x1p5_ASAP7_75t_L g792 ( 
.A(n_563),
.B(n_236),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_544),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_632),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_647),
.B(n_481),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_594),
.B(n_501),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_542),
.A2(n_430),
.B1(n_435),
.B2(n_437),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_595),
.B(n_285),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_622),
.B(n_501),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_586),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_653),
.B(n_285),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_643),
.B(n_344),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_587),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_664),
.B(n_440),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_587),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_624),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_580),
.B(n_304),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_666),
.B(n_243),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_542),
.B(n_344),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_613),
.B(n_562),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_544),
.B(n_454),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_624),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_580),
.B(n_304),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_538),
.A2(n_635),
.B1(n_542),
.B2(n_633),
.Y(n_814)
);

O2A1O1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_542),
.A2(n_481),
.B(n_503),
.C(n_500),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_544),
.B(n_454),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_593),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_538),
.B(n_244),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_671),
.B(n_345),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_544),
.B(n_464),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_593),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_562),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_548),
.B(n_464),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_548),
.B(n_464),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_548),
.B(n_490),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_635),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_627),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_548),
.B(n_490),
.Y(n_828)
);

NAND2x1_ASAP7_75t_L g829 ( 
.A(n_571),
.B(n_465),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_633),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_560),
.B(n_490),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_560),
.B(n_493),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_560),
.B(n_493),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_627),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_632),
.B(n_538),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_634),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_580),
.B(n_304),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_596),
.A2(n_487),
.B(n_503),
.C(n_500),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_568),
.A2(n_457),
.B(n_461),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_635),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_628),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_580),
.B(n_345),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_560),
.B(n_493),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_822),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_680),
.B(n_538),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_764),
.A2(n_603),
.B(n_605),
.C(n_607),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_717),
.B(n_538),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_769),
.A2(n_641),
.B(n_640),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_709),
.A2(n_635),
.B1(n_634),
.B2(n_636),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_676),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_703),
.B(n_628),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_822),
.B(n_640),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_764),
.A2(n_675),
.B1(n_670),
.B2(n_669),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_770),
.B(n_630),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_721),
.B(n_262),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_749),
.B(n_487),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_685),
.B(n_630),
.Y(n_857)
);

AOI33xp33_ASAP7_75t_L g858 ( 
.A1(n_753),
.A2(n_488),
.A3(n_492),
.B1(n_494),
.B2(n_497),
.B3(n_499),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_685),
.B(n_564),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_822),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_676),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_743),
.B(n_564),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_774),
.B(n_248),
.C(n_247),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_743),
.B(n_564),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_810),
.A2(n_569),
.B(n_568),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_755),
.B(n_564),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_755),
.B(n_573),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_784),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_729),
.A2(n_569),
.B(n_568),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_731),
.A2(n_799),
.B(n_822),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_712),
.B(n_573),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_784),
.B(n_573),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_677),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_719),
.B(n_573),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_686),
.B(n_577),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_704),
.B(n_641),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_697),
.A2(n_569),
.B(n_562),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_756),
.A2(n_596),
.B(n_602),
.C(n_603),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_749),
.B(n_488),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_698),
.A2(n_652),
.B(n_651),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_774),
.A2(n_607),
.B(n_602),
.C(n_605),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_720),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_690),
.B(n_577),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_775),
.B(n_352),
.C(n_348),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_733),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_779),
.A2(n_494),
.B(n_497),
.C(n_499),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_730),
.A2(n_636),
.B(n_600),
.C(n_601),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_692),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_577),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_779),
.A2(n_674),
.B(n_277),
.C(n_299),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_709),
.A2(n_652),
.B(n_651),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_692),
.Y(n_892)
);

AO22x1_ASAP7_75t_L g893 ( 
.A1(n_809),
.A2(n_268),
.B1(n_251),
.B2(n_261),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_776),
.A2(n_693),
.B(n_678),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_814),
.B(n_580),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_694),
.B(n_577),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_687),
.A2(n_606),
.B(n_571),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_694),
.B(n_597),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_741),
.B(n_269),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_678),
.A2(n_621),
.B(n_597),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_683),
.B(n_275),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_814),
.B(n_581),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_716),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_716),
.B(n_597),
.Y(n_904)
);

O2A1O1Ixp5_ASAP7_75t_L g905 ( 
.A1(n_769),
.A2(n_693),
.B(n_695),
.C(n_713),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_733),
.B(n_581),
.Y(n_906)
);

AO21x1_ASAP7_75t_L g907 ( 
.A1(n_785),
.A2(n_645),
.B(n_637),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_722),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_771),
.B(n_597),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_795),
.A2(n_637),
.B1(n_670),
.B2(n_669),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_702),
.A2(n_606),
.B(n_571),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_759),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_707),
.A2(n_606),
.B(n_598),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_796),
.A2(n_606),
.B(n_598),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_780),
.B(n_621),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_795),
.B(n_581),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_722),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_785),
.A2(n_675),
.B(n_667),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_728),
.A2(n_667),
.B(n_654),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_SL g920 ( 
.A1(n_695),
.A2(n_660),
.B(n_661),
.C(n_655),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_726),
.B(n_621),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_701),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_780),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_789),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_713),
.A2(n_661),
.B(n_654),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_791),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_744),
.B(n_278),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_682),
.B(n_280),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_732),
.A2(n_665),
.B(n_525),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_708),
.B(n_581),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_708),
.B(n_581),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_747),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_696),
.B(n_621),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_752),
.B(n_623),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_763),
.A2(n_665),
.B(n_525),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_723),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_806),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_684),
.B(n_623),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_757),
.B(n_623),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_766),
.B(n_623),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_767),
.A2(n_665),
.B(n_598),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_699),
.A2(n_662),
.B(n_629),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_777),
.B(n_645),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_778),
.B(n_629),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_723),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_782),
.B(n_629),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_699),
.A2(n_662),
.B(n_629),
.Y(n_947)
);

BUFx12f_ASAP7_75t_L g948 ( 
.A(n_715),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_812),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_786),
.A2(n_290),
.B(n_292),
.C(n_293),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_696),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_734),
.A2(n_662),
.B(n_649),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_689),
.B(n_649),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_794),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_768),
.A2(n_598),
.B(n_525),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_706),
.A2(n_826),
.B1(n_835),
.B2(n_809),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_650),
.B(n_525),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_835),
.A2(n_657),
.B1(n_655),
.B2(n_660),
.Y(n_958)
);

BUFx2_ASAP7_75t_SL g959 ( 
.A(n_739),
.Y(n_959)
);

OAI321xp33_ASAP7_75t_L g960 ( 
.A1(n_783),
.A2(n_367),
.A3(n_258),
.B1(n_313),
.B2(n_220),
.C(n_233),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_797),
.B(n_296),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_691),
.B(n_649),
.Y(n_962)
);

AOI33xp33_ASAP7_75t_L g963 ( 
.A1(n_748),
.A2(n_305),
.A3(n_330),
.B1(n_317),
.B2(n_314),
.B3(n_307),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_816),
.A2(n_650),
.B(n_581),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_705),
.B(n_658),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_710),
.B(n_658),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_840),
.B(n_658),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_734),
.A2(n_658),
.B(n_599),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_827),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_793),
.A2(n_650),
.B(n_631),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_834),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_787),
.B(n_599),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_765),
.A2(n_601),
.B(n_600),
.C(n_608),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_715),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_841),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_748),
.A2(n_608),
.B1(n_220),
.B2(n_233),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_830),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_783),
.B(n_772),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_711),
.A2(n_631),
.B(n_625),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_724),
.A2(n_823),
.B(n_820),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_836),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_798),
.A2(n_348),
.B(n_354),
.C(n_352),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_794),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_824),
.A2(n_650),
.B(n_625),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_815),
.B(n_615),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_738),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_714),
.A2(n_615),
.B(n_457),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_772),
.B(n_234),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_725),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_725),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_740),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_798),
.B(n_238),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_836),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_727),
.A2(n_465),
.B(n_461),
.Y(n_994)
);

AO21x1_ASAP7_75t_L g995 ( 
.A1(n_718),
.A2(n_233),
.B(n_258),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_718),
.B(n_240),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_843),
.A2(n_457),
.B(n_461),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_773),
.A2(n_745),
.B(n_751),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_681),
.B(n_354),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_818),
.A2(n_252),
.B1(n_245),
.B2(n_342),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_804),
.B(n_241),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_700),
.B(n_246),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_L g1003 ( 
.A(n_802),
.B(n_254),
.C(n_249),
.Y(n_1003)
);

BUFx4f_ASAP7_75t_L g1004 ( 
.A(n_754),
.Y(n_1004)
);

CKINVDCx10_ASAP7_75t_R g1005 ( 
.A(n_754),
.Y(n_1005)
);

OAI321xp33_ASAP7_75t_L g1006 ( 
.A1(n_802),
.A2(n_808),
.A3(n_801),
.B1(n_750),
.B2(n_754),
.C(n_819),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_740),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_830),
.B(n_255),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_825),
.A2(n_828),
.B(n_831),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_746),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_746),
.B(n_257),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_792),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_760),
.B(n_265),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_761),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_688),
.B(n_67),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_838),
.A2(n_316),
.B(n_266),
.C(n_291),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_760),
.B(n_297),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_781),
.B(n_298),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_781),
.B(n_334),
.Y(n_1019)
);

OAI321xp33_ASAP7_75t_L g1020 ( 
.A1(n_773),
.A2(n_313),
.A3(n_258),
.B1(n_4),
.B2(n_5),
.C(n_9),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_829),
.A2(n_465),
.B(n_511),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_790),
.A2(n_465),
.B(n_461),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_800),
.B(n_337),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_832),
.A2(n_461),
.B(n_301),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_761),
.A2(n_341),
.B(n_339),
.C(n_329),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_833),
.A2(n_465),
.B(n_511),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_842),
.A2(n_323),
.B(n_322),
.C(n_313),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_735),
.A2(n_465),
.B(n_511),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_736),
.A2(n_461),
.B(n_511),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_927),
.B(n_788),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_870),
.A2(n_865),
.B(n_859),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_885),
.B(n_803),
.Y(n_1032)
);

AO22x1_ASAP7_75t_L g1033 ( 
.A1(n_884),
.A2(n_800),
.B1(n_817),
.B2(n_805),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_873),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_982),
.A2(n_737),
.B(n_742),
.C(n_758),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1003),
.A2(n_762),
.B1(n_805),
.B2(n_821),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_877),
.A2(n_839),
.B(n_790),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_873),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_901),
.B(n_821),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_861),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_850),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_899),
.B(n_817),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_885),
.B(n_803),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_851),
.B(n_837),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_851),
.B(n_813),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_888),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_922),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_884),
.B(n_807),
.C(n_3),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_999),
.B(n_807),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_999),
.B(n_2),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_956),
.A2(n_10),
.B1(n_12),
.B2(n_17),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_1014),
.B(n_151),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_869),
.A2(n_102),
.B(n_150),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_1014),
.B(n_147),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_903),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_978),
.A2(n_12),
.B(n_19),
.C(n_21),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_921),
.B(n_511),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_856),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_959),
.B(n_144),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_932),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_857),
.A2(n_97),
.B(n_137),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_921),
.B(n_511),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1003),
.B(n_22),
.C(n_23),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_954),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_845),
.B(n_847),
.Y(n_1065)
);

OR2x6_ASAP7_75t_SL g1066 ( 
.A(n_961),
.B(n_24),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_928),
.B(n_855),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_854),
.B(n_511),
.Y(n_1068)
);

INVx8_ASAP7_75t_L g1069 ( 
.A(n_933),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_856),
.Y(n_1070)
);

AOI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_992),
.A2(n_25),
.B(n_26),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_951),
.B(n_125),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_868),
.B(n_511),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_982),
.A2(n_25),
.B(n_31),
.C(n_35),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_858),
.B(n_124),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_862),
.A2(n_112),
.B(n_100),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_940),
.B(n_35),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_950),
.A2(n_36),
.B(n_37),
.C(n_40),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_986),
.Y(n_1079)
);

CKINVDCx11_ASAP7_75t_R g1080 ( 
.A(n_948),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_1002),
.A2(n_940),
.B(n_905),
.C(n_863),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_923),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_93),
.B(n_92),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_892),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_849),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_858),
.B(n_91),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_844),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_967),
.B(n_90),
.Y(n_1088)
);

NAND3xp33_ASAP7_75t_SL g1089 ( 
.A(n_1002),
.B(n_50),
.C(n_51),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_954),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_1006),
.B(n_78),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_951),
.B(n_923),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_950),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_879),
.B(n_52),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_879),
.B(n_986),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_912),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_866),
.A2(n_53),
.B(n_56),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1012),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_924),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_926),
.B(n_57),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_867),
.A2(n_947),
.B(n_942),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_933),
.B(n_889),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_882),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_849),
.A2(n_58),
.B1(n_976),
.B2(n_1025),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_894),
.A2(n_58),
.B(n_889),
.C(n_938),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1015),
.B(n_943),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_882),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_937),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_911),
.A2(n_913),
.B(n_952),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_983),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_908),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1001),
.B(n_983),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_949),
.B(n_969),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1025),
.A2(n_960),
.B(n_886),
.C(n_1020),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_893),
.B(n_967),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_974),
.B(n_1015),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_917),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_938),
.A2(n_886),
.B(n_878),
.C(n_971),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_860),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_988),
.A2(n_1000),
.B1(n_916),
.B2(n_996),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_878),
.A2(n_975),
.B(n_963),
.C(n_968),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_963),
.A2(n_881),
.B(n_944),
.C(n_909),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_916),
.A2(n_909),
.B1(n_995),
.B2(n_876),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_993),
.B(n_944),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_890),
.A2(n_881),
.B(n_846),
.C(n_876),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_981),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_976),
.B(n_860),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_993),
.B(n_874),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_915),
.A2(n_902),
.B1(n_895),
.B2(n_998),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_906),
.A2(n_910),
.B1(n_931),
.B2(n_930),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_936),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1004),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_914),
.A2(n_897),
.B(n_852),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_981),
.B(n_934),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_939),
.B(n_946),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_890),
.B(n_1027),
.C(n_902),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_945),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_SL g1138 ( 
.A(n_895),
.B(n_906),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1004),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_977),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1008),
.B(n_1011),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_930),
.B(n_931),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_852),
.A2(n_941),
.B(n_955),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_989),
.B(n_990),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_958),
.B(n_872),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_991),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_935),
.A2(n_957),
.B(n_1009),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1007),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1016),
.A2(n_846),
.B(n_953),
.C(n_973),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_1010),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_962),
.B(n_966),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1013),
.B(n_1017),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_L g1153 ( 
.A(n_1018),
.B(n_1023),
.Y(n_1153)
);

CKINVDCx6p67_ASAP7_75t_R g1154 ( 
.A(n_1005),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1022),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1019),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_875),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_965),
.B(n_871),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_972),
.A2(n_985),
.B(n_920),
.C(n_887),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_953),
.B(n_853),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_907),
.B(n_918),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_883),
.B(n_904),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_848),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_880),
.A2(n_929),
.B(n_980),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_896),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_891),
.A2(n_900),
.B(n_972),
.C(n_985),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_898),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_964),
.A2(n_970),
.B(n_979),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_925),
.A2(n_1024),
.B1(n_920),
.B2(n_1026),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_994),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_919),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_1021),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_984),
.A2(n_987),
.B(n_1028),
.C(n_1029),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_997),
.B(n_770),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_978),
.A2(n_764),
.B(n_680),
.C(n_756),
.Y(n_1175)
);

BUFx4_ASAP7_75t_SL g1176 ( 
.A(n_986),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_978),
.B(n_770),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_856),
.B(n_879),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1014),
.A2(n_679),
.B1(n_680),
.B2(n_717),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_959),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_851),
.B(n_680),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1003),
.A2(n_764),
.B1(n_680),
.B2(n_884),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_922),
.B(n_717),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_1121),
.A2(n_1086),
.B(n_1075),
.C(n_1081),
.Y(n_1184)
);

INVx8_ASAP7_75t_L g1185 ( 
.A(n_1069),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1095),
.B(n_1178),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1181),
.B(n_1177),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1107),
.B(n_1106),
.Y(n_1188)
);

AO21x2_ASAP7_75t_L g1189 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_1031),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1096),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1168),
.A2(n_1147),
.B(n_1161),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_SL g1192 ( 
.A(n_1050),
.B(n_1085),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1182),
.A2(n_1049),
.B(n_1175),
.C(n_1114),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1075),
.A2(n_1086),
.B(n_1125),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1119),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1155),
.A2(n_1159),
.B(n_1174),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1155),
.A2(n_1174),
.B(n_1101),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1162),
.A2(n_1053),
.B(n_1035),
.Y(n_1198)
);

AOI31xp67_ASAP7_75t_L g1199 ( 
.A1(n_1169),
.A2(n_1123),
.A3(n_1065),
.B(n_1120),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1177),
.B(n_1067),
.Y(n_1200)
);

AOI221x1_ASAP7_75t_L g1201 ( 
.A1(n_1104),
.A2(n_1105),
.B1(n_1063),
.B2(n_1089),
.C(n_1051),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1152),
.A2(n_1141),
.B(n_1166),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1042),
.B(n_1039),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1149),
.A2(n_1118),
.B(n_1122),
.Y(n_1204)
);

AOI221x1_ASAP7_75t_L g1205 ( 
.A1(n_1104),
.A2(n_1063),
.B1(n_1085),
.B2(n_1071),
.C(n_1138),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1173),
.A2(n_1158),
.A3(n_1135),
.B(n_1077),
.Y(n_1206)
);

AOI31xp67_ASAP7_75t_L g1207 ( 
.A1(n_1036),
.A2(n_1145),
.A3(n_1088),
.B(n_1127),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1129),
.A2(n_1088),
.B(n_1171),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1183),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1033),
.A2(n_1124),
.B(n_1128),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1178),
.B(n_1094),
.Y(n_1211)
);

AO32x2_ASAP7_75t_L g1212 ( 
.A1(n_1170),
.A2(n_1146),
.A3(n_1136),
.B1(n_1074),
.B2(n_1093),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_1060),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1128),
.A2(n_1153),
.B(n_1044),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1179),
.B(n_1030),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1099),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1134),
.A2(n_1144),
.B(n_1165),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1095),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1110),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1115),
.B(n_1160),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1116),
.B(n_1132),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1071),
.A2(n_1048),
.B1(n_1078),
.B2(n_1056),
.C(n_1082),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1108),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1045),
.A2(n_1068),
.B(n_1062),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1113),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1167),
.B(n_1157),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1047),
.B(n_1112),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1041),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1069),
.B(n_1116),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1119),
.A2(n_1102),
.B(n_1151),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1058),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1068),
.A2(n_1057),
.B(n_1091),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1046),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1055),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1119),
.A2(n_1151),
.B(n_1142),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1142),
.A2(n_1061),
.B(n_1076),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1130),
.A2(n_1083),
.B(n_1097),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1034),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1142),
.A2(n_1054),
.B(n_1052),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1140),
.B(n_1100),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1116),
.A2(n_1150),
.B1(n_1156),
.B2(n_1038),
.Y(n_1241)
);

AOI221xp5_ASAP7_75t_L g1242 ( 
.A1(n_1070),
.A2(n_1079),
.B1(n_1180),
.B2(n_1103),
.C(n_1092),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1163),
.A2(n_1032),
.B(n_1043),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1040),
.B(n_1084),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1069),
.B(n_1117),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1111),
.B(n_1137),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1148),
.A2(n_1072),
.B(n_1131),
.C(n_1073),
.Y(n_1247)
);

BUFx12f_ASAP7_75t_L g1248 ( 
.A(n_1080),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1139),
.B(n_1146),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1176),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1064),
.B(n_1090),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1087),
.A2(n_1163),
.B(n_1172),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1170),
.A2(n_1172),
.B(n_1150),
.Y(n_1253)
);

AO21x1_ASAP7_75t_L g1254 ( 
.A1(n_1172),
.A2(n_1066),
.B(n_1126),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1090),
.B(n_1098),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1059),
.B(n_1154),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1059),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1182),
.A2(n_764),
.B(n_1049),
.C(n_1050),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1259)
);

CKINVDCx16_ASAP7_75t_R g1260 ( 
.A(n_1107),
.Y(n_1260)
);

OR2x6_ASAP7_75t_L g1261 ( 
.A(n_1069),
.B(n_1116),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1064),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1030),
.B(n_476),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1110),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1075),
.A2(n_1086),
.B(n_1125),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1182),
.A2(n_764),
.B(n_1049),
.C(n_1050),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1030),
.B(n_476),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1181),
.B(n_680),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1096),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1047),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1047),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1110),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1179),
.B(n_679),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1121),
.A2(n_1075),
.B(n_1086),
.C(n_1081),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1110),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1149),
.A2(n_1118),
.A3(n_1081),
.B(n_881),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1096),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1182),
.A2(n_1014),
.B1(n_1050),
.B2(n_1104),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1067),
.B(n_741),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1047),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1085),
.A2(n_1050),
.B1(n_1104),
.B2(n_1114),
.C(n_1175),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1050),
.A2(n_1104),
.B1(n_1105),
.B2(n_1063),
.C(n_1003),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1101),
.A2(n_1175),
.B(n_1166),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1164),
.A2(n_1101),
.B(n_1031),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1095),
.B(n_1178),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1096),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1182),
.A2(n_764),
.B(n_1049),
.C(n_1050),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1149),
.A2(n_1118),
.A3(n_1081),
.B(n_881),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1030),
.B(n_476),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1037),
.A2(n_1143),
.B(n_1133),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1182),
.A2(n_1014),
.B1(n_1050),
.B2(n_1104),
.Y(n_1300)
);

AO21x1_ASAP7_75t_L g1301 ( 
.A1(n_1104),
.A2(n_1138),
.B(n_1114),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1067),
.B(n_741),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1182),
.A2(n_1014),
.B1(n_1050),
.B2(n_1104),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_1178),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1128),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1037),
.A2(n_1143),
.B(n_1133),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_SL g1307 ( 
.A(n_1182),
.B(n_679),
.C(n_764),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1181),
.B(n_680),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1149),
.A2(n_1118),
.A3(n_1081),
.B(n_881),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1126),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1311)
);

BUFx2_ASAP7_75t_SL g1312 ( 
.A(n_1064),
.Y(n_1312)
);

NOR4xp25_ASAP7_75t_L g1313 ( 
.A(n_1089),
.B(n_1074),
.C(n_1063),
.D(n_1078),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_SL g1314 ( 
.A1(n_1065),
.A2(n_1071),
.B(n_1161),
.C(n_769),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1050),
.A2(n_764),
.B1(n_884),
.B2(n_1182),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1121),
.A2(n_1075),
.B(n_1086),
.C(n_1081),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1037),
.A2(n_1143),
.B(n_1133),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1119),
.B(n_1106),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1320)
);

AO22x2_ASAP7_75t_L g1321 ( 
.A1(n_1104),
.A2(n_1085),
.B1(n_1063),
.B2(n_1089),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1110),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1080),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_SL g1324 ( 
.A(n_1050),
.B(n_679),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1128),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1064),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1327)
);

BUFx2_ASAP7_75t_R g1328 ( 
.A(n_1060),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_1109),
.B(n_822),
.Y(n_1329)
);

AO32x2_ASAP7_75t_L g1330 ( 
.A1(n_1104),
.A2(n_1085),
.A3(n_826),
.B1(n_1170),
.B2(n_1146),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1264),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1192),
.A2(n_1315),
.B1(n_1284),
.B2(n_1303),
.Y(n_1332)
);

BUFx10_ASAP7_75t_L g1333 ( 
.A(n_1249),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1275),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1219),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1216),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1323),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1227),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1276),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1282),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1244),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1203),
.B(n_1220),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1262),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1192),
.A2(n_1324),
.B1(n_1321),
.B2(n_1303),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1223),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1277),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1324),
.A2(n_1315),
.B1(n_1307),
.B2(n_1300),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1272),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1258),
.A2(n_1269),
.B1(n_1294),
.B2(n_1308),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1262),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1321),
.A2(n_1284),
.B1(n_1300),
.B2(n_1215),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1301),
.A2(n_1222),
.B1(n_1278),
.B2(n_1204),
.Y(n_1352)
);

BUFx8_ASAP7_75t_SL g1353 ( 
.A(n_1248),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1262),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1283),
.Y(n_1355)
);

BUFx8_ASAP7_75t_L g1356 ( 
.A(n_1281),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1204),
.A2(n_1194),
.B1(n_1267),
.B2(n_1187),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1213),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1322),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1271),
.A2(n_1193),
.B1(n_1325),
.B2(n_1305),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1202),
.A2(n_1200),
.B1(n_1254),
.B2(n_1290),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1263),
.A2(n_1270),
.B1(n_1297),
.B2(n_1240),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1293),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1225),
.B(n_1285),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1213),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1290),
.A2(n_1237),
.B1(n_1239),
.B2(n_1302),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1287),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1326),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1237),
.A2(n_1257),
.B1(n_1288),
.B2(n_1256),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1275),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1211),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1326),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1241),
.A2(n_1288),
.B1(n_1188),
.B2(n_1242),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1289),
.A2(n_1201),
.B(n_1205),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1228),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1256),
.A2(n_1226),
.B1(n_1241),
.B2(n_1214),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1218),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1185),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1328),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1233),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1234),
.A2(n_1224),
.B1(n_1221),
.B2(n_1209),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1224),
.A2(n_1221),
.B1(n_1209),
.B2(n_1238),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1218),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1231),
.A2(n_1319),
.B1(n_1261),
.B2(n_1229),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1229),
.A2(n_1261),
.B1(n_1231),
.B2(n_1260),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1330),
.A2(n_1208),
.B1(n_1313),
.B2(n_1312),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1250),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1229),
.A2(n_1261),
.B1(n_1319),
.B2(n_1245),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1217),
.Y(n_1389)
);

INVx6_ASAP7_75t_L g1390 ( 
.A(n_1195),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1186),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1236),
.A2(n_1208),
.B1(n_1232),
.B2(n_1191),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1310),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1186),
.B(n_1292),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1310),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1292),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1184),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1279),
.Y(n_1398)
);

INVx6_ASAP7_75t_L g1399 ( 
.A(n_1185),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1304),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1304),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1230),
.A2(n_1235),
.B1(n_1210),
.B2(n_1251),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1316),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1232),
.A2(n_1191),
.B1(n_1313),
.B2(n_1189),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1255),
.A2(n_1330),
.B1(n_1185),
.B2(n_1243),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1253),
.B(n_1252),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1189),
.A2(n_1196),
.B1(n_1291),
.B2(n_1197),
.Y(n_1407)
);

BUFx8_ASAP7_75t_L g1408 ( 
.A(n_1212),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1291),
.A2(n_1198),
.B1(n_1330),
.B2(n_1280),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1259),
.A2(n_1286),
.B1(n_1327),
.B2(n_1320),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1314),
.Y(n_1411)
);

BUFx4f_ASAP7_75t_SL g1412 ( 
.A(n_1212),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1247),
.A2(n_1295),
.B1(n_1317),
.B2(n_1311),
.Y(n_1413)
);

CKINVDCx14_ASAP7_75t_R g1414 ( 
.A(n_1207),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1265),
.A2(n_1274),
.B1(n_1298),
.B2(n_1273),
.Y(n_1415)
);

BUFx4f_ASAP7_75t_SL g1416 ( 
.A(n_1212),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1329),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1266),
.A2(n_1268),
.B1(n_1199),
.B2(n_1296),
.Y(n_1418)
);

INVx6_ASAP7_75t_L g1419 ( 
.A(n_1206),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1309),
.A2(n_1299),
.B1(n_1306),
.B2(n_1318),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1206),
.B(n_1203),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1246),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1323),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1219),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1192),
.A2(n_1324),
.B1(n_380),
.B2(n_391),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1190),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1190),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1246),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1190),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1275),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1262),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1323),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1323),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1323),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_SL g1440 ( 
.A(n_1213),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1187),
.B(n_1203),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1192),
.A2(n_1050),
.B1(n_1315),
.B2(n_1300),
.Y(n_1443)
);

INVx8_ASAP7_75t_L g1444 ( 
.A(n_1185),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1315),
.A2(n_484),
.B(n_744),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_SL g1446 ( 
.A(n_1213),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1190),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1246),
.Y(n_1448)
);

OAI22x1_ASAP7_75t_L g1449 ( 
.A1(n_1315),
.A2(n_1182),
.B1(n_1050),
.B2(n_1278),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1262),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1190),
.Y(n_1451)
);

BUFx10_ASAP7_75t_L g1452 ( 
.A(n_1249),
.Y(n_1452)
);

BUFx4f_ASAP7_75t_SL g1453 ( 
.A(n_1248),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1315),
.A2(n_604),
.B1(n_1050),
.B2(n_761),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_1340),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1340),
.Y(n_1456)
);

INVx4_ASAP7_75t_SL g1457 ( 
.A(n_1419),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1425),
.A2(n_1432),
.B(n_1429),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1417),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1370),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1412),
.A2(n_1416),
.B1(n_1434),
.B2(n_1439),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1339),
.Y(n_1462)
);

AOI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1413),
.A2(n_1415),
.B(n_1449),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1374),
.A2(n_1402),
.B(n_1389),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1408),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1407),
.A2(n_1410),
.B(n_1409),
.Y(n_1466)
);

INVx4_ASAP7_75t_SL g1467 ( 
.A(n_1419),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1339),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1351),
.B(n_1332),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1454),
.A2(n_1434),
.B1(n_1439),
.B2(n_1441),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1351),
.B(n_1332),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1360),
.B(n_1349),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1437),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1344),
.B(n_1342),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1475)
);

AO21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1425),
.A2(n_1429),
.B(n_1443),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1336),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1409),
.A2(n_1392),
.B(n_1404),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1345),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1348),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1426),
.A2(n_1445),
.B(n_1443),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1404),
.B(n_1369),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1341),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1334),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1366),
.B(n_1414),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1392),
.A2(n_1407),
.B(n_1418),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1366),
.B(n_1432),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1433),
.Y(n_1488)
);

AO21x1_ASAP7_75t_L g1489 ( 
.A1(n_1405),
.A2(n_1402),
.B(n_1397),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1405),
.A2(n_1398),
.B(n_1403),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1377),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1377),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1355),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1441),
.B(n_1352),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1363),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1352),
.B(n_1386),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1410),
.A2(n_1418),
.B(n_1420),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1388),
.A2(n_1373),
.B(n_1427),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1442),
.B(n_1371),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1406),
.B(n_1384),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1406),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1420),
.A2(n_1361),
.B(n_1357),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1375),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1380),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1412),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1428),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_1399),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1416),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1431),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_SL g1510 ( 
.A(n_1423),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1386),
.B(n_1369),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1447),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1451),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1364),
.B(n_1394),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1408),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1411),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1361),
.B(n_1357),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1376),
.A2(n_1382),
.B(n_1381),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1422),
.B(n_1448),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1430),
.B(n_1381),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1388),
.Y(n_1521)
);

BUFx8_ASAP7_75t_SL g1522 ( 
.A(n_1353),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1382),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1385),
.A2(n_1393),
.B(n_1395),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1385),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1376),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1390),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1390),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1378),
.B(n_1396),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1426),
.B(n_1362),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1367),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1331),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1359),
.B(n_1387),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1368),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1368),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1400),
.A2(n_1424),
.B(n_1346),
.Y(n_1536)
);

OAI222xp33_ASAP7_75t_L g1537 ( 
.A1(n_1453),
.A2(n_1379),
.B1(n_1438),
.B2(n_1337),
.C1(n_1436),
.C2(n_1350),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1383),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1383),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1536),
.Y(n_1540)
);

A2O1A1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1481),
.A2(n_1335),
.B(n_1333),
.C(n_1452),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1504),
.B(n_1338),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1481),
.A2(n_1333),
.B(n_1452),
.C(n_1446),
.Y(n_1543)
);

NAND4xp25_ASAP7_75t_L g1544 ( 
.A(n_1530),
.B(n_1450),
.C(n_1350),
.D(n_1354),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1524),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1474),
.B(n_1391),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1472),
.A2(n_1401),
.B(n_1343),
.Y(n_1547)
);

AOI211xp5_ASAP7_75t_L g1548 ( 
.A1(n_1530),
.A2(n_1446),
.B(n_1440),
.C(n_1365),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1458),
.A2(n_1440),
.B(n_1356),
.C(n_1358),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1458),
.A2(n_1356),
.B1(n_1453),
.B2(n_1372),
.C(n_1435),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1477),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1479),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1472),
.A2(n_1343),
.B(n_1372),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1470),
.A2(n_1343),
.B1(n_1435),
.B2(n_1461),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1484),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1455),
.B(n_1483),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1469),
.A2(n_1435),
.B(n_1471),
.C(n_1475),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_SL g1558 ( 
.A1(n_1536),
.A2(n_1489),
.B(n_1461),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1459),
.B(n_1514),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1476),
.A2(n_1475),
.B1(n_1469),
.B2(n_1471),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1489),
.A2(n_1502),
.B(n_1486),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1519),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1494),
.A2(n_1496),
.B1(n_1487),
.B2(n_1465),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1499),
.Y(n_1564)
);

BUFx2_ASAP7_75t_R g1565 ( 
.A(n_1522),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1500),
.B(n_1518),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1512),
.B(n_1460),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

AND2x2_ASAP7_75t_SL g1569 ( 
.A(n_1465),
.B(n_1511),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1494),
.A2(n_1526),
.B(n_1462),
.C(n_1468),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1500),
.B(n_1518),
.Y(n_1571)
);

A2O1A1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1487),
.A2(n_1517),
.B(n_1459),
.C(n_1526),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1459),
.B(n_1537),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1524),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1479),
.B(n_1480),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1517),
.A2(n_1511),
.B1(n_1523),
.B2(n_1482),
.C(n_1485),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1485),
.B(n_1515),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1521),
.B(n_1460),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1457),
.B(n_1467),
.Y(n_1582)
);

NAND2x1_ASAP7_75t_L g1583 ( 
.A(n_1507),
.B(n_1501),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1523),
.A2(n_1498),
.B1(n_1516),
.B2(n_1500),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1463),
.A2(n_1497),
.B(n_1482),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_SL g1586 ( 
.A(n_1498),
.B(n_1500),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1493),
.B(n_1495),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1473),
.A2(n_1510),
.B1(n_1516),
.B2(n_1539),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1502),
.A2(n_1486),
.B(n_1497),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1538),
.B(n_1473),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1516),
.A2(n_1505),
.B(n_1508),
.C(n_1466),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1498),
.A2(n_1516),
.B1(n_1529),
.B2(n_1491),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1559),
.B(n_1492),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1573),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1580),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1551),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1501),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1556),
.B(n_1464),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1577),
.A2(n_1476),
.B1(n_1498),
.B2(n_1502),
.Y(n_1603)
);

NAND3xp33_ASAP7_75t_L g1604 ( 
.A(n_1541),
.B(n_1503),
.C(n_1513),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1571),
.B(n_1478),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1506),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1543),
.B(n_1528),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1554),
.A2(n_1502),
.B1(n_1473),
.B2(n_1464),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1464),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1571),
.B(n_1478),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1576),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1545),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1590),
.B(n_1585),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1592),
.B(n_1501),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1585),
.B(n_1478),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1574),
.B(n_1527),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1587),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1575),
.B(n_1456),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1577),
.A2(n_1490),
.B1(n_1509),
.B2(n_1506),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1568),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1587),
.Y(n_1623)
);

OAI33xp33_ASAP7_75t_L g1624 ( 
.A1(n_1620),
.A2(n_1563),
.A3(n_1542),
.B1(n_1570),
.B2(n_1555),
.B3(n_1588),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1561),
.Y(n_1625)
);

INVx3_ASAP7_75t_SL g1626 ( 
.A(n_1616),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1602),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1597),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1561),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1605),
.B(n_1586),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1608),
.A2(n_1572),
.B1(n_1557),
.B2(n_1560),
.C(n_1549),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1597),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1597),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1599),
.B(n_1589),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1540),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1603),
.A2(n_1563),
.B1(n_1584),
.B2(n_1554),
.Y(n_1637)
);

OAI221xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1621),
.A2(n_1548),
.B1(n_1593),
.B2(n_1550),
.C(n_1547),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1604),
.A2(n_1547),
.B(n_1553),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1605),
.B(n_1589),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1603),
.A2(n_1621),
.B1(n_1558),
.B2(n_1608),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1605),
.B(n_1589),
.Y(n_1645)
);

INVx5_ASAP7_75t_SL g1646 ( 
.A(n_1610),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1595),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1610),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1564),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1578),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1599),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1600),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1490),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1636),
.B(n_1613),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1628),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1609),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1652),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1632),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1648),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1649),
.B(n_1654),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1625),
.B(n_1609),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1626),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1651),
.B(n_1595),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1598),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1652),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1634),
.B(n_1598),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1649),
.B(n_1640),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1596),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1625),
.B(n_1606),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1654),
.B(n_1619),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1623),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1650),
.B(n_1611),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1647),
.B(n_1622),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1655),
.B(n_1643),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1675),
.B(n_1635),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1643),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1670),
.Y(n_1690)
);

OAI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1675),
.A2(n_1644),
.B(n_1638),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1657),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1680),
.B(n_1629),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1686),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1618),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1661),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1680),
.B(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1661),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1677),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1659),
.B(n_1643),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1662),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1677),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1659),
.B(n_1645),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1565),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1671),
.B(n_1634),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1666),
.B(n_1645),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1663),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1660),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1660),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1663),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1666),
.B(n_1645),
.Y(n_1716)
);

NAND2x1_ASAP7_75t_L g1717 ( 
.A(n_1679),
.B(n_1627),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1660),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1679),
.A2(n_1638),
.B(n_1641),
.C(n_1631),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1669),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1669),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1671),
.B(n_1630),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1684),
.B(n_1622),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1674),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1671),
.B(n_1634),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1671),
.B(n_1630),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1678),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1697),
.B(n_1665),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1717),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1719),
.B(n_1684),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1710),
.B(n_1673),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1650),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1713),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1658),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1710),
.B(n_1673),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1717),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1692),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1709),
.A2(n_1635),
.B(n_1641),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1692),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1694),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1729),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1690),
.B(n_1658),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1699),
.Y(n_1752)
);

AND2x2_ASAP7_75t_SL g1753 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1689),
.B(n_1685),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1710),
.A2(n_1631),
.B1(n_1637),
.B2(n_1624),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1702),
.B(n_1681),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1693),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1696),
.A2(n_1637),
.B1(n_1653),
.B2(n_1647),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1707),
.B(n_1685),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1689),
.B(n_1679),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1695),
.B(n_1667),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1725),
.B(n_1656),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1699),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1714),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1727),
.B1(n_1710),
.B2(n_1693),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1733),
.B(n_1703),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1742),
.A2(n_1706),
.B(n_1727),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_L g1769 ( 
.A(n_1755),
.B(n_1679),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1730),
.B(n_1703),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1708),
.Y(n_1771)
);

OAI32xp33_ASAP7_75t_L g1772 ( 
.A1(n_1758),
.A2(n_1742),
.A3(n_1732),
.B1(n_1740),
.B2(n_1735),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1757),
.A2(n_1695),
.B(n_1700),
.C(n_1579),
.Y(n_1773)
);

NAND2x1_ASAP7_75t_L g1774 ( 
.A(n_1740),
.B(n_1706),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1732),
.A2(n_1624),
.B(n_1706),
.C(n_1700),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1761),
.B(n_1708),
.Y(n_1776)
);

OAI311xp33_ASAP7_75t_L g1777 ( 
.A1(n_1731),
.A2(n_1550),
.A3(n_1667),
.B1(n_1544),
.C1(n_1553),
.Y(n_1777)
);

OA21x2_ASAP7_75t_L g1778 ( 
.A1(n_1748),
.A2(n_1718),
.B(n_1704),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1748),
.A2(n_1664),
.B1(n_1653),
.B2(n_1648),
.Y(n_1779)
);

NAND4xp25_ASAP7_75t_L g1780 ( 
.A(n_1757),
.B(n_1706),
.C(n_1591),
.D(n_1727),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1764),
.Y(n_1781)
);

AOI21xp33_ASAP7_75t_SL g1782 ( 
.A1(n_1753),
.A2(n_1565),
.B(n_1727),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1731),
.B(n_1757),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1753),
.A2(n_1615),
.B1(n_1617),
.B2(n_1711),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1753),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1757),
.B(n_1711),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1749),
.A2(n_1664),
.B(n_1701),
.Y(n_1787)
);

AOI32xp33_ASAP7_75t_L g1788 ( 
.A1(n_1761),
.A2(n_1728),
.A3(n_1724),
.B1(n_1716),
.B2(n_1615),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1740),
.B(n_1724),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1716),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1741),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1791),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1766),
.A2(n_1740),
.B1(n_1749),
.B2(n_1739),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1770),
.B(n_1743),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1767),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1774),
.Y(n_1796)
);

OAI322xp33_ASAP7_75t_L g1797 ( 
.A1(n_1775),
.A2(n_1738),
.A3(n_1751),
.B1(n_1744),
.B2(n_1741),
.C1(n_1747),
.C2(n_1752),
.Y(n_1797)
);

INVxp33_ASAP7_75t_L g1798 ( 
.A(n_1786),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1776),
.B(n_1736),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1771),
.B(n_1759),
.Y(n_1800)
);

OAI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1772),
.A2(n_1738),
.B(n_1751),
.C(n_1756),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1782),
.A2(n_1744),
.B(n_1746),
.C(n_1752),
.Y(n_1802)
);

AOI222xp33_ASAP7_75t_L g1803 ( 
.A1(n_1769),
.A2(n_1763),
.B1(n_1615),
.B2(n_1739),
.C1(n_1734),
.C2(n_1747),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1768),
.A2(n_1749),
.B1(n_1734),
.B2(n_1739),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1780),
.A2(n_1734),
.B1(n_1739),
.B2(n_1749),
.Y(n_1805)
);

NAND3x2_ASAP7_75t_L g1806 ( 
.A(n_1789),
.B(n_1734),
.C(n_1762),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1778),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1781),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1778),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1789),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1783),
.B(n_1754),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1790),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1807),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1807),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1809),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1810),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1810),
.B(n_1788),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1796),
.Y(n_1818)
);

O2A1O1Ixp33_ASAP7_75t_SL g1819 ( 
.A1(n_1801),
.A2(n_1795),
.B(n_1798),
.C(n_1808),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1795),
.B(n_1736),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1794),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1792),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1797),
.A2(n_1779),
.B1(n_1787),
.B2(n_1777),
.C(n_1746),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1821),
.B(n_1798),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1813),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1813),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1818),
.B(n_1812),
.Y(n_1827)
);

NAND4xp25_ASAP7_75t_L g1828 ( 
.A(n_1823),
.B(n_1805),
.C(n_1793),
.D(n_1804),
.Y(n_1828)
);

NAND2xp33_ASAP7_75t_SL g1829 ( 
.A(n_1820),
.B(n_1816),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1819),
.B(n_1799),
.Y(n_1830)
);

OAI322xp33_ASAP7_75t_L g1831 ( 
.A1(n_1814),
.A2(n_1800),
.A3(n_1811),
.B1(n_1784),
.B2(n_1806),
.C1(n_1802),
.C2(n_1750),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1817),
.Y(n_1832)
);

AOI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1815),
.B1(n_1819),
.B2(n_1822),
.C1(n_1773),
.C2(n_1803),
.Y(n_1833)
);

OAI211xp5_ASAP7_75t_L g1834 ( 
.A1(n_1828),
.A2(n_1815),
.B(n_1777),
.C(n_1765),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1824),
.A2(n_1745),
.B(n_1762),
.C(n_1760),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1830),
.A2(n_1749),
.B1(n_1745),
.B2(n_1760),
.Y(n_1836)
);

AOI211xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1827),
.A2(n_1765),
.B(n_1760),
.C(n_1750),
.Y(n_1837)
);

AOI21xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1833),
.A2(n_1826),
.B(n_1825),
.Y(n_1838)
);

AOI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1834),
.A2(n_1831),
.B1(n_1829),
.B2(n_1765),
.C(n_1750),
.Y(n_1839)
);

AOI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1835),
.A2(n_1737),
.B(n_1728),
.C(n_1546),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1836),
.B(n_1737),
.C(n_1639),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1837),
.A2(n_1737),
.B(n_1718),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1833),
.A2(n_1704),
.B(n_1701),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1840),
.B(n_1726),
.Y(n_1844)
);

NOR2x1_ASAP7_75t_L g1845 ( 
.A(n_1841),
.B(n_1843),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1842),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1838),
.B(n_1705),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_SL g1848 ( 
.A(n_1839),
.B(n_1705),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1845),
.B(n_1712),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1848),
.B(n_1712),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_SL g1851 ( 
.A(n_1847),
.B(n_1639),
.C(n_1627),
.Y(n_1851)
);

XNOR2xp5_ASAP7_75t_L g1852 ( 
.A(n_1851),
.B(n_1846),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1849),
.B1(n_1850),
.B2(n_1844),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1853),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1853),
.A2(n_1720),
.B(n_1715),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1854),
.A2(n_1726),
.B1(n_1723),
.B2(n_1722),
.Y(n_1856)
);

XNOR2x1_ASAP7_75t_L g1857 ( 
.A(n_1855),
.B(n_1507),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1856),
.A2(n_1723),
.B1(n_1722),
.B2(n_1720),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1857),
.B(n_1715),
.Y(n_1859)
);

AO21x2_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1683),
.B(n_1672),
.Y(n_1860)
);

XNOR2xp5_ASAP7_75t_L g1861 ( 
.A(n_1860),
.B(n_1607),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_R g1862 ( 
.A1(n_1861),
.A2(n_1642),
.B1(n_1682),
.B2(n_1646),
.C(n_1648),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1594),
.B(n_1534),
.C(n_1535),
.Y(n_1863)
);


endmodule