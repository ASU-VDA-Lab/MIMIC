module fake_ariane_2111_n_1152 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1152);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1152;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_1133;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_401;
wire n_485;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_770;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_1080;
wire n_920;
wire n_576;
wire n_843;
wire n_899;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1148;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_608;
wire n_892;
wire n_494;
wire n_959;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_856;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_1069;
wire n_393;
wire n_965;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g221 ( 
.A(n_67),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_11),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_213),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_26),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_171),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_86),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_57),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_158),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_120),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_87),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_71),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_7),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_47),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_30),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_127),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_5),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_103),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_179),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_97),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_62),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_202),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_116),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_107),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_184),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_150),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_174),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_146),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_43),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_22),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_110),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_173),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_145),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_162),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_76),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_68),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_101),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_111),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_83),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_23),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_42),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_125),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_190),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_225),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_222),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_227),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_245),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_221),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_237),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_288),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_230),
.Y(n_310)
);

BUFx6f_ASAP7_75t_SL g311 ( 
.A(n_235),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_230),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_277),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_235),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_234),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_233),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_224),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_224),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_259),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_282),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_236),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_286),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_232),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_232),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_280),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_279),
.B(n_278),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_324),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_334),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_319),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_326),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_336),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_264),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_308),
.A2(n_307),
.B1(n_333),
.B2(n_329),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_322),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_271),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_317),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_304),
.Y(n_373)
);

AND3x2_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_271),
.C(n_290),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_283),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_329),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_333),
.B(n_242),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_320),
.A2(n_284),
.B(n_280),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_297),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_295),
.B(n_228),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_298),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_308),
.A2(n_242),
.B1(n_250),
.B2(n_275),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_337),
.A2(n_286),
.B(n_240),
.Y(n_394)
);

NOR2x1_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_266),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

CKINVDCx8_ASAP7_75t_R g398 ( 
.A(n_323),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_344),
.B(n_339),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_343),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_339),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_310),
.Y(n_406)
);

NOR2x1p5_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_323),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_250),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_344),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_349),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_229),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_371),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_285),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_294),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_355),
.B(n_275),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_355),
.B(n_396),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_276),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_276),
.B1(n_311),
.B2(n_238),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

AOI21x1_ASAP7_75t_L g437 ( 
.A1(n_375),
.A2(n_252),
.B(n_251),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_353),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_371),
.B(n_340),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_368),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_340),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_366),
.B(n_253),
.Y(n_450)
);

AND3x2_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_313),
.C(n_310),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_395),
.B(n_391),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_367),
.B(n_254),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_394),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_372),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_373),
.B(n_255),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_372),
.Y(n_471)
);

AO21x2_ASAP7_75t_L g472 ( 
.A1(n_381),
.A2(n_262),
.B(n_256),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_372),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_377),
.B(n_263),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_411),
.B(n_361),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_424),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_313),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_427),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_377),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_400),
.B(n_383),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_437),
.A2(n_386),
.B(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_410),
.B(n_372),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_414),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g493 ( 
.A(n_401),
.B(n_370),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_397),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_420),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_409),
.B(n_362),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_409),
.B(n_362),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_399),
.B(n_348),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_380),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_439),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_420),
.B(n_397),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_365),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_421),
.B(n_474),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

XOR2x2_ASAP7_75t_L g516 ( 
.A(n_406),
.B(n_451),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_436),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_416),
.B(n_348),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_450),
.B(n_380),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_425),
.B(n_398),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_442),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_408),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g525 ( 
.A1(n_430),
.A2(n_386),
.B(n_394),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

BUFx6f_ASAP7_75t_SL g527 ( 
.A(n_446),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_470),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_406),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_380),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_454),
.B(n_446),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_471),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_423),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_454),
.B(n_398),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_454),
.B(n_387),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_469),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_430),
.B(n_397),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_407),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_446),
.B(n_356),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_380),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_402),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_455),
.B(n_380),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_435),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_435),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_446),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_437),
.B(n_397),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_462),
.B(n_374),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_418),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_475),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_484),
.B(n_356),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_356),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_479),
.Y(n_566)
);

INVx8_ASAP7_75t_L g567 ( 
.A(n_527),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_514),
.B(n_445),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_497),
.B(n_423),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_497),
.B(n_394),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_502),
.B(n_462),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_483),
.B(n_351),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_458),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_492),
.B(n_496),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_513),
.A2(n_472),
.B1(n_458),
.B2(n_465),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_498),
.A2(n_501),
.B1(n_521),
.B2(n_499),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_482),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_477),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_536),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_480),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_485),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_547),
.A2(n_462),
.B(n_412),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_486),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_518),
.B(n_472),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_540),
.B(n_462),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_540),
.B(n_462),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_547),
.A2(n_412),
.B(n_405),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_499),
.A2(n_472),
.B1(n_382),
.B2(n_369),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_535),
.B(n_465),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_552),
.A2(n_382),
.B1(n_369),
.B2(n_405),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_478),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_534),
.B(n_465),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_492),
.B(n_496),
.Y(n_594)
);

AND2x6_ASAP7_75t_SL g595 ( 
.A(n_531),
.B(n_0),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_552),
.B(n_415),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_488),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_560),
.B(n_465),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_478),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_537),
.A2(n_351),
.B(n_461),
.C(n_408),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_554),
.A2(n_382),
.B1(n_461),
.B2(n_408),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_534),
.B(n_473),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_529),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_415),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_473),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_541),
.B(n_351),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_490),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_527),
.B(n_369),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_543),
.B(n_473),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_487),
.B(n_473),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_487),
.B(n_473),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_543),
.B(n_402),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_SL g616 ( 
.A(n_522),
.B(n_270),
.C(n_267),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_529),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_500),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_481),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_558),
.B(n_461),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_541),
.B(n_438),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_402),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_511),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_560),
.B(n_402),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_522),
.B(n_438),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_491),
.B(n_503),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_SL g627 ( 
.A1(n_523),
.A2(n_449),
.B(n_438),
.C(n_447),
.Y(n_627)
);

AND2x6_ASAP7_75t_SL g628 ( 
.A(n_516),
.B(n_0),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_481),
.B(n_449),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_476),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_505),
.B(n_449),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_526),
.A2(n_369),
.B1(n_453),
.B2(n_448),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_538),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_617),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_579),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_585),
.B(n_556),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_576),
.B(n_476),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_538),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_SL g640 ( 
.A(n_569),
.B(n_525),
.C(n_519),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_577),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_580),
.B(n_476),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_563),
.Y(n_643)
);

AOI221xp5_ASAP7_75t_L g644 ( 
.A1(n_564),
.A2(n_510),
.B1(n_506),
.B2(n_509),
.C(n_533),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_581),
.B(n_512),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_566),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_592),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_562),
.B(n_545),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_621),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_600),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_582),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_568),
.B(n_545),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_616),
.B(n_605),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_619),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_567),
.A2(n_494),
.B1(n_507),
.B2(n_530),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_SL g659 ( 
.A(n_625),
.B(n_281),
.C(n_274),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_573),
.B(n_508),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_630),
.B(n_523),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_572),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_626),
.B(n_508),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_603),
.B(n_556),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_565),
.B(n_544),
.Y(n_668)
);

AND3x2_ASAP7_75t_SL g669 ( 
.A(n_595),
.B(n_559),
.C(n_447),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_612),
.B(n_545),
.Y(n_670)
);

AND3x1_ASAP7_75t_L g671 ( 
.A(n_610),
.B(n_539),
.C(n_546),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_613),
.B(n_545),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_590),
.B(n_528),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_532),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_623),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_593),
.B(n_604),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_614),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_618),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_599),
.B(n_548),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_628),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_620),
.B(n_550),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_557),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

NAND2x1p5_ASAP7_75t_L g685 ( 
.A(n_596),
.B(n_551),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_597),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_606),
.B(n_561),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_629),
.Y(n_688)
);

AND2x2_ASAP7_75t_SL g689 ( 
.A(n_610),
.B(n_553),
.Y(n_689)
);

AOI21x1_ASAP7_75t_L g690 ( 
.A1(n_602),
.A2(n_489),
.B(n_555),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_629),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_606),
.Y(n_692)
);

BUFx4f_ASAP7_75t_L g693 ( 
.A(n_630),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_589),
.B(n_524),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_624),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_SL g696 ( 
.A(n_571),
.B(n_292),
.C(n_289),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_635),
.B(n_608),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_SL g698 ( 
.A1(n_676),
.A2(n_611),
.B(n_615),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_655),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_647),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_650),
.A2(n_570),
.B(n_611),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_644),
.A2(n_631),
.B(n_601),
.C(n_622),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_690),
.A2(n_583),
.B(n_588),
.Y(n_703)
);

AOI221xp5_ASAP7_75t_SL g704 ( 
.A1(n_644),
.A2(n_602),
.B1(n_632),
.B2(n_520),
.C(n_515),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_693),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_693),
.Y(n_706)
);

NOR2x1_ASAP7_75t_SL g707 ( 
.A(n_638),
.B(n_586),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_SL g708 ( 
.A(n_659),
.B(n_293),
.C(n_607),
.Y(n_708)
);

OAI22x1_ASAP7_75t_L g709 ( 
.A1(n_669),
.A2(n_587),
.B1(n_607),
.B2(n_596),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_634),
.A2(n_627),
.B(n_591),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_637),
.B(n_517),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_654),
.A2(n_448),
.B(n_443),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_666),
.A2(n_460),
.B(n_453),
.C(n_443),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_647),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_660),
.A2(n_460),
.B(n_494),
.Y(n_715)
);

AOI21x1_ASAP7_75t_L g716 ( 
.A1(n_660),
.A2(n_507),
.B(n_494),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_647),
.B(n_494),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_651),
.B(n_369),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_651),
.B(n_369),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_636),
.A2(n_507),
.B1(n_494),
.B2(n_417),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_640),
.A2(n_507),
.B(n_417),
.Y(n_721)
);

AOI21x1_ASAP7_75t_SL g722 ( 
.A1(n_634),
.A2(n_1),
.B(n_2),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_639),
.A2(n_507),
.B(n_417),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_675),
.B(n_667),
.Y(n_725)
);

AO31x2_ASAP7_75t_L g726 ( 
.A1(n_683),
.A2(n_417),
.A3(n_106),
.B(n_108),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_639),
.A2(n_417),
.B(n_35),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_668),
.A2(n_674),
.B(n_673),
.C(n_696),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_665),
.A2(n_37),
.B(n_33),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_665),
.A2(n_40),
.B(n_39),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_689),
.B(n_2),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_687),
.A2(n_44),
.B(n_41),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_687),
.A2(n_46),
.B(n_45),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_673),
.A2(n_3),
.B(n_5),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_643),
.B(n_3),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_646),
.B(n_6),
.Y(n_736)
);

AO31x2_ASAP7_75t_L g737 ( 
.A1(n_683),
.A2(n_684),
.A3(n_686),
.B(n_692),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_645),
.Y(n_738)
);

BUFx6f_ASAP7_75t_SL g739 ( 
.A(n_642),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_670),
.A2(n_50),
.B(n_48),
.Y(n_740)
);

OAI21x1_ASAP7_75t_SL g741 ( 
.A1(n_674),
.A2(n_691),
.B(n_688),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_648),
.B(n_6),
.Y(n_742)
);

AOI21x1_ASAP7_75t_L g743 ( 
.A1(n_672),
.A2(n_52),
.B(n_51),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_695),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_653),
.B(n_9),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_671),
.A2(n_658),
.B(n_685),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_671),
.A2(n_54),
.B(n_53),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_661),
.B(n_10),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_677),
.B(n_10),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_685),
.A2(n_58),
.B(n_55),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_657),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_678),
.B(n_11),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_694),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_633),
.A2(n_60),
.B(n_59),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_633),
.A2(n_130),
.B(n_214),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_641),
.A2(n_129),
.B(n_212),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_642),
.B(n_682),
.Y(n_757)
);

OA22x2_ASAP7_75t_L g758 ( 
.A1(n_669),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_641),
.A2(n_132),
.B(n_211),
.Y(n_759)
);

AO31x2_ASAP7_75t_L g760 ( 
.A1(n_710),
.A2(n_649),
.A3(n_652),
.B(n_656),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_738),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_724),
.Y(n_762)
);

OAI22x1_ASAP7_75t_L g763 ( 
.A1(n_731),
.A2(n_657),
.B1(n_679),
.B2(n_680),
.Y(n_763)
);

AO21x2_ASAP7_75t_L g764 ( 
.A1(n_701),
.A2(n_679),
.B(n_663),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_SL g765 ( 
.A(n_753),
.B(n_681),
.C(n_662),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_SL g766 ( 
.A1(n_744),
.A2(n_663),
.B(n_657),
.C(n_18),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_741),
.Y(n_767)
);

INVx6_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

AO31x2_ASAP7_75t_L g769 ( 
.A1(n_709),
.A2(n_681),
.A3(n_662),
.B(n_663),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_705),
.B(n_663),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_698),
.A2(n_723),
.B(n_727),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_702),
.A2(n_15),
.B(n_17),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_711),
.B(n_15),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_703),
.A2(n_131),
.B(n_210),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_728),
.A2(n_17),
.B(n_18),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_720),
.A2(n_19),
.B(n_20),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_758),
.B(n_19),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_714),
.B(n_20),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_757),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_725),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_720),
.A2(n_21),
.B(n_22),
.Y(n_781)
);

AO31x2_ASAP7_75t_L g782 ( 
.A1(n_746),
.A2(n_135),
.A3(n_209),
.B(n_208),
.Y(n_782)
);

AOI221x1_ASAP7_75t_L g783 ( 
.A1(n_734),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.C(n_25),
.Y(n_783)
);

AOI31xp67_ASAP7_75t_L g784 ( 
.A1(n_722),
.A2(n_217),
.A3(n_134),
.B(n_136),
.Y(n_784)
);

BUFx12f_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_715),
.A2(n_721),
.B(n_716),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_697),
.B(n_24),
.Y(n_787)
);

BUFx12f_ASAP7_75t_L g788 ( 
.A(n_705),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_706),
.B(n_700),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_717),
.A2(n_25),
.B(n_26),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_706),
.B(n_27),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_707),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_704),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

AO31x2_ASAP7_75t_L g795 ( 
.A1(n_713),
.A2(n_140),
.A3(n_206),
.B(n_205),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_750),
.A2(n_133),
.A3(n_204),
.B(n_201),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_732),
.A2(n_28),
.B(n_29),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_735),
.B(n_30),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_751),
.Y(n_799)
);

AO21x2_ASAP7_75t_L g800 ( 
.A1(n_747),
.A2(n_139),
.B(n_200),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_704),
.A2(n_31),
.B(n_32),
.C(n_61),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_708),
.A2(n_32),
.B1(n_63),
.B2(n_64),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_737),
.B(n_65),
.Y(n_804)
);

AO32x2_ASAP7_75t_L g805 ( 
.A1(n_726),
.A2(n_66),
.A3(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_R g806 ( 
.A(n_736),
.B(n_73),
.Y(n_806)
);

OAI22x1_ASAP7_75t_L g807 ( 
.A1(n_742),
.A2(n_745),
.B1(n_748),
.B2(n_749),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_752),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_733),
.A2(n_729),
.B(n_754),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_739),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_718),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_811)
);

AOI31xp67_ASAP7_75t_L g812 ( 
.A1(n_719),
.A2(n_207),
.A3(n_79),
.B(n_80),
.Y(n_812)
);

BUFx10_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_726),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_759),
.B(n_78),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_730),
.A2(n_81),
.B(n_84),
.Y(n_816)
);

NAND3xp33_ASAP7_75t_L g817 ( 
.A(n_726),
.B(n_85),
.C(n_88),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_740),
.A2(n_90),
.A3(n_91),
.B(n_92),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_712),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_756),
.A2(n_755),
.B(n_743),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_725),
.Y(n_821)
);

NOR4xp25_ASAP7_75t_L g822 ( 
.A(n_744),
.B(n_94),
.C(n_95),
.D(n_96),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_698),
.A2(n_199),
.B(n_99),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_753),
.B(n_98),
.C(n_100),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_728),
.A2(n_102),
.B(n_104),
.Y(n_825)
);

BUFx12f_ASAP7_75t_L g826 ( 
.A(n_785),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_105),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_777),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_769),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_SL g830 ( 
.A1(n_775),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_761),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_SL g832 ( 
.A1(n_808),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_779),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_780),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_813),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_788),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_798),
.A2(n_126),
.B1(n_128),
.B2(n_141),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_807),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_825),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_787),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_783),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_799),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_821),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_SL g844 ( 
.A1(n_763),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_772),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_845)
);

INVx6_ASAP7_75t_L g846 ( 
.A(n_794),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_768),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_817),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_789),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_768),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_802),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_824),
.A2(n_168),
.B1(n_170),
.B2(n_172),
.Y(n_852)
);

CKINVDCx14_ASAP7_75t_R g853 ( 
.A(n_794),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_778),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_804),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_778),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_810),
.B(n_175),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_783),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_859)
);

CKINVDCx6p67_ASAP7_75t_R g860 ( 
.A(n_789),
.Y(n_860)
);

CKINVDCx6p67_ASAP7_75t_R g861 ( 
.A(n_770),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_767),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_806),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_773),
.Y(n_864)
);

BUFx2_ASAP7_75t_R g865 ( 
.A(n_764),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_805),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_776),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_781),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_805),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_792),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_791),
.B(n_192),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_SL g873 ( 
.A1(n_790),
.A2(n_193),
.B(n_194),
.Y(n_873)
);

CKINVDCx6p67_ASAP7_75t_R g874 ( 
.A(n_770),
.Y(n_874)
);

INVx6_ASAP7_75t_L g875 ( 
.A(n_769),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_815),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_805),
.A2(n_771),
.B1(n_823),
.B2(n_816),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_811),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_797),
.Y(n_879)
);

BUFx2_ASAP7_75t_SL g880 ( 
.A(n_809),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_875),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_834),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_866),
.B(n_819),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_SL g884 ( 
.A1(n_870),
.A2(n_800),
.B1(n_793),
.B2(n_801),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_831),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_857),
.B(n_766),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_829),
.A2(n_786),
.B(n_820),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_843),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_871),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_855),
.Y(n_890)
);

AO21x2_ASAP7_75t_L g891 ( 
.A1(n_841),
.A2(n_822),
.B(n_765),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_856),
.B(n_782),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_857),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_829),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_864),
.B(n_782),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_862),
.B(n_795),
.Y(n_896)
);

BUFx4f_ASAP7_75t_SL g897 ( 
.A(n_826),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_869),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_875),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_851),
.B(n_795),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_875),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_833),
.B(n_818),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_849),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_880),
.Y(n_904)
);

AO21x2_ASAP7_75t_L g905 ( 
.A1(n_841),
.A2(n_774),
.B(n_784),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_879),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_865),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_827),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_827),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_842),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_877),
.B(n_796),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_849),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_877),
.B(n_796),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_859),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_838),
.A2(n_803),
.B(n_784),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_846),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_859),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_846),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_858),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_846),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_858),
.A2(n_847),
.B(n_835),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_850),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_872),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_860),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_840),
.B(n_812),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_906),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_898),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_885),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_885),
.B(n_853),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_904),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_898),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

OA21x2_ASAP7_75t_L g933 ( 
.A1(n_887),
.A2(n_838),
.B(n_873),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_889),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_898),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_911),
.A2(n_863),
.B(n_812),
.Y(n_936)
);

AO21x2_ASAP7_75t_L g937 ( 
.A1(n_911),
.A2(n_839),
.B(n_848),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_910),
.B(n_853),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_889),
.B(n_836),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_890),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_890),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_883),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_883),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_882),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_910),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_894),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_882),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_918),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_888),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_918),
.Y(n_950)
);

NOR2x1_ASAP7_75t_SL g951 ( 
.A(n_921),
.B(n_854),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_918),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_887),
.A2(n_867),
.B(n_868),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_928),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_926),
.B(n_929),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_926),
.B(n_904),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_932),
.B(n_922),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_940),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_934),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_929),
.B(n_904),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_942),
.B(n_913),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_928),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_946),
.B(n_893),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_940),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_944),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_946),
.B(n_893),
.Y(n_968)
);

OR2x2_ASAP7_75t_SL g969 ( 
.A(n_933),
.B(n_914),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_945),
.B(n_922),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_942),
.B(n_893),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_930),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_930),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_943),
.B(n_893),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_941),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_941),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_927),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_956),
.B(n_953),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_967),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_955),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_963),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_960),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_956),
.B(n_953),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_962),
.B(n_943),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_962),
.B(n_939),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_972),
.A2(n_937),
.B(n_891),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_969),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_958),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_977),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_977),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_957),
.B(n_944),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_982),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_979),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_964),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_985),
.B(n_969),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_980),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_984),
.B(n_964),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_989),
.B(n_971),
.Y(n_999)
);

AND2x2_ASAP7_75t_SL g1000 ( 
.A(n_988),
.B(n_933),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_986),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_981),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_983),
.B(n_968),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_990),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_991),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_994),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1003),
.B(n_987),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_995),
.B(n_968),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_997),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_993),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_996),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1003),
.B(n_987),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1002),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1004),
.B(n_1001),
.Y(n_1014)
);

AO221x2_ASAP7_75t_L g1015 ( 
.A1(n_1014),
.A2(n_999),
.B1(n_938),
.B2(n_897),
.C(n_993),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1010),
.B(n_1000),
.Y(n_1017)
);

OAI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_1007),
.A2(n_996),
.B1(n_914),
.B2(n_917),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_1014),
.B(n_1005),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_1011),
.B(n_995),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1006),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1009),
.B(n_1000),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1021),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_1019),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1017),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_1020),
.Y(n_1026)
);

NOR2x1_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_1013),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1016),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_1015),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1018),
.A2(n_1012),
.B(n_925),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1020),
.B(n_998),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1020),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1020),
.B(n_998),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1027),
.A2(n_1005),
.B(n_917),
.Y(n_1034)
);

XNOR2x1_ASAP7_75t_L g1035 ( 
.A(n_1025),
.B(n_924),
.Y(n_1035)
);

NOR2x1_ASAP7_75t_L g1036 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1030),
.A2(n_937),
.B1(n_913),
.B2(n_936),
.Y(n_1037)
);

OAI221xp5_ASAP7_75t_L g1038 ( 
.A1(n_1025),
.A2(n_886),
.B1(n_907),
.B2(n_828),
.C(n_830),
.Y(n_1038)
);

AOI32xp33_ASAP7_75t_L g1039 ( 
.A1(n_1023),
.A2(n_828),
.A3(n_953),
.B1(n_907),
.B2(n_884),
.Y(n_1039)
);

AOI32xp33_ASAP7_75t_L g1040 ( 
.A1(n_1026),
.A2(n_884),
.A3(n_915),
.B1(n_830),
.B2(n_909),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1031),
.B(n_924),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_971),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_836),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1041),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_SL g1046 ( 
.A1(n_1034),
.A2(n_1024),
.B(n_1028),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1042),
.B(n_1029),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1024),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_1036),
.B(n_837),
.C(n_839),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1037),
.B(n_974),
.Y(n_1050)
);

INVxp33_ASAP7_75t_L g1051 ( 
.A(n_1038),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1039),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_1045),
.A2(n_832),
.B(n_891),
.C(n_837),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1044),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1046),
.A2(n_936),
.B1(n_891),
.B2(n_937),
.C(n_895),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1049),
.A2(n_840),
.B1(n_936),
.B2(n_891),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1053),
.A2(n_936),
.B1(n_908),
.B2(n_909),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1048),
.B(n_992),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1052),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1052),
.A2(n_908),
.B1(n_909),
.B2(n_933),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1050),
.B(n_992),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1059),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1060),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1055),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_1058),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_1062),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1057),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_1054),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1056),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1065),
.A2(n_1047),
.B(n_1051),
.Y(n_1072)
);

NOR3x1_ASAP7_75t_L g1073 ( 
.A(n_1063),
.B(n_939),
.C(n_973),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1064),
.B(n_876),
.C(n_921),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1067),
.B(n_985),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_L g1076 ( 
.A(n_1069),
.B(n_974),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1068),
.B(n_957),
.Y(n_1077)
);

NAND5xp2_ASAP7_75t_L g1078 ( 
.A(n_1071),
.B(n_876),
.C(n_845),
.D(n_852),
.E(n_848),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_973),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_L g1080 ( 
.A(n_1070),
.B(n_961),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1080),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1076),
.B(n_1070),
.Y(n_1082)
);

NOR4xp25_ASAP7_75t_L g1083 ( 
.A(n_1075),
.B(n_1066),
.C(n_868),
.D(n_867),
.Y(n_1083)
);

OAI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_1072),
.A2(n_845),
.B1(n_844),
.B2(n_909),
.C(n_852),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1073),
.A2(n_972),
.B1(n_961),
.B2(n_930),
.C(n_919),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1079),
.A2(n_951),
.B(n_878),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1078),
.B(n_905),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1083),
.B(n_1077),
.Y(n_1088)
);

NAND4xp25_ASAP7_75t_L g1089 ( 
.A(n_1082),
.B(n_1074),
.C(n_919),
.D(n_916),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1081),
.B(n_923),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_1086),
.B(n_1084),
.C(n_1087),
.Y(n_1091)
);

OAI211xp5_ASAP7_75t_L g1092 ( 
.A1(n_1085),
.A2(n_933),
.B(n_930),
.C(n_915),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1082),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_SL g1094 ( 
.A(n_1082),
.B(n_951),
.C(n_923),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1082),
.A2(n_905),
.B(n_923),
.C(n_895),
.Y(n_1095)
);

AOI221x1_ASAP7_75t_L g1096 ( 
.A1(n_1081),
.A2(n_916),
.B1(n_920),
.B2(n_947),
.C(n_949),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1088),
.B(n_1093),
.C(n_1090),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1089),
.Y(n_1098)
);

NOR2x1p5_ASAP7_75t_L g1099 ( 
.A(n_1091),
.B(n_861),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1094),
.Y(n_1100)
);

NOR2x1p5_ASAP7_75t_L g1101 ( 
.A(n_1092),
.B(n_874),
.Y(n_1101)
);

NOR2x1_ASAP7_75t_L g1102 ( 
.A(n_1095),
.B(n_905),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_1096),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1091),
.A2(n_905),
.B1(n_915),
.B2(n_975),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1093),
.B(n_916),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1088),
.Y(n_1106)
);

AND3x4_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_903),
.C(n_912),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1106),
.B(n_976),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1103),
.Y(n_1109)
);

AND4x1_ASAP7_75t_L g1110 ( 
.A(n_1098),
.B(n_899),
.C(n_901),
.D(n_949),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1099),
.Y(n_1111)
);

XOR2x2_ASAP7_75t_L g1112 ( 
.A(n_1097),
.B(n_903),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1101),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1100),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1102),
.B(n_1104),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1097),
.B(n_976),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_1097),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_L g1118 ( 
.A(n_1106),
.B(n_903),
.C(n_912),
.D(n_916),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_SL g1119 ( 
.A(n_1106),
.B(n_975),
.C(n_966),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_1117),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1109),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1114),
.B(n_912),
.Y(n_1122)
);

NAND4xp25_ASAP7_75t_L g1123 ( 
.A(n_1116),
.B(n_920),
.C(n_894),
.D(n_881),
.Y(n_1123)
);

NAND5xp2_ASAP7_75t_L g1124 ( 
.A(n_1108),
.B(n_901),
.C(n_899),
.D(n_818),
.E(n_947),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1112),
.Y(n_1125)
);

NAND4xp25_ASAP7_75t_L g1126 ( 
.A(n_1113),
.B(n_920),
.C(n_881),
.D(n_896),
.Y(n_1126)
);

XOR2xp5_ASAP7_75t_L g1127 ( 
.A(n_1111),
.B(n_892),
.Y(n_1127)
);

NOR2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1118),
.B(n_881),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_1121),
.A2(n_1115),
.B1(n_1107),
.B2(n_1119),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_1120),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1122),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_L g1132 ( 
.A1(n_1125),
.A2(n_1110),
.B1(n_952),
.B2(n_950),
.Y(n_1132)
);

AO22x2_ASAP7_75t_L g1133 ( 
.A1(n_1127),
.A2(n_966),
.B1(n_965),
.B2(n_959),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1128),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1124),
.A2(n_948),
.B1(n_965),
.B2(n_959),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1123),
.Y(n_1136)
);

XNOR2xp5_ASAP7_75t_L g1137 ( 
.A(n_1129),
.B(n_1126),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1130),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1131),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1138),
.B(n_1134),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1140),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1141),
.B(n_1139),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1142),
.A2(n_1137),
.B1(n_1136),
.B2(n_1132),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_1135),
.B1(n_1133),
.B2(n_954),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1142),
.A2(n_881),
.B1(n_888),
.B2(n_927),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1143),
.B(n_931),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_954),
.B(n_892),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1145),
.B(n_902),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_902),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1148),
.B(n_935),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_1147),
.B1(n_935),
.B2(n_927),
.Y(n_1151)
);

AOI211xp5_ASAP7_75t_L g1152 ( 
.A1(n_1151),
.A2(n_1149),
.B(n_896),
.C(n_900),
.Y(n_1152)
);


endmodule