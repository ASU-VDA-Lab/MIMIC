module fake_ariane_2203_n_1990 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1990);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1990;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g196 ( 
.A(n_16),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx4_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_130),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

INVx4_ASAP7_75t_R g205 ( 
.A(n_122),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_9),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_29),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_109),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_126),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_18),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_29),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_90),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_0),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_20),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_19),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_124),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_159),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_33),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_151),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_123),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_25),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_73),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_35),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_186),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_161),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_88),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_71),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_83),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_79),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_108),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_34),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_74),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_114),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_32),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_82),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_61),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_38),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_78),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_157),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_187),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_80),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_35),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_24),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_16),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_107),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_24),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_160),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_117),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_168),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_62),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_101),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_96),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_98),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_60),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_191),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_145),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_173),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_19),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_125),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_44),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_110),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_0),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_62),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_25),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_193),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_167),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_111),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_75),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_69),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_85),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_118),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_22),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_77),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_97),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_51),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_94),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_28),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_169),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_147),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_7),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_52),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_32),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_165),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_43),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_150),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_103),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_23),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_128),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_153),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_182),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_93),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_142),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_59),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_41),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_7),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_5),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_45),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_84),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_76),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_10),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_105),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_154),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_170),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_65),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_44),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_8),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_104),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_61),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_21),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_57),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_30),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_50),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_86),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_58),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_81),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_158),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_91),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_131),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_49),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_40),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_64),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_195),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_21),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_11),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_45),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_8),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_140),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_27),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_59),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_171),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_20),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_127),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_2),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_42),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_192),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_64),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_113),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_11),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_95),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_15),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_47),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_9),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_46),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_52),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_1),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_26),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_51),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_56),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_143),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_100),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_27),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_68),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_132),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_175),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_17),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_115),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_37),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_149),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_141),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_33),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_181),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_112),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_232),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_209),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_310),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_334),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_330),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_215),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_207),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_207),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_207),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_310),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_207),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_280),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_284),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_294),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_310),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_298),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_207),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_206),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_306),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_302),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_306),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_306),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_306),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_206),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_306),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_216),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_196),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_198),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_225),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_226),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_234),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_253),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_261),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_290),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_337),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_296),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_309),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_210),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_398),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_398),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_216),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_316),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_348),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_224),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_361),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_362),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_284),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_398),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_373),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_250),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_349),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_236),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_201),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_349),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_201),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_230),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_270),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_230),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_269),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_218),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_383),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_236),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_202),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_204),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_202),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_204),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_304),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_248),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_248),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_332),
.Y(n_493)
);

BUFx2_ASAP7_75t_SL g494 ( 
.A(n_222),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_203),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_351),
.Y(n_496)
);

INVxp33_ASAP7_75t_SL g497 ( 
.A(n_218),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_270),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_299),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_356),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_366),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_203),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_299),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_347),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_471),
.B(n_231),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_SL g509 ( 
.A(n_403),
.B(n_219),
.Y(n_509)
);

BUFx8_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_222),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_389),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_450),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_405),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_389),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_437),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_197),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_308),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_406),
.A2(n_211),
.B(n_199),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_308),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_458),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_214),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_418),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_409),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_410),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_414),
.B(n_220),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_466),
.A2(n_368),
.B1(n_394),
.B2(n_479),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_490),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_468),
.B(n_347),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_493),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_429),
.B(n_221),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_472),
.B(n_347),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_419),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_408),
.B(n_227),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_470),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_403),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_471),
.B(n_474),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_400),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_237),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_395),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_426),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_475),
.B(n_219),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_404),
.B(n_417),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_404),
.B(n_244),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_411),
.A2(n_254),
.B(n_252),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_421),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_428),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_395),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_417),
.B(n_266),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_478),
.B(n_223),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_422),
.B(n_272),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_496),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_425),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_423),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_422),
.B(n_275),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_430),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_430),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_432),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_432),
.Y(n_583)
);

AOI22x1_ASAP7_75t_SL g584 ( 
.A1(n_500),
.A2(n_363),
.B1(n_397),
.B2(n_223),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_427),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_447),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_559),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_557),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_505),
.B(n_474),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_512),
.B(n_514),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_557),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_532),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_559),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_512),
.B(n_451),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_512),
.B(n_451),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_506),
.B(n_412),
.C(n_485),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_530),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_506),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_511),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_552),
.B(n_485),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_566),
.B(n_571),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_537),
.B(n_420),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_534),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_531),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_534),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_512),
.B(n_452),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_565),
.B(n_488),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_537),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_488),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_542),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_541),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_511),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_542),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_546),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_543),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_577),
.B(n_495),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_509),
.A2(n_327),
.B1(n_497),
.B2(n_346),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_513),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_543),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_551),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_516),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_551),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_546),
.B(n_456),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_401),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_510),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_495),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_585),
.Y(n_634)
);

CKINVDCx6p67_ASAP7_75t_R g635 ( 
.A(n_515),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_502),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_579),
.B(n_502),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_519),
.B(n_452),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_563),
.B(n_462),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_517),
.A2(n_491),
.B(n_489),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_522),
.B(n_461),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_517),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_553),
.B(n_431),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_519),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_519),
.B(n_462),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_518),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_518),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_564),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_524),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_524),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_526),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_SL g659 ( 
.A1(n_572),
.A2(n_497),
.B(n_504),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_526),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_529),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_580),
.A2(n_327),
.B1(n_561),
.B2(n_525),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_525),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_529),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_581),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_510),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_578),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_578),
.Y(n_668)
);

AOI21x1_ASAP7_75t_L g669 ( 
.A1(n_523),
.A2(n_492),
.B(n_491),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_532),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_582),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_582),
.B(n_492),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_507),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_519),
.B(n_499),
.Y(n_675)
);

AND2x2_ASAP7_75t_SL g676 ( 
.A(n_558),
.B(n_236),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_583),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_507),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_510),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_508),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_583),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_513),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_508),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_520),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_579),
.B(n_481),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_513),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_575),
.A2(n_239),
.B1(n_480),
.B2(n_433),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_544),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_555),
.A2(n_370),
.B1(n_375),
.B2(n_363),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_545),
.B(n_499),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_523),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_572),
.B(n_208),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_520),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_547),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_563),
.B(n_208),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_510),
.B(n_212),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_560),
.B(n_503),
.Y(n_697)
);

INVx8_ASAP7_75t_L g698 ( 
.A(n_522),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_522),
.B(n_212),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_522),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_525),
.B(n_482),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_550),
.A2(n_375),
.B1(n_377),
.B2(n_370),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_547),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_548),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_525),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_550),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_548),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_561),
.B(n_570),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_538),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_538),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_561),
.B(n_439),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_538),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_544),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_561),
.B(n_213),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_570),
.B(n_213),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_544),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_544),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_570),
.Y(n_721)
);

AOI21x1_ASAP7_75t_L g722 ( 
.A1(n_567),
.A2(n_503),
.B(n_435),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_549),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_584),
.A2(n_379),
.B1(n_382),
.B2(n_377),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_567),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_549),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_586),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_549),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_568),
.B(n_217),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_584),
.A2(n_486),
.B1(n_483),
.B2(n_441),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_549),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_554),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_554),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_568),
.B(n_217),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_576),
.B(n_228),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_554),
.B(n_440),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_554),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_535),
.A2(n_382),
.B1(n_388),
.B2(n_379),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_590),
.B(n_228),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_659),
.B(n_397),
.C(n_388),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_634),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_602),
.B(n_233),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_650),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_676),
.B(n_229),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_676),
.A2(n_443),
.B1(n_445),
.B2(n_442),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_659),
.A2(n_459),
.B(n_476),
.C(n_473),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_604),
.B(n_576),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_650),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_599),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_621),
.A2(n_341),
.B1(n_293),
.B2(n_295),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_598),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_611),
.B(n_229),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_636),
.B(n_633),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_598),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_630),
.B(n_245),
.C(n_235),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_676),
.A2(n_372),
.B1(n_364),
.B2(n_367),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_611),
.B(n_249),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_618),
.B(n_303),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_600),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_654),
.B(n_303),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_654),
.B(n_364),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_654),
.B(n_367),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_600),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_711),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_601),
.A2(n_446),
.B(n_469),
.C(n_467),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_592),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_716),
.A2(n_448),
.B1(n_449),
.B2(n_465),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_594),
.B(n_256),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_596),
.B(n_257),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_618),
.B(n_369),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_608),
.B(n_369),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_616),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_663),
.B(n_267),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_603),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_656),
.B(n_374),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_663),
.B(n_289),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_663),
.B(n_324),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_616),
.A2(n_277),
.B(n_276),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_711),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_605),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_629),
.B(n_586),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_629),
.B(n_685),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_656),
.B(n_374),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_691),
.B(n_236),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_597),
.A2(n_376),
.B1(n_386),
.B2(n_387),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_620),
.B(n_259),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_663),
.B(n_387),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_656),
.B(n_391),
.Y(n_793)
);

NAND2x1_ASAP7_75t_L g794 ( 
.A(n_664),
.B(n_200),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_605),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_700),
.B(n_391),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_727),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_664),
.B(n_587),
.Y(n_798)
);

OAI221xp5_ASAP7_75t_L g799 ( 
.A1(n_621),
.A2(n_318),
.B1(n_273),
.B2(n_271),
.C(n_268),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_610),
.B(n_260),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_626),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_662),
.B(n_646),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_607),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_685),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_700),
.B(n_396),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_631),
.B(n_454),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_716),
.B(n_399),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_664),
.B(n_399),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_626),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_638),
.B(n_279),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_635),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_662),
.B(n_283),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_685),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_645),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_607),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_685),
.B(n_501),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_685),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_646),
.B(n_639),
.Y(n_819)
);

AND2x6_ASAP7_75t_SL g820 ( 
.A(n_592),
.B(n_455),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_613),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_646),
.B(n_292),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_671),
.B(n_536),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_698),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_597),
.A2(n_278),
.B(n_288),
.C(n_339),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_646),
.B(n_297),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_705),
.B(n_311),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_647),
.B(n_314),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_695),
.B(n_315),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_613),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_617),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_705),
.B(n_321),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_637),
.B(n_329),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_721),
.B(n_331),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_640),
.B(n_614),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_614),
.B(n_721),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_644),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_617),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_587),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_619),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_702),
.B(n_336),
.C(n_335),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_619),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_589),
.B(n_340),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_624),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_690),
.B(n_342),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_614),
.B(n_345),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_631),
.B(n_540),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_692),
.A2(n_307),
.B1(n_313),
.B2(n_319),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_644),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_666),
.B(n_457),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_643),
.B(n_574),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_649),
.Y(n_852)
);

BUFx5_ASAP7_75t_L g853 ( 
.A(n_691),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_614),
.B(n_357),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_587),
.B(n_352),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_624),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_697),
.B(n_360),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_625),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_625),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_708),
.B(n_238),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_587),
.B(n_240),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_593),
.B(n_241),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_671),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_593),
.B(n_390),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_606),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_628),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_628),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_649),
.A2(n_463),
.B1(n_460),
.B2(n_464),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_593),
.B(n_242),
.Y(n_869)
);

INVx8_ASAP7_75t_L g870 ( 
.A(n_698),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_593),
.B(n_243),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_699),
.B(n_393),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_643),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_729),
.B(n_434),
.C(n_435),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_735),
.B(n_434),
.C(n_265),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_658),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_725),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_698),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_712),
.B(n_246),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_666),
.B(n_2),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_247),
.Y(n_881)
);

AOI22x1_ASAP7_75t_L g882 ( 
.A1(n_658),
.A2(n_556),
.B1(n_554),
.B2(n_312),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_679),
.B(n_236),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_588),
.B(n_251),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_632),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_588),
.B(n_255),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_612),
.A2(n_701),
.B1(n_698),
.B2(n_715),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_660),
.B(n_258),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_632),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_591),
.B(n_262),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_660),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_661),
.B(n_263),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_648),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_661),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_591),
.B(n_264),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_648),
.Y(n_896)
);

NOR2xp67_ASAP7_75t_L g897 ( 
.A(n_645),
.B(n_696),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_651),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_706),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_706),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_651),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_595),
.B(n_274),
.Y(n_902)
);

NAND2x1_ASAP7_75t_L g903 ( 
.A(n_622),
.B(n_205),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_653),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_674),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_675),
.B(n_281),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_674),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_653),
.A2(n_484),
.B1(n_325),
.B2(n_359),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_750),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_751),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_814),
.B(n_679),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_755),
.B(n_736),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_743),
.B(n_717),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_741),
.A2(n_739),
.B1(n_730),
.B2(n_657),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_768),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_743),
.B(n_701),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_753),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_846),
.B(n_701),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_835),
.A2(n_668),
.B(n_681),
.C(n_672),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_846),
.B(n_701),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_823),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_804),
.B(n_701),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_804),
.B(n_673),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_854),
.B(n_655),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_818),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_854),
.B(n_772),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_766),
.B(n_655),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_766),
.B(n_725),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_756),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_765),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_772),
.B(n_657),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_773),
.B(n_667),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_742),
.Y(n_933)
);

OR2x2_ASAP7_75t_SL g934 ( 
.A(n_752),
.B(n_739),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_761),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_778),
.A2(n_681),
.B1(n_677),
.B2(n_672),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_870),
.B(n_730),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_784),
.Y(n_938)
);

AND2x4_ASAP7_75t_SL g939 ( 
.A(n_806),
.B(n_615),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_773),
.B(n_668),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_795),
.A2(n_677),
.B1(n_710),
.B2(n_713),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_836),
.B(n_710),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_873),
.B(n_835),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_767),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_776),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_766),
.B(n_622),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_823),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_824),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_803),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_818),
.B(n_673),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_824),
.B(n_622),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_783),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_816),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_821),
.Y(n_954)
);

BUFx8_ASAP7_75t_L g955 ( 
.A(n_770),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_787),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_845),
.B(n_665),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_830),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_831),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_786),
.B(n_615),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_838),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_863),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_801),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_798),
.A2(n_688),
.B(n_622),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_899),
.Y(n_965)
);

NAND2x1p5_ASAP7_75t_L g966 ( 
.A(n_824),
.B(n_709),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_824),
.B(n_641),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_741),
.A2(n_709),
.B(n_665),
.C(n_670),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_746),
.A2(n_745),
.B1(n_752),
.B2(n_841),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_857),
.B(n_670),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_878),
.B(n_641),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_810),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_851),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_746),
.B(n_737),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_840),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_878),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_842),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_844),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_856),
.B(n_704),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_858),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_812),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_859),
.B(n_704),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_820),
.Y(n_983)
);

CKINVDCx14_ASAP7_75t_R g984 ( 
.A(n_817),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_866),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_867),
.B(n_707),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_900),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_878),
.B(n_615),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_798),
.A2(n_686),
.B(n_682),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_878),
.B(n_641),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_870),
.Y(n_991)
);

OAI22xp33_ASAP7_75t_L g992 ( 
.A1(n_758),
.A2(n_799),
.B1(n_848),
.B2(n_887),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_748),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_885),
.B(n_889),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_806),
.B(n_623),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_762),
.A2(n_686),
.B(n_682),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_853),
.B(n_877),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_870),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_837),
.Y(n_999)
);

CKINVDCx8_ASAP7_75t_R g1000 ( 
.A(n_806),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_853),
.B(n_877),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_839),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_815),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_850),
.B(n_623),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_893),
.B(n_896),
.Y(n_1005)
);

INVx4_ASAP7_75t_SL g1006 ( 
.A(n_789),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_898),
.B(n_707),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_762),
.A2(n_686),
.B(n_682),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_901),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_745),
.A2(n_730),
.B1(n_687),
.B2(n_724),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_785),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_850),
.B(n_689),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_904),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_678),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_763),
.A2(n_788),
.B(n_764),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_849),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_852),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_759),
.B(n_680),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_880),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_839),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_883),
.B(n_623),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_891),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_777),
.B(n_680),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_780),
.B(n_683),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_894),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_905),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_744),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_797),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_791),
.A2(n_731),
.B(n_726),
.C(n_733),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_781),
.B(n_683),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_749),
.B(n_684),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_841),
.A2(n_730),
.B1(n_724),
.B2(n_627),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_880),
.B(n_627),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_808),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_883),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_763),
.A2(n_641),
.B(n_682),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_879),
.B(n_684),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_881),
.B(n_693),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_897),
.B(n_802),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_907),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_794),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_769),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_771),
.B(n_693),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_791),
.A2(n_627),
.B1(n_652),
.B2(n_733),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_807),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_827),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_865),
.B(n_694),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_855),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_764),
.A2(n_686),
.B(n_688),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_809),
.A2(n_792),
.B1(n_788),
.B2(n_800),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_771),
.B(n_694),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_832),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_834),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_864),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_800),
.A2(n_829),
.B1(n_793),
.B2(n_779),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_796),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_829),
.A2(n_652),
.B1(n_726),
.B2(n_731),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_SL g1059 ( 
.A1(n_847),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_703),
.Y(n_1060)
);

XNOR2xp5_ASAP7_75t_L g1061 ( 
.A(n_813),
.B(n_757),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_740),
.B(n_703),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_789),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_833),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_789),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_805),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_754),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_789),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_843),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_903),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_864),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_853),
.B(n_609),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_890),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_747),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_819),
.B(n_652),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_895),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_906),
.B(n_728),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_SL g1078 ( 
.A1(n_875),
.A2(n_738),
.B(n_734),
.C(n_732),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_789),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_902),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_790),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_884),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_825),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_775),
.B(n_728),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_886),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_782),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_828),
.B(n_718),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_868),
.B(n_718),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_868),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_811),
.A2(n_353),
.B1(n_291),
.B2(n_300),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_875),
.B(n_719),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_822),
.B(n_642),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_861),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_931),
.A2(n_862),
.B(n_869),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_932),
.A2(n_871),
.B(n_877),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_952),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_913),
.A2(n_874),
.B(n_826),
.C(n_888),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_962),
.B(n_760),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_917),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_912),
.B(n_774),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_912),
.B(n_908),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_955),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_991),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_913),
.B(n_908),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_956),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_926),
.A2(n_874),
.B(n_892),
.C(n_888),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_SL g1107 ( 
.A(n_987),
.B(n_892),
.C(n_355),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_940),
.A2(n_877),
.B(n_853),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_929),
.Y(n_1109)
);

BUFx4f_ASAP7_75t_L g1110 ( 
.A(n_947),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1056),
.A2(n_732),
.B(n_719),
.C(n_738),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_916),
.A2(n_734),
.B(n_723),
.C(n_720),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_930),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_924),
.A2(n_720),
.B(n_723),
.C(n_5),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_909),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_965),
.B(n_642),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_SL g1117 ( 
.A(n_921),
.B(n_1011),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_918),
.B(n_877),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_920),
.B(n_609),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_609),
.B(n_714),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1051),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_955),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_SL g1123 ( 
.A(n_1081),
.B(n_969),
.C(n_1059),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_997),
.A2(n_609),
.B(n_714),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_948),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_938),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_910),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1003),
.A2(n_722),
.B1(n_669),
.B2(n_287),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_943),
.B(n_609),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1001),
.A2(n_714),
.B(n_882),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_948),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_981),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_922),
.B(n_669),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_949),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1059),
.B(n_714),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_969),
.A2(n_714),
.B(n_338),
.C(n_333),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1001),
.A2(n_326),
.B(n_305),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_915),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1020),
.B(n_484),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_983),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_943),
.A2(n_343),
.B(n_317),
.C(n_354),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_SL g1143 ( 
.A1(n_994),
.A2(n_6),
.B(n_12),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1012),
.B(n_1003),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1005),
.A2(n_301),
.B1(n_320),
.B2(n_322),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_L g1146 ( 
.A(n_1047),
.B(n_556),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_993),
.B(n_12),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1046),
.B(n_13),
.Y(n_1148)
);

INVx4_ASAP7_75t_SL g1149 ( 
.A(n_937),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1057),
.B(n_14),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_934),
.B(n_323),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_952),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_953),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_944),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_922),
.B(n_15),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1057),
.B(n_17),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1020),
.B(n_22),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_915),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1072),
.A2(n_350),
.B(n_344),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1054),
.B(n_23),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1035),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_954),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1072),
.A2(n_556),
.B(n_484),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_973),
.B(n_26),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_942),
.A2(n_556),
.B(n_484),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1000),
.B(n_30),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1029),
.B(n_31),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1015),
.A2(n_556),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1066),
.B(n_31),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1010),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_958),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_995),
.B(n_48),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_925),
.B(n_49),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_991),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_925),
.B(n_1074),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_959),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1082),
.B(n_50),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1085),
.B(n_53),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1064),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_933),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_945),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_948),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_911),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1015),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_992),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_995),
.B(n_60),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_933),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_948),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_960),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_963),
.Y(n_1190)
);

NOR3xp33_ASAP7_75t_L g1191 ( 
.A(n_992),
.B(n_63),
.C(n_65),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_976),
.B(n_70),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_961),
.B(n_72),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_960),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_R g1195 ( 
.A(n_984),
.B(n_87),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_975),
.B(n_89),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_SL g1197 ( 
.A(n_1069),
.B(n_120),
.C(n_121),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_977),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_972),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_968),
.A2(n_135),
.B(n_136),
.C(n_139),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_SL g1201 ( 
.A(n_914),
.B(n_144),
.C(n_156),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_978),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_980),
.B(n_174),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_985),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1009),
.B(n_1013),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1053),
.B(n_176),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1076),
.A2(n_179),
.B(n_180),
.C(n_188),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1004),
.B(n_194),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1016),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_914),
.A2(n_1010),
.B1(n_1083),
.B2(n_936),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1036),
.A2(n_1089),
.B1(n_937),
.B2(n_1018),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_919),
.A2(n_1007),
.B1(n_986),
.B2(n_982),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1004),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_979),
.A2(n_974),
.B1(n_941),
.B2(n_1043),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1073),
.B(n_1080),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_988),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1077),
.A2(n_928),
.B(n_957),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_923),
.A2(n_950),
.B1(n_1033),
.B2(n_1067),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1030),
.B(n_970),
.C(n_1093),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_928),
.A2(n_1060),
.B(n_989),
.Y(n_1220)
);

AND2x6_ASAP7_75t_L g1221 ( 
.A(n_1079),
.B(n_976),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_923),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1061),
.A2(n_1040),
.B1(n_1067),
.B2(n_1022),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_998),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1017),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1034),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_950),
.B(n_1034),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1040),
.B(n_1019),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_999),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1055),
.A2(n_1071),
.B(n_1039),
.C(n_1038),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_998),
.Y(n_1231)
);

AND2x2_ASAP7_75t_SL g1232 ( 
.A(n_1068),
.B(n_1079),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_927),
.A2(n_1068),
.B1(n_1022),
.B2(n_1052),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1023),
.Y(n_1234)
);

OA22x2_ASAP7_75t_L g1235 ( 
.A1(n_937),
.A2(n_1028),
.B1(n_939),
.B2(n_1049),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_988),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1002),
.B(n_1021),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_946),
.A2(n_990),
.B(n_951),
.C(n_971),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1048),
.B(n_1002),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1026),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1027),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_964),
.A2(n_989),
.B(n_1050),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_964),
.A2(n_1050),
.B(n_1008),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1091),
.A2(n_1092),
.B(n_1086),
.C(n_1037),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_927),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1044),
.A2(n_1014),
.B1(n_1021),
.B2(n_1084),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1058),
.A2(n_1041),
.B1(n_1045),
.B2(n_1075),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1042),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_996),
.A2(n_1037),
.B(n_1008),
.C(n_1062),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1024),
.B(n_1031),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1108),
.A2(n_1095),
.B(n_1094),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1216),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1105),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1212),
.A2(n_946),
.B(n_951),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1144),
.B(n_1090),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1099),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1102),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1242),
.A2(n_996),
.B(n_1070),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1243),
.A2(n_1070),
.B(n_1042),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_1219),
.B(n_1063),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1123),
.B(n_1087),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1214),
.A2(n_967),
.B(n_971),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1132),
.Y(n_1263)
);

AOI31xp67_ASAP7_75t_L g1264 ( 
.A1(n_1119),
.A2(n_967),
.A3(n_990),
.B(n_1025),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1170),
.A2(n_1088),
.B1(n_1032),
.B2(n_1079),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1104),
.A2(n_1078),
.B(n_966),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1096),
.B(n_966),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1101),
.A2(n_1078),
.B(n_1075),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_1219),
.B(n_1063),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1214),
.A2(n_1063),
.B(n_1065),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1161),
.B(n_1079),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1170),
.A2(n_1063),
.B1(n_1065),
.B2(n_1006),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1110),
.B(n_1065),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1220),
.A2(n_1006),
.B(n_1065),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1152),
.B(n_1183),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1130),
.A2(n_1006),
.B(n_1165),
.Y(n_1276)
);

NAND3x1_ASAP7_75t_L g1277 ( 
.A(n_1151),
.B(n_1166),
.C(n_1191),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1216),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1100),
.A2(n_1210),
.B(n_1143),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1120),
.A2(n_1124),
.B(n_1163),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1116),
.B(n_1155),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1180),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1109),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1244),
.A2(n_1249),
.A3(n_1246),
.B(n_1247),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1158),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1217),
.A2(n_1238),
.B(n_1233),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1183),
.B(n_1175),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1222),
.B(n_1187),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1106),
.A2(n_1246),
.B(n_1137),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1097),
.A2(n_1111),
.B(n_1112),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1213),
.B(n_1226),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1210),
.A2(n_1142),
.B1(n_1205),
.B2(n_1110),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1230),
.A2(n_1233),
.A3(n_1168),
.B(n_1200),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1139),
.B(n_1232),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1113),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1118),
.A2(n_1129),
.B(n_1250),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1223),
.A2(n_1196),
.A3(n_1203),
.B(n_1193),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1215),
.B(n_1239),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1126),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1184),
.A2(n_1201),
.B1(n_1171),
.B2(n_1228),
.C(n_1207),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1209),
.A2(n_1225),
.A3(n_1234),
.B(n_1190),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1134),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1155),
.B(n_1153),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1149),
.B(n_1189),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1237),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1216),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1179),
.B(n_1227),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1162),
.B(n_1176),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1198),
.B(n_1202),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1195),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1127),
.A2(n_1154),
.A3(n_1229),
.B(n_1199),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1178),
.B(n_1169),
.Y(n_1312)
);

NOR2xp67_ASAP7_75t_L g1313 ( 
.A(n_1103),
.B(n_1174),
.Y(n_1313)
);

NAND3xp33_ASAP7_75t_L g1314 ( 
.A(n_1121),
.B(n_1185),
.C(n_1143),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1235),
.A2(n_1218),
.B1(n_1211),
.B2(n_1240),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1171),
.A2(n_1177),
.B(n_1160),
.C(n_1148),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1204),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1218),
.B(n_1173),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1150),
.B(n_1156),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1192),
.A2(n_1135),
.B(n_1146),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1167),
.A2(n_1164),
.B(n_1114),
.C(n_1145),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1172),
.B(n_1186),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1159),
.A2(n_1245),
.B(n_1138),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1189),
.B(n_1194),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1208),
.B(n_1186),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1107),
.A2(n_1098),
.B(n_1206),
.C(n_1208),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1192),
.A2(n_1231),
.B(n_1224),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_SL g1328 ( 
.A(n_1147),
.B(n_1197),
.C(n_1117),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1236),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1224),
.A2(n_1231),
.B(n_1174),
.Y(n_1330)
);

AOI21xp33_ASAP7_75t_L g1331 ( 
.A1(n_1136),
.A2(n_1181),
.B(n_1241),
.Y(n_1331)
);

AOI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1172),
.A2(n_1122),
.B1(n_1157),
.B2(n_1248),
.C(n_1194),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1157),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1133),
.A2(n_1140),
.B(n_1103),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1221),
.A2(n_1125),
.B(n_1131),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1125),
.B(n_1131),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1189),
.B(n_1194),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1236),
.B(n_1149),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1221),
.A2(n_1125),
.B(n_1131),
.Y(n_1339)
);

INVxp67_ASAP7_75t_SL g1340 ( 
.A(n_1182),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1182),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1221),
.A2(n_1182),
.B(n_1188),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1236),
.B(n_1188),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1140),
.Y(n_1344)
);

NAND3x1_ASAP7_75t_L g1345 ( 
.A(n_1141),
.B(n_1221),
.C(n_1140),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1099),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1144),
.B(n_743),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1152),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1104),
.A2(n_755),
.B1(n_926),
.B2(n_743),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1102),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1151),
.A2(n_913),
.B(n_926),
.C(n_755),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1099),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1099),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1108),
.A2(n_1001),
.B(n_997),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1104),
.B(n_926),
.Y(n_1357)
);

OAI22x1_ASAP7_75t_L g1358 ( 
.A1(n_1210),
.A2(n_739),
.B1(n_1033),
.B2(n_724),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1151),
.A2(n_913),
.B(n_926),
.C(n_755),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1144),
.B(n_743),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1115),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1099),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1096),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1123),
.A2(n_1170),
.B1(n_743),
.B2(n_913),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1191),
.B(n_926),
.C(n_913),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1144),
.B(n_1096),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1104),
.A2(n_926),
.B(n_913),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1123),
.B(n_592),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1099),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1151),
.A2(n_913),
.B(n_926),
.C(n_755),
.Y(n_1373)
);

O2A1O1Ixp5_ASAP7_75t_SL g1374 ( 
.A1(n_1135),
.A2(n_1119),
.B(n_1246),
.C(n_489),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_SL g1375 ( 
.A(n_1117),
.B(n_926),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1123),
.B(n_592),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1099),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1115),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1216),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1212),
.A2(n_1068),
.B(n_916),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1158),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1244),
.A2(n_1249),
.A3(n_1246),
.B(n_1243),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1104),
.A2(n_926),
.B(n_913),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1099),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1096),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1390)
);

OAI22x1_ASAP7_75t_L g1391 ( 
.A1(n_1210),
.A2(n_739),
.B1(n_1033),
.B2(n_724),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1123),
.B(n_592),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1144),
.B(n_604),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1105),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1244),
.A2(n_1249),
.A3(n_1246),
.B(n_1243),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1151),
.A2(n_913),
.B(n_926),
.C(n_755),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1149),
.B(n_922),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1105),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1152),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1244),
.A2(n_1249),
.A3(n_1246),
.B(n_1243),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1242),
.A2(n_1243),
.B(n_1220),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1151),
.A2(n_913),
.B(n_926),
.C(n_755),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1243),
.A2(n_1242),
.B(n_1249),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1108),
.A2(n_1001),
.B(n_997),
.Y(n_1405)
);

OAI21xp33_ASAP7_75t_L g1406 ( 
.A1(n_1104),
.A2(n_743),
.B(n_755),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1099),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1144),
.B(n_743),
.Y(n_1408)
);

OAI22x1_ASAP7_75t_L g1409 ( 
.A1(n_1210),
.A2(n_739),
.B1(n_1033),
.B2(n_724),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1108),
.A2(n_1001),
.B(n_997),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1108),
.A2(n_1001),
.B(n_997),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1123),
.B(n_676),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1104),
.B(n_926),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1365),
.A2(n_1406),
.B(n_1279),
.C(n_1359),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1365),
.A2(n_1391),
.B1(n_1409),
.B2(n_1358),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1350),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1316),
.A2(n_1289),
.B(n_1292),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1367),
.B(n_1275),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1325),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1308),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1382),
.A2(n_1349),
.B(n_1406),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1309),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1289),
.A2(n_1251),
.B(n_1268),
.Y(n_1425)
);

CKINVDCx6p67_ASAP7_75t_R g1426 ( 
.A(n_1257),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1370),
.A2(n_1376),
.B(n_1371),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1380),
.A2(n_1389),
.B(n_1386),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1397),
.B(n_1364),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1364),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1270),
.A2(n_1373),
.B(n_1351),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1412),
.A2(n_1392),
.B1(n_1377),
.B2(n_1369),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1279),
.A2(n_1396),
.B1(n_1403),
.B2(n_1321),
.C(n_1368),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1412),
.A2(n_1325),
.B1(n_1265),
.B2(n_1408),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1301),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1385),
.A2(n_1254),
.B(n_1262),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1390),
.A2(n_1402),
.B(n_1399),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_SL g1438 ( 
.A(n_1366),
.B(n_1385),
.C(n_1326),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1366),
.A2(n_1314),
.B(n_1265),
.C(n_1261),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1280),
.A2(n_1276),
.B(n_1286),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1290),
.A2(n_1413),
.B(n_1357),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1258),
.A2(n_1259),
.B(n_1410),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1268),
.A2(n_1266),
.B(n_1290),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1356),
.A2(n_1411),
.B(n_1405),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1256),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1311),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1311),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1253),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1283),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1318),
.B(n_1295),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1274),
.A2(n_1320),
.B(n_1374),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1304),
.B(n_1397),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1304),
.B(n_1336),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1296),
.A2(n_1404),
.B(n_1375),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1281),
.B(n_1322),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1327),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1266),
.A2(n_1404),
.B(n_1305),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1260),
.A2(n_1269),
.B(n_1314),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1323),
.A2(n_1335),
.B(n_1342),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1339),
.A2(n_1334),
.B(n_1260),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1299),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1302),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1310),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1277),
.A2(n_1272),
.B1(n_1312),
.B2(n_1319),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1269),
.A2(n_1330),
.B(n_1300),
.Y(n_1465)
);

OR3x4_ASAP7_75t_SL g1466 ( 
.A(n_1348),
.B(n_1400),
.C(n_1340),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1255),
.A2(n_1303),
.B(n_1328),
.C(n_1333),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1252),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1315),
.A2(n_1393),
.B1(n_1379),
.B2(n_1362),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1345),
.A2(n_1344),
.B(n_1355),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1282),
.A2(n_1388),
.B1(n_1307),
.B2(n_1263),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1317),
.A2(n_1363),
.B(n_1353),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1264),
.A2(n_1388),
.B(n_1287),
.Y(n_1473)
);

A2O1A1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1298),
.A2(n_1332),
.B(n_1387),
.C(n_1378),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1346),
.A2(n_1407),
.B1(n_1372),
.B2(n_1288),
.C(n_1383),
.Y(n_1475)
);

NAND2x1_ASAP7_75t_L g1476 ( 
.A(n_1313),
.B(n_1336),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1293),
.A2(n_1284),
.A3(n_1297),
.B(n_1267),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1253),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1343),
.A2(n_1294),
.B(n_1273),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1284),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1284),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1291),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1313),
.A2(n_1341),
.B(n_1395),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1394),
.Y(n_1484)
);

AOI21xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1271),
.A2(n_1324),
.B(n_1337),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1331),
.A2(n_1297),
.B(n_1338),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1278),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1285),
.A2(n_1398),
.B1(n_1381),
.B2(n_1306),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1293),
.A2(n_1384),
.B(n_1395),
.C(n_1401),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1384),
.A2(n_1401),
.B(n_1306),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1278),
.Y(n_1491)
);

NAND2xp33_ASAP7_75t_SL g1492 ( 
.A(n_1329),
.B(n_1381),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1329),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1329),
.A2(n_1123),
.B1(n_1365),
.B2(n_1358),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1384),
.Y(n_1495)
);

BUFx2_ASAP7_75t_R g1496 ( 
.A(n_1350),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1289),
.A2(n_1251),
.B(n_1268),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1382),
.A2(n_1349),
.B(n_1406),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1325),
.B(n_1304),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1325),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_1350),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1365),
.A2(n_755),
.B(n_743),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1325),
.B(n_1304),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1365),
.A2(n_1123),
.B1(n_1377),
.B2(n_1369),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1253),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_926),
.B1(n_1359),
.B2(n_1351),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1308),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1289),
.A2(n_1251),
.B(n_1268),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1325),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1512)
);

CKINVDCx6p67_ASAP7_75t_R g1513 ( 
.A(n_1257),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1308),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1308),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1365),
.A2(n_1123),
.B1(n_1391),
.B2(n_1358),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1301),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1253),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1365),
.B(n_1123),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1301),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1365),
.A2(n_926),
.B1(n_1359),
.B2(n_1351),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1365),
.A2(n_926),
.B1(n_1359),
.B2(n_1351),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1367),
.B(n_1275),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1365),
.A2(n_1406),
.B(n_913),
.C(n_1279),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1301),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1325),
.B(n_1368),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1347),
.B(n_1360),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1289),
.A2(n_1251),
.B(n_1268),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1382),
.A2(n_1349),
.B(n_1406),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1253),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1393),
.B(n_1144),
.Y(n_1539)
);

AO31x2_ASAP7_75t_L g1540 ( 
.A1(n_1251),
.A2(n_1244),
.A3(n_1246),
.B(n_1249),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1365),
.A2(n_1123),
.B1(n_1391),
.B2(n_1358),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1308),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1382),
.A2(n_1349),
.B(n_1406),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1364),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1308),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1308),
.Y(n_1552)
);

BUFx2_ASAP7_75t_R g1553 ( 
.A(n_1350),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1365),
.A2(n_755),
.B(n_743),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1365),
.B(n_1123),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1301),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1352),
.A2(n_1361),
.B(n_1354),
.Y(n_1560)
);

AO31x2_ASAP7_75t_L g1561 ( 
.A1(n_1251),
.A2(n_1244),
.A3(n_1246),
.B(n_1249),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1365),
.B(n_1359),
.C(n_1351),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1365),
.A2(n_926),
.B1(n_1359),
.B2(n_1351),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1347),
.B(n_1360),
.Y(n_1564)
);

CKINVDCx16_ASAP7_75t_R g1565 ( 
.A(n_1257),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1364),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1504),
.A2(n_1557),
.B1(n_1562),
.B2(n_1524),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1508),
.A2(n_1528),
.B(n_1563),
.C(n_1527),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1509),
.B(n_1514),
.Y(n_1571)
);

BUFx12f_ASAP7_75t_L g1572 ( 
.A(n_1417),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1421),
.B(n_1517),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1516),
.B(n_1542),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1529),
.B(n_1482),
.Y(n_1575)
);

O2A1O1Ixp5_ASAP7_75t_L g1576 ( 
.A1(n_1530),
.A2(n_1414),
.B(n_1439),
.C(n_1423),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1548),
.B(n_1552),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1450),
.B(n_1533),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1530),
.A2(n_1439),
.B(n_1414),
.C(n_1418),
.Y(n_1579)
);

AOI21x1_ASAP7_75t_SL g1580 ( 
.A1(n_1564),
.A2(n_1547),
.B(n_1430),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1445),
.Y(n_1581)
);

O2A1O1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1524),
.A2(n_1558),
.B(n_1438),
.C(n_1433),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1450),
.B(n_1566),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1415),
.A2(n_1428),
.B(n_1427),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1558),
.A2(n_1544),
.B(n_1498),
.C(n_1536),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1506),
.A2(n_1432),
.B1(n_1519),
.B2(n_1541),
.Y(n_1587)
);

AND2x2_ASAP7_75t_SL g1588 ( 
.A(n_1416),
.B(n_1494),
.Y(n_1588)
);

AOI221x1_ASAP7_75t_SL g1589 ( 
.A1(n_1471),
.A2(n_1464),
.B1(n_1434),
.B2(n_1449),
.C(n_1461),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1462),
.B(n_1517),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1518),
.B(n_1522),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1435),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1518),
.B(n_1522),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1475),
.B(n_1441),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1436),
.A2(n_1431),
.B(n_1454),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1455),
.B(n_1429),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1525),
.B(n_1532),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1525),
.B(n_1532),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1467),
.A2(n_1474),
.B1(n_1489),
.B2(n_1473),
.C(n_1455),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1467),
.A2(n_1474),
.B1(n_1488),
.B2(n_1469),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1415),
.A2(n_1545),
.B(n_1551),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1425),
.A2(n_1510),
.B(n_1497),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1429),
.B(n_1487),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1420),
.A2(n_1511),
.B1(n_1502),
.B2(n_1521),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1443),
.B(n_1477),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1443),
.B(n_1477),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1491),
.B(n_1485),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1453),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1426),
.A2(n_1513),
.B1(n_1565),
.B2(n_1538),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1426),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1490),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1495),
.A2(n_1481),
.B1(n_1480),
.B2(n_1510),
.C(n_1425),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_SL g1613 ( 
.A1(n_1535),
.A2(n_1466),
.B(n_1444),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_SL g1614 ( 
.A(n_1458),
.B(n_1466),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1513),
.A2(n_1478),
.B1(n_1448),
.B2(n_1538),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1437),
.A2(n_1500),
.B(n_1556),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1535),
.A2(n_1448),
.B(n_1478),
.C(n_1507),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1493),
.B(n_1458),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1507),
.B(n_1486),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1463),
.Y(n_1620)
);

AND2x2_ASAP7_75t_SL g1621 ( 
.A(n_1520),
.B(n_1559),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1486),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1463),
.A2(n_1484),
.B1(n_1496),
.B2(n_1553),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1468),
.B(n_1452),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1452),
.B(n_1470),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1470),
.B(n_1490),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1479),
.B(n_1476),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1456),
.A2(n_1520),
.B(n_1526),
.C(n_1531),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1503),
.B(n_1483),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1456),
.A2(n_1523),
.B1(n_1515),
.B2(n_1534),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1632)
);

AOI211xp5_ASAP7_75t_L g1633 ( 
.A1(n_1457),
.A2(n_1465),
.B(n_1492),
.C(n_1451),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1465),
.B(n_1561),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1492),
.A2(n_1561),
.B1(n_1540),
.B2(n_1526),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1460),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_R g1637 ( 
.A(n_1531),
.B(n_1559),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1540),
.B(n_1561),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1451),
.A2(n_1459),
.B(n_1440),
.C(n_1442),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1540),
.B(n_1534),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1540),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1501),
.A2(n_1537),
.B(n_1555),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1512),
.A2(n_1543),
.B(n_1554),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1446),
.A2(n_1447),
.B(n_1440),
.C(n_1442),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1546),
.B(n_1560),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1549),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1550),
.B(n_1419),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1524),
.A2(n_1365),
.B(n_1558),
.C(n_1557),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1504),
.A2(n_1365),
.B1(n_1557),
.B2(n_1562),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1472),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1473),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1654)
);

NOR2xp67_ASAP7_75t_L g1655 ( 
.A(n_1438),
.B(n_1484),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1524),
.A2(n_934),
.B1(n_1558),
.B2(n_1506),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1484),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1504),
.A2(n_1365),
.B1(n_1557),
.B2(n_1562),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1436),
.A2(n_1498),
.B(n_1423),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1417),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1592),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1590),
.B(n_1647),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1581),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1651),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1618),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1652),
.B(n_1648),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1645),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1652),
.Y(n_1673)
);

AO21x2_ASAP7_75t_L g1674 ( 
.A1(n_1595),
.A2(n_1602),
.B(n_1662),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1638),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1648),
.B(n_1568),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1634),
.B(n_1641),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1617),
.B(n_1629),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1583),
.B(n_1575),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1569),
.B(n_1650),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1614),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1628),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1605),
.B(n_1606),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1622),
.A2(n_1644),
.B(n_1631),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1573),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1620),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1619),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1625),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1593),
.B(n_1597),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1636),
.B(n_1646),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1567),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1571),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1582),
.A2(n_1570),
.B(n_1576),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1591),
.B(n_1598),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1611),
.B(n_1639),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1584),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1617),
.B(n_1629),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1656),
.A2(n_1588),
.B1(n_1600),
.B2(n_1587),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1585),
.B(n_1570),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1584),
.B(n_1601),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1574),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1616),
.B(n_1643),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1577),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1582),
.B(n_1594),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1599),
.A2(n_1607),
.B(n_1653),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1658),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1616),
.B(n_1642),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1699),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1695),
.A2(n_1579),
.B(n_1649),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1708),
.A2(n_1579),
.B1(n_1589),
.B2(n_1660),
.C(n_1659),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1683),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1672),
.B(n_1691),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1673),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1673),
.B(n_1661),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1633),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1691),
.B(n_1642),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1668),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1691),
.B(n_1637),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1665),
.B(n_1596),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1687),
.B(n_1621),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1676),
.B(n_1615),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1665),
.B(n_1603),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1681),
.B(n_1655),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1680),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1704),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1664),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1704),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1683),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1679),
.B(n_1604),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1676),
.A2(n_1588),
.B1(n_1623),
.B2(n_1608),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1671),
.B(n_1624),
.Y(n_1736)
);

AO21x2_ASAP7_75t_L g1737 ( 
.A1(n_1674),
.A2(n_1613),
.B(n_1580),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1713),
.A2(n_1702),
.B1(n_1701),
.B2(n_1695),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1688),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1713),
.A2(n_1708),
.B1(n_1702),
.B2(n_1703),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1723),
.B(n_1679),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1715),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1719),
.A2(n_1698),
.B1(n_1690),
.B2(n_1666),
.C(n_1609),
.Y(n_1745)
);

OAI332xp33_ASAP7_75t_L g1746 ( 
.A1(n_1725),
.A2(n_1705),
.A3(n_1694),
.B1(n_1693),
.B2(n_1707),
.B3(n_1710),
.C1(n_1690),
.C2(n_1667),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1727),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_R g1748 ( 
.A(n_1727),
.B(n_1610),
.Y(n_1748)
);

AOI33xp33_ASAP7_75t_L g1749 ( 
.A1(n_1714),
.A2(n_1698),
.A3(n_1667),
.B1(n_1697),
.B2(n_1684),
.B3(n_1693),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1735),
.A2(n_1703),
.B1(n_1709),
.B2(n_1675),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1722),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1721),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1714),
.A2(n_1697),
.B1(n_1705),
.B2(n_1710),
.C(n_1694),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1735),
.A2(n_1697),
.B1(n_1709),
.B2(n_1703),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1736),
.A2(n_1709),
.B1(n_1703),
.B2(n_1678),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1736),
.A2(n_1709),
.B1(n_1678),
.B2(n_1700),
.C(n_1707),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1717),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1734),
.A2(n_1703),
.B1(n_1675),
.B2(n_1678),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1712),
.A2(n_1698),
.B1(n_1669),
.B2(n_1689),
.C(n_1677),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1737),
.A2(n_1686),
.B(n_1711),
.Y(n_1762)
);

OAI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1734),
.A2(n_1700),
.B1(n_1678),
.B2(n_1696),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1734),
.A2(n_1700),
.B1(n_1678),
.B2(n_1677),
.Y(n_1764)
);

OAI31xp33_ASAP7_75t_L g1765 ( 
.A1(n_1715),
.A2(n_1669),
.A3(n_1685),
.B(n_1689),
.Y(n_1765)
);

NOR2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1717),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1718),
.Y(n_1769)
);

AND2x2_ASAP7_75t_SL g1770 ( 
.A(n_1733),
.B(n_1586),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1723),
.B(n_1726),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1682),
.Y(n_1773)
);

CKINVDCx16_ASAP7_75t_R g1774 ( 
.A(n_1724),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1730),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1731),
.Y(n_1776)
);

NAND4xp25_ASAP7_75t_L g1777 ( 
.A(n_1720),
.B(n_1692),
.C(n_1711),
.D(n_1706),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1737),
.A2(n_1700),
.B1(n_1677),
.B2(n_1675),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1720),
.B(n_1682),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1762),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1752),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1745),
.A2(n_1732),
.B(n_1729),
.Y(n_1782)
);

NOR2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1747),
.B(n_1688),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1762),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1744),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1738),
.B(n_1730),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1767),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1770),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1770),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1772),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1766),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1775),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1744),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1768),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1776),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1771),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1756),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.B(n_1729),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1756),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1747),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1739),
.B(n_1572),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1743),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1779),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1743),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1784),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1800),
.B(n_1740),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1788),
.B(n_1774),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1788),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_L g1809 ( 
.A(n_1782),
.B(n_1753),
.C(n_1749),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1773),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1794),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1800),
.B(n_1746),
.Y(n_1812)
);

INVx4_ASAP7_75t_L g1813 ( 
.A(n_1793),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1788),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1782),
.B(n_1742),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1794),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1802),
.B(n_1760),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1802),
.B(n_1769),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1786),
.B(n_1726),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_1804),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1804),
.B(n_1769),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1794),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1784),
.A2(n_1750),
.B1(n_1757),
.B2(n_1754),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1782),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1784),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1783),
.Y(n_1827)
);

BUFx6f_ASAP7_75t_L g1828 ( 
.A(n_1784),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1780),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1782),
.B(n_1761),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1781),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1789),
.B(n_1751),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1804),
.B(n_1765),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1796),
.B(n_1758),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1780),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1793),
.B(n_1751),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1795),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1782),
.B(n_1803),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1780),
.Y(n_1839)
);

INVx1_ASAP7_75t_SL g1840 ( 
.A(n_1785),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1780),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1807),
.B(n_1791),
.Y(n_1842)
);

A2O1A1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1812),
.A2(n_1801),
.B(n_1778),
.C(n_1755),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1817),
.B(n_1797),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1787),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1840),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1828),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1809),
.B(n_1787),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1809),
.B(n_1797),
.Y(n_1849)
);

NOR2xp67_ASAP7_75t_SL g1850 ( 
.A(n_1827),
.B(n_1657),
.Y(n_1850)
);

OAI21xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1815),
.A2(n_1783),
.B(n_1798),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1824),
.A2(n_1801),
.B(n_1741),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1797),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1818),
.B(n_1799),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1823),
.A2(n_1763),
.B1(n_1759),
.B2(n_1764),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1818),
.B(n_1799),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1831),
.Y(n_1857)
);

INVx1_ASAP7_75t_SL g1858 ( 
.A(n_1806),
.Y(n_1858)
);

NAND3xp33_ASAP7_75t_L g1859 ( 
.A(n_1828),
.B(n_1793),
.C(n_1785),
.Y(n_1859)
);

NAND2xp33_ASAP7_75t_R g1860 ( 
.A(n_1814),
.B(n_1748),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1821),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1821),
.B(n_1799),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1833),
.B(n_1790),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1833),
.B(n_1834),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1807),
.B(n_1791),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1834),
.B(n_1790),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1831),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1828),
.Y(n_1869)
);

AND2x4_ASAP7_75t_SL g1870 ( 
.A(n_1836),
.B(n_1791),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1820),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1828),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1811),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1819),
.B(n_1792),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1828),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1828),
.B(n_1793),
.C(n_1785),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1813),
.B(n_1803),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1811),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1864),
.B(n_1819),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1838),
.Y(n_1880)
);

NOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1859),
.B(n_1813),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1848),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1878),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1878),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1867),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1849),
.B(n_1820),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1867),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1870),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1877),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1846),
.B(n_1838),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1842),
.B(n_1827),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1873),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1870),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1851),
.A2(n_1826),
.B1(n_1824),
.B2(n_1863),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_SL g1897 ( 
.A1(n_1844),
.A2(n_1824),
.B1(n_1826),
.B2(n_1828),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1842),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_L g1899 ( 
.A(n_1876),
.B(n_1813),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1865),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1853),
.B(n_1874),
.Y(n_1901)
);

INVx1_ASAP7_75t_SL g1902 ( 
.A(n_1865),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1857),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1853),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1845),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1882),
.A2(n_1843),
.B1(n_1852),
.B2(n_1826),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1905),
.B(n_1871),
.Y(n_1908)
);

OAI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1895),
.A2(n_1843),
.B(n_1868),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1900),
.B(n_1850),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1881),
.A2(n_1826),
.B(n_1824),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1883),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1882),
.A2(n_1860),
.B1(n_1855),
.B2(n_1850),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1880),
.A2(n_1866),
.B(n_1825),
.Y(n_1914)
);

INVxp33_ASAP7_75t_L g1915 ( 
.A(n_1891),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1884),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1898),
.B(n_1854),
.Y(n_1917)
);

CKINVDCx14_ASAP7_75t_R g1918 ( 
.A(n_1891),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1900),
.B(n_1877),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1902),
.B(n_1856),
.Y(n_1920)
);

O2A1O1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1906),
.A2(n_1886),
.B(n_1901),
.C(n_1887),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1894),
.B(n_1862),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1897),
.B(n_1813),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1896),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1896),
.B(n_1815),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1894),
.B(n_1836),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1885),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1904),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1928),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1918),
.B(n_1888),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1928),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1924),
.Y(n_1932)
);

OAI222xp33_ASAP7_75t_L g1933 ( 
.A1(n_1907),
.A2(n_1886),
.B1(n_1890),
.B2(n_1893),
.C1(n_1879),
.C2(n_1899),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1908),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1917),
.B(n_1889),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1919),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1921),
.B(n_1904),
.Y(n_1937)
);

INVxp67_ASAP7_75t_SL g1938 ( 
.A(n_1909),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1919),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1912),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1918),
.B(n_1904),
.Y(n_1941)
);

AOI21xp33_ASAP7_75t_L g1942 ( 
.A1(n_1938),
.A2(n_1915),
.B(n_1911),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1933),
.A2(n_1914),
.B1(n_1913),
.B2(n_1915),
.C(n_1925),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_SL g1944 ( 
.A1(n_1938),
.A2(n_1920),
.B1(n_1910),
.B2(n_1889),
.C(n_1927),
.Y(n_1944)
);

NAND3x1_ASAP7_75t_L g1945 ( 
.A(n_1937),
.B(n_1941),
.C(n_1930),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1936),
.B(n_1922),
.Y(n_1946)
);

OAI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1933),
.A2(n_1923),
.B(n_1926),
.Y(n_1947)
);

NOR2xp67_ASAP7_75t_L g1948 ( 
.A(n_1939),
.B(n_1923),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1929),
.Y(n_1949)
);

OAI21xp33_ASAP7_75t_L g1950 ( 
.A1(n_1934),
.A2(n_1903),
.B(n_1916),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1935),
.B(n_1836),
.Y(n_1951)
);

AOI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1932),
.A2(n_1892),
.B(n_1875),
.C(n_1872),
.Y(n_1952)
);

OR3x1_ASAP7_75t_L g1953 ( 
.A(n_1931),
.B(n_1822),
.C(n_1816),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1945),
.B(n_1940),
.Y(n_1954)
);

OAI21xp33_ASAP7_75t_L g1955 ( 
.A1(n_1947),
.A2(n_1869),
.B(n_1847),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1942),
.B(n_1869),
.C(n_1847),
.Y(n_1956)
);

AOI22x1_ASAP7_75t_L g1957 ( 
.A1(n_1949),
.A2(n_1875),
.B1(n_1872),
.B2(n_1814),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1953),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1946),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1948),
.B(n_1836),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1960),
.B(n_1943),
.Y(n_1961)
);

AOI221x1_ASAP7_75t_L g1962 ( 
.A1(n_1959),
.A2(n_1950),
.B1(n_1944),
.B2(n_1805),
.C(n_1825),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1954),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1958),
.B(n_1951),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1954),
.B(n_1952),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1956),
.Y(n_1966)
);

NAND3xp33_ASAP7_75t_L g1967 ( 
.A(n_1957),
.B(n_1825),
.C(n_1805),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1961),
.A2(n_1955),
.B1(n_1805),
.B2(n_1815),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1963),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1966),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_R g1971 ( 
.A(n_1965),
.B(n_1663),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_R g1972 ( 
.A(n_1964),
.B(n_1627),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1961),
.B(n_1832),
.Y(n_1973)
);

AOI21xp33_ASAP7_75t_SL g1974 ( 
.A1(n_1973),
.A2(n_1967),
.B(n_1962),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1969),
.B(n_1832),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1970),
.B(n_1832),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_1976),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1977),
.Y(n_1978)
);

XOR2xp5_ASAP7_75t_L g1979 ( 
.A(n_1978),
.B(n_1968),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1978),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1980),
.Y(n_1981)
);

OAI22x1_ASAP7_75t_L g1982 ( 
.A1(n_1979),
.A2(n_1971),
.B1(n_1974),
.B2(n_1972),
.Y(n_1982)
);

NAND4xp75_ASAP7_75t_L g1983 ( 
.A(n_1981),
.B(n_1830),
.C(n_1829),
.D(n_1839),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1982),
.Y(n_1984)
);

AO22x2_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1835),
.B1(n_1808),
.B2(n_1839),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1983),
.B(n_1835),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1986),
.B(n_1829),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1808),
.B1(n_1829),
.B2(n_1841),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1808),
.B1(n_1816),
.B2(n_1837),
.Y(n_1989)
);

AOI211xp5_ASAP7_75t_L g1990 ( 
.A1(n_1989),
.A2(n_1839),
.B(n_1841),
.C(n_1808),
.Y(n_1990)
);


endmodule