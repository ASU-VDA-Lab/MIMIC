module real_jpeg_33700_n_32 (n_17, n_232, n_8, n_0, n_21, n_2, n_229, n_226, n_29, n_10, n_31, n_9, n_12, n_24, n_6, n_221, n_223, n_28, n_230, n_231, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_224, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_222, n_228, n_30, n_227, n_220, n_16, n_15, n_13, n_225, n_32);

input n_17;
input n_232;
input n_8;
input n_0;
input n_21;
input n_2;
input n_229;
input n_226;
input n_29;
input n_10;
input n_31;
input n_9;
input n_12;
input n_24;
input n_6;
input n_221;
input n_223;
input n_28;
input n_230;
input n_231;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_224;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_222;
input n_228;
input n_30;
input n_227;
input n_220;
input n_16;
input n_15;
input n_13;
input n_225;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_203;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_80;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_138;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_67),
.C(n_205),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_2),
.B(n_134),
.Y(n_133)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_2),
.B(n_180),
.CON(n_179),
.SN(n_179)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_119),
.A3(n_121),
.B1(n_126),
.B2(n_183),
.C1(n_185),
.C2(n_230),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_6),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_6),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_7),
.Y(n_99)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_105),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_11),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_13),
.B(n_98),
.Y(n_203)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_14),
.A2(n_16),
.B1(n_148),
.B2(n_152),
.C(n_154),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_148),
.C(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_15),
.A2(n_69),
.B1(n_189),
.B2(n_204),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_17),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_18),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_19),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_19),
.A2(n_211),
.B(n_216),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_19),
.B(n_211),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_21),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_21),
.B(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_23),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_24),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_28),
.B(n_128),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_31),
.B(n_92),
.Y(n_200)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_47),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_44),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_50),
.B(n_52),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_46),
.B(n_50),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_63),
.B(n_210),
.C(n_217),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_62),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_110),
.B(n_188),
.Y(n_67)
);

NAND4xp25_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.C(n_96),
.D(n_103),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_70),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_80),
.C(n_84),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_75),
.B(n_198),
.C(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_76),
.B(n_79),
.Y(n_192)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

OAI322xp33_ASAP7_75t_L g196 ( 
.A1(n_80),
.A2(n_86),
.A3(n_197),
.B1(n_200),
.B2(n_201),
.C1(n_202),
.C2(n_232),
.Y(n_196)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g190 ( 
.A1(n_85),
.A2(n_191),
.A3(n_192),
.B1(n_193),
.B2(n_196),
.C(n_231),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_91),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_97),
.A2(n_190),
.B(n_203),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI31xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_138),
.A3(n_170),
.B(n_177),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_125),
.C(n_133),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_112),
.A2(n_178),
.B(n_182),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_133),
.C(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_221),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OA21x2_ASAP7_75t_SL g178 ( 
.A1(n_125),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_165),
.C(n_166),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_158),
.B(n_164),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_226),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_163),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_179),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_220),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_222),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_223),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_224),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_225),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_227),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_228),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_229),
.Y(n_173)
);


endmodule