module fake_jpeg_16281_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_40),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_31),
.B1(n_21),
.B2(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_47),
.B1(n_34),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_15),
.B1(n_30),
.B2(n_23),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_31),
.B1(n_21),
.B2(n_20),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_31),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_34),
.B(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_31),
.B1(n_21),
.B2(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_18),
.B1(n_35),
.B2(n_38),
.Y(n_75)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_40),
.B1(n_36),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_64),
.B1(n_78),
.B2(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_72),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_64)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_34),
.A3(n_25),
.B1(n_30),
.B2(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_18),
.B1(n_35),
.B2(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_79),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_19),
.CON(n_77),
.SN(n_77)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_37),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_37),
.B1(n_27),
.B2(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_17),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_27),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_37),
.B1(n_54),
.B2(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_63),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_52),
.B1(n_46),
.B2(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_89),
.B1(n_96),
.B2(n_80),
.Y(n_128)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_71),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_46),
.B1(n_56),
.B2(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_61),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_67),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_109),
.B(n_81),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_65),
.A2(n_46),
.B1(n_56),
.B2(n_49),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_68),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_37),
.B1(n_56),
.B2(n_27),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_82),
.B1(n_60),
.B2(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_83),
.C(n_79),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_127),
.C(n_119),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_119),
.B1(n_137),
.B2(n_103),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_118),
.B(n_135),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_93),
.B1(n_102),
.B2(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_16),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_98),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_64),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_67),
.B1(n_73),
.B2(n_43),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_138),
.B1(n_87),
.B2(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_100),
.B(n_88),
.C(n_101),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_43),
.B1(n_16),
.B2(n_27),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_22),
.B1(n_14),
.B2(n_11),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_33),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_144),
.C(n_151),
.Y(n_178)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_147),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_146),
.B1(n_153),
.B2(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_92),
.B1(n_99),
.B2(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_170),
.B1(n_132),
.B2(n_131),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_160),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_84),
.A3(n_131),
.B1(n_24),
.B2(n_19),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_33),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_92),
.B1(n_106),
.B2(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_117),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_161),
.C(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_24),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_33),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_125),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_22),
.B(n_28),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_22),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_115),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_123),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_114),
.A2(n_55),
.B1(n_19),
.B2(n_17),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_55),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_185),
.C(n_194),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_19),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_187),
.B(n_199),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_55),
.C(n_84),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_164),
.B(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_198),
.B1(n_200),
.B2(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_197),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_28),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_28),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_196),
.C(n_170),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_22),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_164),
.B(n_159),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_184),
.B(n_199),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_216),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_153),
.B1(n_163),
.B2(n_141),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_211),
.B1(n_224),
.B2(n_225),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_202),
.A2(n_140),
.B1(n_166),
.B2(n_165),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_19),
.C(n_24),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_217),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_14),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_1),
.C(n_2),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_172),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_228),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_186),
.B1(n_192),
.B2(n_176),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_212),
.B1(n_221),
.B2(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_238),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_236),
.A2(n_237),
.B(n_239),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_190),
.B(n_180),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_190),
.B(n_200),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_186),
.B(n_173),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_243),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_205),
.B1(n_181),
.B2(n_188),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_209),
.B(n_178),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_185),
.C(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_254),
.C(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_214),
.C(n_213),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_219),
.B1(n_207),
.B2(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_194),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_217),
.C(n_211),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_210),
.B1(n_224),
.B2(n_195),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_236),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_196),
.C(n_6),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_239),
.C(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_275),
.C(n_278),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_276),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_11),
.B(n_13),
.Y(n_293)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_237),
.B(n_230),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_231),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_262),
.B1(n_257),
.B2(n_249),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_250),
.C(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_290),
.C(n_292),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_265),
.B1(n_238),
.B2(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_267),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_253),
.CI(n_238),
.CON(n_288),
.SN(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_10),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_253),
.C(n_6),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_5),
.C(n_7),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_7),
.C(n_8),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_277),
.B1(n_269),
.B2(n_274),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_12),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_13),
.B1(n_14),
.B2(n_9),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.C(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_282),
.CI(n_283),
.CON(n_307),
.SN(n_307)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_303),
.C(n_296),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_295),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.C(n_307),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_305),
.B(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_306),
.B(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_281),
.Y(n_318)
);

OAI321xp33_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_281),
.A3(n_290),
.B1(n_304),
.B2(n_288),
.C(n_9),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_9),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_9),
.B(n_304),
.Y(n_321)
);


endmodule