module fake_jpeg_8558_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_5),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_21),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_7),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_24),
.C(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_2),
.Y(n_21)
);

OR2x2_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_3),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_11),
.B(n_9),
.C(n_16),
.D(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVxp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_19),
.B(n_4),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_30),
.B1(n_29),
.B2(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_14),
.B1(n_9),
.B2(n_5),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_14),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_42)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_29),
.B1(n_27),
.B2(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_32),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_42),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_47),
.B1(n_40),
.B2(n_41),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_50),
.B(n_48),
.C(n_44),
.Y(n_52)
);

OAI21x1_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_43),
.B(n_46),
.Y(n_53)
);


endmodule