module real_jpeg_31255_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_0),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_0),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_0),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_2),
.B(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_2),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_5),
.B(n_101),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_5),
.B(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_6),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_7),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_7),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_8),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_8),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_8),
.B(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_10),
.B(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_13),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_13),
.Y(n_225)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_14),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_14),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_14),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_15),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_15),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_193),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_143),
.B(n_192),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_96),
.B(n_142),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_L g142 ( 
.A(n_21),
.B(n_63),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.C(n_53),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_23),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_36),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_36),
.C(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_27),
.B(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_35),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_38),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_44),
.A2(n_53),
.B1(n_54),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_47),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_48),
.Y(n_153)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_57),
.Y(n_186)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_81),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_79),
.B2(n_80),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_R g146 ( 
.A(n_67),
.B(n_71),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_67),
.B(n_190),
.C(n_191),
.Y(n_189)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2x1_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_72),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_145),
.C(n_146),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_84),
.C(n_91),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

AOI21x1_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_113),
.B(n_141),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_109),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.C(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_102),
.Y(n_236)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_134),
.B(n_140),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_129),
.B(n_133),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_120),
.Y(n_133)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_126),
.Y(n_135)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_147),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_169),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_168),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_168),
.C(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_167),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_160),
.C(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_152),
.B(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_160),
.B1(n_161),
.B2(n_166),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_183),
.C(n_189),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_178),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_176),
.C(n_179),
.Y(n_217)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_243),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_219),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_213),
.B2(n_218),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_242),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_228),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_226),
.Y(n_228)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_235),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);


endmodule