module fake_netlist_5_1486_n_1089 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1089);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1089;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_1073;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_1020;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_897;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1075;
wire n_1069;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_989;
wire n_1041;
wire n_852;
wire n_1039;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_952;
wire n_809;
wire n_931;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_868;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_1032;
wire n_1056;
wire n_960;
wire n_890;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_45),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_5),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_33),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_17),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_130),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_198),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_84),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_112),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_49),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_94),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_87),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_67),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_77),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_124),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_160),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_71),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_151),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_172),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_153),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_57),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_152),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_61),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_5),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_76),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_69),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_136),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_38),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_95),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_68),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_41),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_51),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_189),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_163),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_23),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_116),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_79),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_103),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_203),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_213),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_236),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_208),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_228),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_246),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_233),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_260),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_218),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_262),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_209),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_223),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_210),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_211),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_302),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

OAI22x1_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_266),
.B1(n_265),
.B2(n_238),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_303),
.A2(n_275),
.B1(n_262),
.B2(n_272),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_215),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_216),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_217),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_222),
.B(n_221),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_224),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_280),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_225),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_227),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_279),
.B(n_275),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_283),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_249),
.B1(n_271),
.B2(n_270),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_231),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_320),
.B(n_232),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_300),
.A2(n_274),
.B1(n_269),
.B2(n_267),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_314),
.A2(n_264),
.B1(n_263),
.B2(n_253),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_234),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

NAND2x1_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_235),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_320),
.B(n_237),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_277),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_281),
.A2(n_287),
.B(n_286),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_276),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_286),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_250),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_281),
.Y(n_379)
);

BUFx8_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_335),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_287),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

OR2x6_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_299),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_313),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_312),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_305),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_363),
.B(n_319),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

AND3x2_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_323),
.C(n_291),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_289),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_349),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_338),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_330),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_330),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_289),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_291),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_348),
.B(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_349),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

NAND3xp33_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_323),
.C(n_296),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_329),
.A2(n_308),
.B1(n_299),
.B2(n_316),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_369),
.B(n_239),
.Y(n_426)
);

INVx8_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_316),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_342),
.B(n_292),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_369),
.B(n_242),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_327),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_364),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_327),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_361),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_317),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_328),
.B(n_317),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_346),
.Y(n_443)
);

AND3x1_ASAP7_75t_L g444 ( 
.A(n_358),
.B(n_296),
.C(n_292),
.Y(n_444)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_371),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_361),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_341),
.B(n_298),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_343),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_328),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_343),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_333),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_404),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_381),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_398),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_414),
.B(n_343),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_381),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_357),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_389),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_404),
.B(n_326),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_336),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_391),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_412),
.B(n_357),
.Y(n_484)
);

XNOR2x2_ASAP7_75t_L g485 ( 
.A(n_405),
.B(n_298),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_371),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_341),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_337),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_383),
.B(n_333),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_399),
.B(n_245),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_397),
.B(n_451),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_424),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_R g499 ( 
.A(n_437),
.B(n_413),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_430),
.B(n_341),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_413),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_442),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_441),
.B(n_376),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_436),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_426),
.B(n_346),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_445),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_440),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_392),
.B(n_362),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_446),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_447),
.Y(n_519)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_442),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_445),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_448),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_428),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_346),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_396),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_463),
.B(n_385),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_455),
.A2(n_451),
.B1(n_416),
.B2(n_437),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_385),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_464),
.B(n_385),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_416),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_495),
.B(n_397),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_502),
.B(n_416),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_525),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_456),
.B(n_416),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_495),
.B(n_416),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_427),
.Y(n_547)
);

NAND2x1_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_406),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_498),
.Y(n_549)
);

NOR3xp33_ASAP7_75t_L g550 ( 
.A(n_458),
.B(n_311),
.C(n_339),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_478),
.B(n_385),
.Y(n_551)
);

AND2x6_ASAP7_75t_SL g552 ( 
.A(n_516),
.B(n_311),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_495),
.B(n_397),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_469),
.B(n_427),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_465),
.A2(n_427),
.B1(n_444),
.B2(n_395),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_455),
.B(n_427),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_503),
.B(n_511),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_466),
.A2(n_395),
.B1(n_425),
.B2(n_403),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_395),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_489),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_530),
.B(n_448),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_522),
.B(n_445),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_476),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_445),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_520),
.A2(n_410),
.B1(n_431),
.B2(n_422),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_527),
.B(n_475),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_454),
.B(n_362),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_520),
.B(n_362),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_380),
.C(n_248),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_475),
.B(n_390),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_497),
.A2(n_521),
.B1(n_504),
.B2(n_471),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_453),
.B(n_390),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_468),
.B(n_376),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

AND2x6_ASAP7_75t_SL g582 ( 
.A(n_516),
.B(n_380),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_472),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_533),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_522),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_533),
.B(n_402),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_488),
.A2(n_411),
.B1(n_431),
.B2(n_422),
.Y(n_588)
);

AND2x6_ASAP7_75t_SL g589 ( 
.A(n_484),
.B(n_380),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_473),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_521),
.B(n_402),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_376),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_493),
.A2(n_410),
.B1(n_406),
.B2(n_418),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_494),
.A2(n_344),
.B(n_347),
.C(n_354),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_474),
.A2(n_375),
.B1(n_409),
.B2(n_418),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_488),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

OAI221xp5_ASAP7_75t_L g598 ( 
.A1(n_526),
.A2(n_376),
.B1(n_353),
.B2(n_379),
.C(n_375),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_496),
.B(n_402),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_528),
.Y(n_600)
);

AND2x4_ASAP7_75t_SL g601 ( 
.A(n_497),
.B(n_448),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_597),
.B(n_494),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_SL g604 ( 
.A(n_591),
.B(n_499),
.C(n_529),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_563),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_SL g606 ( 
.A(n_591),
.B(n_531),
.C(n_532),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_566),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_538),
.B(n_534),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_541),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_536),
.B(n_500),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_536),
.B(n_509),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_596),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_501),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_SL g614 ( 
.A(n_567),
.B(n_506),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_535),
.B(n_601),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_538),
.B(n_507),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_554),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_583),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_571),
.B(n_508),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_539),
.B(n_510),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_581),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_586),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_545),
.B(n_547),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_542),
.B(n_513),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_555),
.B(n_512),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_557),
.A2(n_448),
.B(n_514),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_565),
.B(n_515),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_601),
.B(n_524),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_R g634 ( 
.A(n_537),
.B(n_517),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_558),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_573),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_544),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_579),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_586),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_549),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_549),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_596),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_537),
.A2(n_492),
.B1(n_491),
.B2(n_483),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

NOR2x1_ASAP7_75t_L g645 ( 
.A(n_575),
.B(n_518),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_576),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_580),
.B(n_519),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_556),
.B(n_481),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_580),
.B(n_523),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_R g650 ( 
.A(n_560),
.B(n_477),
.Y(n_650)
);

OR2x2_ASAP7_75t_SL g651 ( 
.A(n_552),
.B(n_375),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_600),
.B(n_479),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_551),
.B(n_480),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_550),
.B(n_407),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_570),
.B(n_421),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_544),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_551),
.B(n_421),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_550),
.B(n_407),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_578),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_612),
.Y(n_662)
);

AOI21xp33_ASAP7_75t_L g663 ( 
.A1(n_634),
.A2(n_572),
.B(n_574),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_657),
.B(n_592),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_657),
.B(n_574),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_630),
.A2(n_564),
.B(n_548),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_613),
.B(n_540),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_646),
.B(n_540),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_607),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_624),
.A2(n_598),
.B(n_564),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_615),
.B(n_553),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_620),
.B(n_553),
.Y(n_672)
);

OAI21x1_ASAP7_75t_SL g673 ( 
.A1(n_655),
.A2(n_561),
.B(n_562),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_611),
.A2(n_546),
.B(n_588),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_606),
.B(n_604),
.C(n_634),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_610),
.A2(n_595),
.B1(n_580),
.B2(n_599),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_624),
.A2(n_595),
.B(n_569),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_594),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_621),
.A2(n_593),
.B(n_411),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_621),
.A2(n_409),
.B(n_421),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_629),
.A2(n_368),
.B(n_366),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_611),
.A2(n_368),
.B(n_366),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_652),
.B(n_582),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_632),
.B(n_366),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_614),
.A2(n_368),
.B(n_366),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_622),
.A2(n_589),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_648),
.A2(n_36),
.B(n_34),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_661),
.B(n_0),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_656),
.B(n_638),
.Y(n_689)
);

AOI21xp33_ASAP7_75t_L g690 ( 
.A1(n_659),
.A2(n_2),
.B(n_3),
.Y(n_690)
);

NAND2x1p5_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_37),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_610),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_648),
.A2(n_645),
.B(n_660),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_623),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_637),
.B(n_39),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_654),
.A2(n_44),
.B(n_40),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_654),
.A2(n_48),
.B(n_47),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_659),
.A2(n_52),
.B(n_50),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_650),
.B(n_4),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_604),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_643),
.A2(n_55),
.B(n_53),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_644),
.Y(n_702)
);

AO31x2_ASAP7_75t_L g703 ( 
.A1(n_609),
.A2(n_8),
.A3(n_9),
.B(n_10),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_625),
.A2(n_58),
.B(n_56),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_618),
.A2(n_60),
.B(n_59),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_607),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_653),
.B(n_9),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_625),
.A2(n_606),
.B(n_603),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_647),
.A2(n_118),
.B(n_204),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_647),
.A2(n_649),
.B(n_616),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_625),
.A2(n_206),
.B(n_117),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_625),
.A2(n_202),
.B(n_115),
.Y(n_713)
);

AO221x2_ASAP7_75t_L g714 ( 
.A1(n_628),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_714)
);

AO31x2_ASAP7_75t_L g715 ( 
.A1(n_640),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_663),
.A2(n_602),
.B(n_605),
.C(n_649),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_694),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_693),
.A2(n_641),
.B(n_619),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_711),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_665),
.B(n_639),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_710),
.B(n_612),
.Y(n_721)
);

INVx3_ASAP7_75t_SL g722 ( 
.A(n_662),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_683),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_699),
.B(n_608),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_698),
.A2(n_647),
.B(n_608),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_666),
.A2(n_680),
.B(n_679),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_688),
.B(n_617),
.Y(n_729)
);

OAI22x1_ASAP7_75t_L g730 ( 
.A1(n_675),
.A2(n_627),
.B1(n_633),
.B2(n_635),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_674),
.A2(n_602),
.B(n_612),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_690),
.A2(n_636),
.B(n_644),
.C(n_658),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_692),
.A2(n_658),
.B(n_651),
.C(n_650),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_L g734 ( 
.A1(n_678),
.A2(n_625),
.B(n_631),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_682),
.A2(n_631),
.B(n_642),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_702),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_689),
.B(n_642),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_706),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_670),
.A2(n_642),
.B(n_121),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_702),
.Y(n_740)
);

AOI221x1_ASAP7_75t_L g741 ( 
.A1(n_700),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_17),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_670),
.A2(n_122),
.B(n_197),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_691),
.B(n_62),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_664),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_667),
.B(n_15),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_715),
.Y(n_746)
);

AOI21x1_ASAP7_75t_L g747 ( 
.A1(n_677),
.A2(n_123),
.B(n_194),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_715),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_708),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_684),
.Y(n_750)
);

AO31x2_ASAP7_75t_L g751 ( 
.A1(n_676),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_707),
.B(n_20),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_671),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_672),
.A2(n_126),
.B(n_192),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_673),
.A2(n_125),
.B(n_191),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_675),
.A2(n_21),
.B(n_22),
.Y(n_756)
);

AO32x2_ASAP7_75t_L g757 ( 
.A1(n_714),
.A2(n_21),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_757)
);

AOI221x1_ASAP7_75t_L g758 ( 
.A1(n_704),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_704),
.A2(n_199),
.B(n_129),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_712),
.A2(n_188),
.B(n_128),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_668),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_712),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_703),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_681),
.A2(n_132),
.B(n_186),
.Y(n_765)
);

AO31x2_ASAP7_75t_L g766 ( 
.A1(n_685),
.A2(n_29),
.A3(n_30),
.B(n_31),
.Y(n_766)
);

AO32x2_ASAP7_75t_L g767 ( 
.A1(n_714),
.A2(n_703),
.A3(n_708),
.B1(n_713),
.B2(n_705),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_701),
.A2(n_131),
.B(n_185),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_713),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_687),
.Y(n_770)
);

INVx3_ASAP7_75t_SL g771 ( 
.A(n_691),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_695),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_686),
.B(n_63),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_695),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_703),
.B(n_709),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_697),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_776)
);

AO31x2_ASAP7_75t_L g777 ( 
.A1(n_696),
.A2(n_32),
.A3(n_65),
.B(n_66),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_753),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_720),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_773),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_758),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_719),
.Y(n_782)
);

CKINVDCx8_ASAP7_75t_R g783 ( 
.A(n_725),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_726),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_SL g785 ( 
.A1(n_756),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_717),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_743),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_764),
.Y(n_789)
);

BUFx4f_ASAP7_75t_SL g790 ( 
.A(n_722),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_752),
.B(n_88),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_746),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_738),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_769),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_723),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_758),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_SL g797 ( 
.A1(n_759),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_748),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_737),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_760),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_736),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_763),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_761),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_744),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_762),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_718),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_724),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_776),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_SL g810 ( 
.A1(n_741),
.A2(n_114),
.B(n_119),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_745),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_771),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_723),
.Y(n_813)
);

BUFx2_ASAP7_75t_SL g814 ( 
.A(n_723),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_751),
.Y(n_815)
);

INVx5_ASAP7_75t_L g816 ( 
.A(n_743),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_734),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_750),
.B(n_140),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_772),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_751),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_716),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_772),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_751),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_742),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_721),
.B(n_155),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_730),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_721),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_727),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_828)
);

INVx8_ASAP7_75t_L g829 ( 
.A(n_774),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_731),
.B(n_159),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_757),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_831)
);

INVx6_ASAP7_75t_L g832 ( 
.A(n_775),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_739),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_792),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_832),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_807),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_782),
.Y(n_837)
);

AO21x1_ASAP7_75t_L g838 ( 
.A1(n_831),
.A2(n_757),
.B(n_755),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_788),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_798),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_800),
.Y(n_841)
);

INVx8_ASAP7_75t_L g842 ( 
.A(n_829),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_827),
.B(n_770),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_789),
.Y(n_844)
);

OAI21xp33_ASAP7_75t_SL g845 ( 
.A1(n_831),
.A2(n_780),
.B(n_811),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_795),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_815),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_826),
.B(n_728),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_804),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_799),
.B(n_766),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_804),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_806),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_820),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_823),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_832),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_785),
.A2(n_733),
.B1(n_754),
.B2(n_732),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_799),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_830),
.A2(n_747),
.B(n_768),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_828),
.A2(n_747),
.B(n_765),
.Y(n_859)
);

OAI211xp5_ASAP7_75t_L g860 ( 
.A1(n_810),
.A2(n_757),
.B(n_767),
.C(n_749),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_828),
.A2(n_735),
.B(n_767),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_813),
.Y(n_864)
);

OA21x2_ASAP7_75t_L g865 ( 
.A1(n_810),
.A2(n_767),
.B(n_766),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_793),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_813),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_783),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_813),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_825),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_784),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_779),
.B(n_766),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_780),
.A2(n_777),
.B(n_169),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_781),
.B(n_796),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_838),
.A2(n_802),
.B(n_821),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_834),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_834),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_840),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_836),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_857),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_840),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_873),
.B(n_784),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_835),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_841),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_857),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_842),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_835),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_861),
.B(n_787),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_841),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_842),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_873),
.B(n_777),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_847),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_861),
.B(n_777),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_851),
.B(n_787),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_844),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_844),
.B(n_787),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_847),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_854),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_837),
.B(n_816),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_894),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_892),
.B(n_865),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_884),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_894),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_892),
.B(n_865),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_894),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_899),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_899),
.B(n_848),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_899),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_900),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_900),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_900),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_880),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_880),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_889),
.B(n_872),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_877),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_884),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_881),
.B(n_850),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_877),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_888),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_883),
.B(n_865),
.Y(n_922)
);

OAI221xp5_ASAP7_75t_SL g923 ( 
.A1(n_875),
.A2(n_845),
.B1(n_860),
.B2(n_794),
.C(n_811),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_875),
.A2(n_856),
.B1(n_816),
.B2(n_797),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_922),
.B(n_888),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_917),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_904),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_917),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_905),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_905),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_905),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_922),
.B(n_883),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_909),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_922),
.B(n_898),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_903),
.B(n_898),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_920),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_903),
.B(n_886),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_912),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_912),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_929),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_927),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_928),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_919),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_927),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_932),
.B(n_919),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_935),
.B(n_903),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_929),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_932),
.B(n_916),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_934),
.B(n_906),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_934),
.B(n_904),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_906),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_R g954 ( 
.A(n_952),
.B(n_947),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_946),
.B(n_938),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_944),
.B(n_950),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_952),
.B(n_925),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_943),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_949),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_942),
.B(n_938),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_945),
.B(n_936),
.Y(n_961)
);

AO221x2_ASAP7_75t_L g962 ( 
.A1(n_954),
.A2(n_961),
.B1(n_959),
.B2(n_958),
.C(n_866),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_956),
.A2(n_923),
.B1(n_924),
.B2(n_952),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_961),
.B(n_945),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_957),
.Y(n_965)
);

NAND2xp33_ASAP7_75t_SL g966 ( 
.A(n_960),
.B(n_812),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_955),
.B(n_868),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_962),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_964),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_965),
.B(n_947),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_966),
.B(n_778),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_963),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_967),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_963),
.A2(n_923),
.B1(n_951),
.B2(n_925),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_964),
.B(n_953),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_964),
.B(n_953),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_966),
.A2(n_785),
.B(n_868),
.C(n_846),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_951),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_973),
.B(n_790),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_933),
.Y(n_980)
);

OAI322xp33_ASAP7_75t_L g981 ( 
.A1(n_968),
.A2(n_974),
.A3(n_972),
.B1(n_969),
.B2(n_976),
.C1(n_975),
.C2(n_941),
.Y(n_981)
);

NOR4xp75_ASAP7_75t_L g982 ( 
.A(n_969),
.B(n_896),
.C(n_933),
.D(n_901),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_977),
.B(n_933),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_971),
.A2(n_875),
.B(n_941),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_948),
.B(n_855),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_985),
.B(n_979),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_983),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_980),
.B(n_948),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_981),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_982),
.Y(n_991)
);

INVxp33_ASAP7_75t_L g992 ( 
.A(n_984),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_937),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_918),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_993),
.Y(n_995)
);

AOI221xp5_ASAP7_75t_L g996 ( 
.A1(n_990),
.A2(n_918),
.B1(n_904),
.B2(n_921),
.C(n_876),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

AOI211xp5_ASAP7_75t_L g998 ( 
.A1(n_988),
.A2(n_846),
.B(n_869),
.C(n_786),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_SL g999 ( 
.A1(n_991),
.A2(n_869),
.B1(n_921),
.B2(n_816),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_987),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_994),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_1000),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_995),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_999),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_998),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_996),
.Y(n_1007)
);

INVxp33_ASAP7_75t_SL g1008 ( 
.A(n_1000),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_994),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_994),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_994),
.Y(n_1011)
);

NAND4xp25_ASAP7_75t_L g1012 ( 
.A(n_1006),
.B(n_992),
.C(n_791),
.D(n_817),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_1005),
.B(n_803),
.C(n_824),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_1009),
.B(n_921),
.Y(n_1015)
);

AOI211x1_ASAP7_75t_L g1016 ( 
.A1(n_1007),
.A2(n_863),
.B(n_906),
.C(n_855),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1010),
.Y(n_1017)
);

NAND4xp75_ASAP7_75t_L g1018 ( 
.A(n_1002),
.B(n_1004),
.C(n_1011),
.D(n_1001),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1003),
.Y(n_1019)
);

AOI211x1_ASAP7_75t_L g1020 ( 
.A1(n_1008),
.A2(n_910),
.B(n_902),
.C(n_907),
.Y(n_1020)
);

OAI211xp5_ASAP7_75t_SL g1021 ( 
.A1(n_1006),
.A2(n_809),
.B(n_833),
.C(n_818),
.Y(n_1021)
);

XNOR2x1_ASAP7_75t_SL g1022 ( 
.A(n_1002),
.B(n_867),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1022),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_L g1024 ( 
.A(n_1013),
.B(n_887),
.C(n_891),
.Y(n_1024)
);

NAND4xp25_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_891),
.C(n_887),
.D(n_801),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1017),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1019),
.B(n_822),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1012),
.B(n_822),
.C(n_839),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_1014),
.B(n_822),
.C(n_819),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_1023),
.A2(n_1021),
.B(n_1018),
.C(n_1016),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_1027),
.A2(n_1020),
.B(n_940),
.Y(n_1031)
);

CKINVDCx6p67_ASAP7_75t_R g1032 ( 
.A(n_1026),
.Y(n_1032)
);

NAND4xp25_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1024),
.C(n_1028),
.D(n_1025),
.Y(n_1033)
);

NAND4xp25_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_891),
.C(n_887),
.D(n_871),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1026),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_1026),
.B(n_891),
.C(n_887),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_940),
.B(n_939),
.C(n_931),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_1026),
.B(n_939),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_1035),
.B(n_931),
.Y(n_1039)
);

NAND4xp75_ASAP7_75t_L g1040 ( 
.A(n_1038),
.B(n_930),
.C(n_864),
.D(n_871),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

OAI22x1_ASAP7_75t_SL g1042 ( 
.A1(n_1030),
.A2(n_930),
.B1(n_864),
.B2(n_870),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1036),
.A2(n_867),
.B1(n_870),
.B2(n_893),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_L g1044 ( 
.A(n_1033),
.B(n_870),
.Y(n_1044)
);

AO22x2_ASAP7_75t_L g1045 ( 
.A1(n_1031),
.A2(n_867),
.B1(n_915),
.B2(n_913),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_1034),
.B(n_842),
.Y(n_1046)
);

NAND4xp75_ASAP7_75t_L g1047 ( 
.A(n_1037),
.B(n_865),
.C(n_902),
.D(n_907),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_1041),
.B(n_837),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1049)
);

OR3x1_ASAP7_75t_L g1050 ( 
.A(n_1042),
.B(n_910),
.C(n_879),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_1039),
.B(n_858),
.C(n_859),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1043),
.B(n_895),
.C(n_170),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_858),
.C(n_859),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1045),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1047),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1041),
.B(n_915),
.Y(n_1056)
);

AOI31xp33_ASAP7_75t_L g1057 ( 
.A1(n_1044),
.A2(n_895),
.A3(n_911),
.B(n_842),
.Y(n_1057)
);

OAI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_1041),
.A2(n_911),
.B1(n_908),
.B2(n_915),
.C(n_914),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1041),
.B(n_914),
.Y(n_1059)
);

NOR4xp25_ASAP7_75t_L g1060 ( 
.A(n_1041),
.B(n_914),
.C(n_913),
.D(n_912),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1056),
.B(n_914),
.Y(n_1061)
);

XNOR2xp5_ASAP7_75t_L g1062 ( 
.A(n_1049),
.B(n_168),
.Y(n_1062)
);

AOI211xp5_ASAP7_75t_L g1063 ( 
.A1(n_1055),
.A2(n_908),
.B(n_175),
.C(n_176),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1054),
.B(n_913),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1048),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1059),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1052),
.A2(n_876),
.B1(n_897),
.B2(n_890),
.C(n_885),
.Y(n_1067)
);

XOR2xp5_ASAP7_75t_L g1068 ( 
.A(n_1050),
.B(n_171),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_1057),
.A2(n_909),
.B(n_897),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1068),
.A2(n_1053),
.B1(n_1058),
.B2(n_1051),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_SL g1072 ( 
.A1(n_1062),
.A2(n_1060),
.B1(n_909),
.B2(n_890),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1066),
.A2(n_909),
.B1(n_876),
.B2(n_829),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_1065),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1063),
.A2(n_829),
.B1(n_885),
.B2(n_882),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1074),
.B(n_1070),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1071),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1075),
.A2(n_1064),
.B1(n_1067),
.B2(n_1069),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1076),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1079),
.Y(n_1080)
);

AOI222xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1080),
.A2(n_1077),
.B1(n_1078),
.B2(n_1072),
.C1(n_1073),
.C2(n_181),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_L g1082 ( 
.A(n_1081),
.B(n_177),
.C(n_178),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1081),
.A2(n_882),
.B1(n_879),
.B2(n_878),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1082),
.B(n_179),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1083),
.B(n_180),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_1084),
.B(n_182),
.Y(n_1086)
);

OAI221xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1085),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.C(n_878),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_1087),
.A2(n_854),
.B1(n_853),
.B2(n_848),
.C(n_843),
.Y(n_1088)
);

AOI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1088),
.A2(n_1086),
.B(n_862),
.C(n_852),
.Y(n_1089)
);


endmodule