module fake_jpeg_1079_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_0),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_41),
.B(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_50),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_28),
.B(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_28),
.B(n_9),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_58),
.B1(n_72),
.B2(n_46),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_16),
.C(n_32),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_42),
.B1(n_52),
.B2(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_32),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_17),
.B(n_16),
.C(n_4),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_74),
.B(n_15),
.C(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_34),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_23),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

XNOR2x2_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_70),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_35),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_97),
.B(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_98),
.Y(n_112)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_101),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_46),
.B1(n_37),
.B2(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_0),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_64),
.B(n_68),
.C(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_0),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_61),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_62),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_61),
.C(n_79),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_117),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_115),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_70),
.B(n_68),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_120),
.B(n_102),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_65),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_79),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_95),
.C(n_91),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_39),
.B(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_2),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_87),
.B(n_82),
.Y(n_136)
);

NOR4xp25_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_80),
.C(n_83),
.D(n_81),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_122),
.B(n_117),
.C(n_121),
.D(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_96),
.B1(n_80),
.B2(n_81),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_135),
.B1(n_105),
.B2(n_121),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_86),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.C(n_132),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_99),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_90),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_133),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_100),
.B(n_85),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_138),
.B(n_122),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_136),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_102),
.C(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_145),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_107),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_75),
.B1(n_5),
.B2(n_6),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_119),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_130),
.C(n_104),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

AO221x1_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_114),
.B1(n_113),
.B2(n_104),
.C(n_137),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

OAI321xp33_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_130),
.A3(n_132),
.B1(n_133),
.B2(n_113),
.C(n_114),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_158),
.B1(n_160),
.B2(n_149),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_146),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_75),
.B1(n_71),
.B2(n_6),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_159),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_141),
.C(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_167),
.B1(n_169),
.B2(n_163),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_143),
.B1(n_141),
.B2(n_145),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_156),
.B1(n_151),
.B2(n_162),
.Y(n_174)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_159),
.B(n_157),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_8),
.B(n_171),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_173),
.A2(n_161),
.B(n_7),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_169),
.C(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_170),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_178),
.B(n_177),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_8),
.Y(n_182)
);


endmodule