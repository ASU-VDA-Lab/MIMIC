module fake_jpeg_22298_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_17),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_52),
.B(n_17),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_9),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_67),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_34),
.B1(n_39),
.B2(n_31),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_28),
.C(n_18),
.Y(n_104)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_71),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_26),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_39),
.B1(n_31),
.B2(n_20),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_81),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_36),
.B1(n_32),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_90),
.Y(n_152)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_30),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_27),
.B1(n_37),
.B2(n_35),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_28),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_117),
.B(n_119),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_120),
.B(n_38),
.C(n_22),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_57),
.B(n_51),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_28),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_28),
.C(n_50),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_62),
.C(n_50),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_21),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_30),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_65),
.Y(n_136)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_76),
.B1(n_68),
.B2(n_66),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_143),
.B1(n_99),
.B2(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_132),
.Y(n_186)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_139),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_138),
.C(n_104),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_65),
.C(n_23),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_99),
.B1(n_123),
.B2(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_100),
.B(n_38),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_147),
.Y(n_192)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_24),
.B1(n_33),
.B2(n_29),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_95),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_24),
.B1(n_33),
.B2(n_29),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_26),
.B1(n_25),
.B2(n_35),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_25),
.B(n_10),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_13),
.C(n_16),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_111),
.B(n_115),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_173),
.B(n_180),
.C(n_1),
.D(n_4),
.Y(n_220)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_166),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_184),
.B1(n_147),
.B2(n_141),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_93),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_176),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_126),
.A2(n_117),
.B1(n_91),
.B2(n_87),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_132),
.C(n_110),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_117),
.B(n_91),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_119),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_190),
.B1(n_137),
.B2(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_135),
.B(n_120),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_101),
.B1(n_103),
.B2(n_114),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_143),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_12),
.B(n_15),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_107),
.B1(n_110),
.B2(n_3),
.Y(n_190)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_198),
.B1(n_200),
.B2(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_215),
.B1(n_191),
.B2(n_175),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_149),
.B1(n_154),
.B2(n_124),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_146),
.B1(n_127),
.B2(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_169),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_176),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_209),
.C(n_213),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_224),
.B(n_181),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_130),
.B1(n_134),
.B2(n_0),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_173),
.B(n_180),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_194),
.B(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_130),
.C(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_9),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_220),
.C(n_179),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_1),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_191),
.B1(n_161),
.B2(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_237),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_238),
.B(n_242),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_244),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_195),
.B1(n_223),
.B2(n_198),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_204),
.B(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_162),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_246),
.C(n_220),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_165),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_182),
.C(n_170),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_166),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_6),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_185),
.B1(n_193),
.B2(n_8),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_222),
.B1(n_185),
.B2(n_204),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_210),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_258),
.C(n_260),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_215),
.B1(n_232),
.B2(n_241),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_246),
.C(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

NOR4xp25_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_208),
.C(n_213),
.D(n_196),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_264),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_227),
.A2(n_238),
.B1(n_237),
.B2(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_233),
.B1(n_249),
.B2(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_217),
.C(n_201),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_277),
.B1(n_286),
.B2(n_11),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_281),
.B1(n_283),
.B2(n_287),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_248),
.B(n_218),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_248),
.B1(n_214),
.B2(n_9),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_6),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_258),
.C(n_254),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_260),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

FAx1_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_265),
.CI(n_251),
.CON(n_291),
.SN(n_291)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_275),
.B(n_282),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_256),
.C(n_257),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.C(n_299),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_256),
.C(n_257),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_276),
.C(n_271),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_14),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_285),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_291),
.C(n_286),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_305),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_270),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_298),
.C(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.C(n_284),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_16),
.B1(n_291),
.B2(n_304),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_281),
.C(n_270),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_296),
.B1(n_292),
.B2(n_290),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_319),
.C(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_272),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_277),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_306),
.B(n_16),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_319),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_321),
.B(n_327),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_315),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_314),
.C(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_330),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_326),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_329),
.Y(n_334)
);


endmodule