module fake_jpeg_26148_n_68 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_11),
.B(n_22),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2x1_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_0),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_9),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_23),
.B(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_2),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_3),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_19),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_6),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_54),
.C(n_59),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_5),
.B1(n_15),
.B2(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_56),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_52),
.C(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_57),
.Y(n_68)
);


endmodule