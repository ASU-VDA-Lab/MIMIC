module fake_aes_30_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NOR2xp33_ASAP7_75t_L g4 ( .A(n_1), .B(n_2), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
AOI221xp5_ASAP7_75t_SL g7 ( .A1(n_3), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_4), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
AOI21xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .B(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_3), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_12), .B(n_10), .Y(n_14) );
OAI21xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_13), .B(n_10), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_15), .B(n_14), .Y(n_16) );
endmodule