module fake_jpeg_17653_n_44 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_1),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g26 ( 
.A(n_5),
.B(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_15),
.B1(n_14),
.B2(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_24),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_23),
.Y(n_38)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.A3(n_18),
.B1(n_35),
.B2(n_13),
.C(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_16),
.CI(n_18),
.CON(n_43),
.SN(n_43)
);

OAI31xp33_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_35),
.A3(n_41),
.B(n_40),
.Y(n_44)
);


endmodule