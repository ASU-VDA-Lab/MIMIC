module fake_jpeg_30144_n_437 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_14),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_46),
.B(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_60),
.Y(n_98)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_72),
.Y(n_107)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_74),
.Y(n_131)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_80),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_77),
.Y(n_130)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_79),
.Y(n_138)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_82),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_41),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_33),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_89),
.B(n_43),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_44),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_94),
.B(n_116),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_129),
.Y(n_179)
);

BUFx2_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_30),
.B1(n_17),
.B2(n_45),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_114),
.B1(n_117),
.B2(n_50),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_30),
.B1(n_45),
.B2(n_41),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_45),
.B1(n_22),
.B2(n_32),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_136),
.B1(n_43),
.B2(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_22),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_44),
.B1(n_23),
.B2(n_41),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_20),
.B1(n_36),
.B2(n_40),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_125),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_64),
.A2(n_44),
.B(n_41),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_27),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_27),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_36),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_32),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_43),
.B1(n_37),
.B2(n_28),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_58),
.B(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_159),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_91),
.B1(n_61),
.B2(n_75),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_158),
.B(n_106),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_64),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_162),
.Y(n_200)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_139),
.B(n_100),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_78),
.B1(n_72),
.B2(n_67),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_164),
.A2(n_175),
.B1(n_181),
.B2(n_186),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_63),
.B1(n_40),
.B2(n_44),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_180),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_44),
.B1(n_41),
.B2(n_23),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_191),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_173),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_122),
.B(n_2),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_183),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_97),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_185),
.Y(n_230)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_96),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_192),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_94),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_193),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_111),
.A2(n_10),
.B1(n_11),
.B2(n_115),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_122),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_221),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_102),
.B(n_127),
.C(n_113),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_196),
.A2(n_231),
.B(n_184),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_154),
.B(n_132),
.CI(n_113),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_202),
.B(n_139),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_190),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_138),
.C(n_132),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_226),
.C(n_183),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_217),
.B(n_232),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_156),
.A2(n_138),
.B(n_140),
.C(n_135),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_159),
.B(n_135),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_156),
.A2(n_152),
.B1(n_169),
.B2(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_229),
.B1(n_164),
.B2(n_186),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_225),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_100),
.C(n_103),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_99),
.B1(n_106),
.B2(n_103),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_143),
.B1(n_153),
.B2(n_192),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_158),
.A2(n_118),
.B1(n_112),
.B2(n_108),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_159),
.A2(n_113),
.B(n_139),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_143),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_112),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_206),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_238),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_239),
.A2(n_244),
.B1(n_268),
.B2(n_211),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_247),
.B1(n_224),
.B2(n_227),
.Y(n_282)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_212),
.B(n_210),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_246),
.B(n_253),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_203),
.B1(n_210),
.B2(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_252),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_157),
.B(n_151),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_202),
.A2(n_158),
.B1(n_162),
.B2(n_145),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_248),
.B(n_274),
.Y(n_279)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_197),
.A2(n_179),
.A3(n_175),
.B1(n_99),
.B2(n_176),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_214),
.Y(n_286)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_187),
.B1(n_150),
.B2(n_120),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_185),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

NAND2x1_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_139),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_118),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_134),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_225),
.B(n_134),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_265),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_201),
.B(n_199),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_267),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_210),
.A2(n_148),
.B1(n_155),
.B2(n_161),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_182),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_200),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_200),
.B(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_198),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_218),
.A2(n_232),
.B(n_236),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_243),
.A2(n_214),
.B(n_229),
.C(n_196),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_276),
.A2(n_252),
.B(n_261),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_226),
.C(n_222),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_293),
.C(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_199),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_299),
.C(n_256),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_260),
.C(n_241),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_237),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_215),
.C(n_198),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_253),
.B(n_215),
.C(n_221),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_234),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_256),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_194),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_306),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_240),
.A2(n_204),
.B1(n_211),
.B2(n_195),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_239),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_216),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_242),
.C(n_269),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_247),
.B1(n_261),
.B2(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_311),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_SL g344 ( 
.A1(n_313),
.A2(n_276),
.B(n_308),
.C(n_266),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_289),
.B(n_270),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_314),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_316),
.Y(n_338)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_321),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_323),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g320 ( 
.A(n_296),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_291),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_325),
.B1(n_268),
.B2(n_292),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_273),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_306),
.B(n_281),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_324),
.A2(n_335),
.B(n_337),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_271),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_328),
.C(n_331),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_246),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_330),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_291),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_332),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_237),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_248),
.B1(n_267),
.B2(n_275),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_292),
.B1(n_276),
.B2(n_290),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_277),
.A2(n_257),
.B(n_272),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_279),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_336),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_251),
.B(n_266),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_347),
.B(n_313),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_284),
.B1(n_282),
.B2(n_295),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_345),
.A2(n_350),
.B1(n_322),
.B2(n_310),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_320),
.A2(n_295),
.B(n_276),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_284),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_359),
.Y(n_362)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_302),
.B(n_287),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_349),
.B(n_319),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_320),
.A2(n_300),
.B1(n_276),
.B2(n_302),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_351),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_328),
.C(n_283),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_356),
.C(n_361),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_358),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_290),
.C(n_298),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_332),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_287),
.C(n_303),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_363),
.A2(n_344),
.B(n_352),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_365),
.B1(n_358),
.B2(n_341),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_345),
.A2(n_310),
.B1(n_311),
.B2(n_329),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_323),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_367),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_331),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_335),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_316),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_372),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_329),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_380),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_249),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_376),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_334),
.B1(n_337),
.B2(n_305),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_352),
.B1(n_354),
.B2(n_341),
.Y(n_386)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_312),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_301),
.C(n_250),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_361),
.C(n_354),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_342),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_389),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_385),
.A2(n_379),
.B1(n_344),
.B2(n_369),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_386),
.A2(n_364),
.B1(n_377),
.B2(n_370),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_390),
.B(n_391),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_347),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_394),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_338),
.C(n_346),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_397),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_365),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_382),
.B(n_362),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_401),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_396),
.B(n_343),
.Y(n_401)
);

OAI321xp33_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_379),
.A3(n_377),
.B1(n_363),
.B2(n_376),
.C(n_373),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_402),
.A2(n_405),
.B1(n_385),
.B2(n_388),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_371),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_389),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_343),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_406),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_378),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_387),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_409),
.A2(n_393),
.B1(n_383),
.B2(n_305),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_414),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_412),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_378),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_390),
.B(n_258),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_415),
.A2(n_417),
.B(n_413),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_403),
.A2(n_266),
.B1(n_255),
.B2(n_259),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_409),
.C(n_408),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_398),
.A2(n_238),
.B(n_384),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_418),
.B(n_419),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_425),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_415),
.A2(n_399),
.B(n_398),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_423),
.A2(n_238),
.B(n_195),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_387),
.C(n_216),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_418),
.C(n_235),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_427),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_429),
.B(n_238),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_422),
.B(n_238),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_430),
.A2(n_421),
.B(n_424),
.Y(n_432)
);

O2A1O1Ixp5_ASAP7_75t_SL g435 ( 
.A1(n_434),
.A2(n_432),
.B(n_424),
.C(n_433),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_204),
.B(n_208),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_208),
.B(n_204),
.Y(n_437)
);


endmodule