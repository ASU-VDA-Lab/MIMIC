module fake_ariane_119_n_122 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_122);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_122;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_117;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_112;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

AOI22x1_ASAP7_75t_SL g41 ( 
.A1(n_25),
.A2(n_10),
.B1(n_30),
.B2(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_1),
.Y(n_50)
);

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_16),
.B(n_3),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_11),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_14),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_17),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_18),
.C(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_38),
.B(n_50),
.C(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_41),
.B1(n_34),
.B2(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_63),
.Y(n_73)
);

OAI21x1_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_35),
.B(n_64),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_51),
.B(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_51),
.B(n_41),
.C(n_43),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_48),
.B(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_48),
.B1(n_43),
.B2(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_61),
.B1(n_56),
.B2(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_39),
.B(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_45),
.B(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_69),
.B1(n_78),
.B2(n_80),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_81),
.B1(n_98),
.B2(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_100),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_94),
.B1(n_92),
.B2(n_87),
.Y(n_105)
);

XOR2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_81),
.Y(n_106)
);

NOR2x1_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_102),
.Y(n_111)
);

NOR4xp25_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_79),
.C(n_91),
.D(n_85),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_94),
.B1(n_45),
.B2(n_96),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_96),
.B1(n_45),
.B2(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_115),
.B1(n_86),
.B2(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_107),
.B1(n_91),
.B2(n_47),
.Y(n_119)
);

AOI31xp33_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_60),
.A3(n_46),
.B(n_47),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_39),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_46),
.B1(n_47),
.B2(n_89),
.C(n_121),
.Y(n_122)
);


endmodule