module real_jpeg_17901_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_445),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_0),
.B(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_1),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_62),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_1),
.B(n_296),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_1),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_1),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_1),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_3),
.B(n_58),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_3),
.B(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_4),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_4),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_5),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_5),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_5),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_6),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_8),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_8),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_8),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_8),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_8),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_8),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_9),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_9),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_9),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_9),
.B(n_373),
.Y(n_372)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_10),
.Y(n_92)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_10),
.Y(n_418)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_11),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_17),
.B1(n_41),
.B2(n_45),
.Y(n_40)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_12),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_12),
.B(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_14),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_14),
.B(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_14),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_17),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_17),
.B(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_402),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_214),
.B(n_400),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_166),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_23),
.B(n_166),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_102),
.C(n_142),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_24),
.A2(n_25),
.B1(n_102),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_65),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_39),
.C(n_50),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_27),
.B(n_51),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_32),
.C(n_35),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_35),
.B(n_198),
.Y(n_240)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

XNOR2x1_ASAP7_75t_SL g248 ( 
.A(n_38),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_40),
.A2(n_273),
.B(n_275),
.Y(n_272)
);

XOR2x2_ASAP7_75t_SL g388 ( 
.A(n_40),
.B(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_43),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_45),
.Y(n_274)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_47),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_49),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_49),
.Y(n_442)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_61),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_52),
.B(n_61),
.Y(n_145)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_56),
.B(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_79),
.B1(n_100),
.B2(n_101),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_73),
.B(n_76),
.C(n_78),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_86),
.C(n_97),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_80),
.A2(n_83),
.B1(n_98),
.B2(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_82),
.Y(n_362)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_86),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_93),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_87),
.A2(n_93),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_87),
.Y(n_281)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_91),
.B(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_93),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_93),
.Y(n_282)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_168),
.C(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_102),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_132),
.C(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_104),
.B(n_108),
.C(n_112),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_111),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_114),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_132),
.Y(n_115)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_117),
.B(n_124),
.C(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_118),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_118),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_131),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_124),
.A2(n_125),
.B1(n_148),
.B2(n_149),
.Y(n_226)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_127),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_128),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_129),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_129),
.A2(n_131),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_129),
.B(n_256),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_130),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_131),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_131),
.B(n_193),
.C(n_198),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_138),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_134),
.B1(n_138),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_136),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_135),
.A2(n_136),
.B1(n_430),
.B2(n_434),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_142),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_158),
.C(n_163),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_143),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_151),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_144),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_150),
.Y(n_375)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_151),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_152),
.A2(n_155),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_153),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_155),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_155),
.A2(n_198),
.B1(n_200),
.B2(n_224),
.Y(n_436)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_157),
.Y(n_303)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_159),
.B(n_164),
.Y(n_386)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_167),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_191),
.B1(n_212),
.B2(n_213),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_190),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_172),
.B(n_176),
.C(n_189),
.Y(n_407)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_189),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_181),
.B(n_184),
.C(n_188),
.Y(n_413)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_185),
.B(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_191),
.B(n_212),
.C(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_201),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_192),
.B(n_202),
.C(n_203),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_211),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_205),
.B(n_211),
.C(n_282),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_382),
.B(n_397),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_283),
.B(n_381),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_261),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_218),
.B(n_261),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_239),
.C(n_247),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_219),
.A2(n_220),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_226),
.C(n_227),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_235),
.Y(n_305)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_239),
.B(n_247),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.C(n_255),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_255),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_263),
.B(n_268),
.C(n_269),
.Y(n_391)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_270),
.B(n_272),
.C(n_279),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21x1_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_309),
.B(n_380),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_306),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_285),
.B(n_306),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_304),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_304),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.C(n_301),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_314),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_301),
.Y(n_314)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_328),
.B(n_379),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_326),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_311),
.B(n_326),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.C(n_324),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_312),
.A2(n_313),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_324),
.B1(n_325),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_315),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_342),
.B(n_378),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_338),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_330),
.B(n_338),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.C(n_336),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_355),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_336),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_339),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_357),
.B(n_377),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_354),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_344),
.B(n_354),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_351),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_351),
.Y(n_363)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_364),
.B(n_376),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_359),
.B(n_363),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_372),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_391),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_391),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_388),
.C(n_390),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

OAI21x1_ASAP7_75t_SL g397 ( 
.A1(n_392),
.A2(n_398),
.B(n_399),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_394),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_443),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_406),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_423),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_422),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

AO22x1_ASAP7_75t_SL g414 ( 
.A1(n_415),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_414)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_415),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_419),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_435),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_430),
.Y(n_434)
);

INVx5_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);


endmodule