module fake_jpeg_14561_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_42),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_28),
.B1(n_32),
.B2(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_45),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_21),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_65),
.B1(n_73),
.B2(n_47),
.Y(n_80)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_66),
.B1(n_28),
.B2(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_35),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_48),
.B1(n_40),
.B2(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_0),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_28),
.B1(n_22),
.B2(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_27),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_71),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_34),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_20),
.B1(n_30),
.B2(n_17),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_77),
.Y(n_118)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_100),
.B1(n_23),
.B2(n_61),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_93),
.B1(n_71),
.B2(n_69),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_20),
.B1(n_43),
.B2(n_36),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_98),
.B(n_24),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_36),
.B1(n_43),
.B2(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_101),
.B1(n_65),
.B2(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_23),
.B1(n_22),
.B2(n_38),
.Y(n_98)
);

OA22x2_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_38),
.B1(n_44),
.B2(n_46),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_46),
.B1(n_23),
.B2(n_22),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_46),
.B1(n_34),
.B2(n_26),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_55),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_83),
.B(n_88),
.C(n_87),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_105),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_68),
.C(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_119),
.B1(n_84),
.B2(n_91),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_68),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_67),
.B1(n_53),
.B2(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_53),
.B1(n_51),
.B2(n_72),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_127),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_132),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_57),
.C(n_63),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_61),
.B1(n_62),
.B2(n_51),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_54),
.B1(n_19),
.B2(n_18),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_91),
.B1(n_76),
.B2(n_84),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_74),
.A2(n_66),
.B(n_73),
.C(n_18),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_66),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_24),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_19),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_97),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_79),
.A2(n_49),
.B1(n_34),
.B2(n_26),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_117),
.B1(n_119),
.B2(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_141),
.B1(n_145),
.B2(n_154),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_139),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_82),
.B(n_81),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_157),
.B(n_159),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_153),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_102),
.B1(n_90),
.B2(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_94),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_79),
.B1(n_100),
.B2(n_99),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_163),
.B1(n_132),
.B2(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_131),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_126),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_99),
.B1(n_100),
.B2(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_160),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_84),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_116),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_76),
.B1(n_96),
.B2(n_85),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_166),
.A2(n_178),
.B1(n_190),
.B2(n_157),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_108),
.B(n_105),
.C(n_106),
.D(n_130),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_171),
.B(n_128),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_116),
.C(n_108),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_176),
.C(n_184),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_122),
.C(n_105),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_129),
.B1(n_113),
.B2(n_119),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_183),
.Y(n_214)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_111),
.C(n_103),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_157),
.C(n_140),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_138),
.A2(n_106),
.B1(n_129),
.B2(n_103),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_106),
.B(n_118),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_159),
.B(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_118),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_140),
.B1(n_150),
.B2(n_155),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_155),
.B1(n_145),
.B2(n_133),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_201),
.A2(n_224),
.B1(n_169),
.B2(n_26),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_146),
.B(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_211),
.C(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_168),
.B1(n_181),
.B2(n_186),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_141),
.B(n_133),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_195),
.B(n_174),
.C(n_186),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_R g209 ( 
.A1(n_190),
.A2(n_154),
.B(n_152),
.C(n_149),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_179),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_163),
.C(n_153),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_144),
.B1(n_139),
.B2(n_135),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_136),
.B1(n_77),
.B2(n_75),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_77),
.B1(n_75),
.B2(n_101),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_220),
.B1(n_222),
.B2(n_182),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_70),
.C(n_49),
.Y(n_219)
);

XOR2x2_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_44),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_31),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_184),
.C(n_179),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_164),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_185),
.A2(n_34),
.B1(n_26),
.B2(n_29),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_231),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_226),
.A2(n_245),
.B1(n_213),
.B2(n_196),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_168),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_242),
.C(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_232),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_248),
.B1(n_249),
.B2(n_224),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_29),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_174),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_243),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_188),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_167),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_205),
.B1(n_216),
.B2(n_218),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_172),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_3),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_193),
.C(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_177),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_204),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_177),
.B1(n_169),
.B2(n_2),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_208),
.A2(n_169),
.B(n_49),
.C(n_70),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_24),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_31),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_221),
.C(n_31),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_253),
.B1(n_259),
.B2(n_267),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_200),
.B1(n_211),
.B2(n_206),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_263),
.C(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_201),
.B1(n_219),
.B2(n_215),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_270),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_217),
.B(n_222),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_249),
.B(n_250),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_229),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_29),
.C(n_24),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_24),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_269),
.C(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_44),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_1),
.C(n_3),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_226),
.B(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_233),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_285),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_266),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_247),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_229),
.B(n_233),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_242),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_249),
.B(n_268),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_252),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_287),
.B(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_249),
.C(n_4),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_273),
.C(n_267),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_292),
.B1(n_4),
.B2(n_5),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_3),
.B(n_4),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_253),
.B1(n_259),
.B2(n_256),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_280),
.B1(n_9),
.B2(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_304),
.C(n_305),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_292),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_263),
.C(n_264),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_7),
.C(n_8),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_16),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_283),
.B(n_276),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.Y(n_325)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_290),
.B(n_278),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_317),
.B(n_9),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_285),
.B(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_278),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_316),
.B(n_320),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_280),
.B(n_277),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_304),
.A3(n_298),
.B1(n_295),
.B2(n_302),
.C1(n_300),
.C2(n_306),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_321),
.B(n_322),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_303),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_308),
.B1(n_311),
.B2(n_310),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_327)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_334),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_311),
.B(n_310),
.C(n_315),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_336),
.B(n_324),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_11),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_15),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_337),
.B(n_330),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_339),
.A2(n_341),
.B(n_342),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_327),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_340),
.B(n_331),
.CI(n_325),
.CON(n_344),
.SN(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_335),
.B(n_338),
.C(n_15),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_343),
.C(n_15),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_15),
.Y(n_347)
);


endmodule