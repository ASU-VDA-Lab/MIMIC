module fake_aes_1820_n_864 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_864);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_864;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_21), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_70), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_16), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_89), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_48), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_102), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_65), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_59), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_49), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_98), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_56), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_57), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_8), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_74), .B(n_28), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_19), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_20), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_78), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_36), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_1), .Y(n_135) );
XOR2xp5_ASAP7_75t_L g136 ( .A(n_94), .B(n_12), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_12), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_101), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_47), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_58), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_126), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_111), .A2(n_43), .B(n_99), .Y(n_143) );
CKINVDCx8_ASAP7_75t_R g144 ( .A(n_138), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_126), .Y(n_145) );
BUFx12f_ASAP7_75t_L g146 ( .A(n_118), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVxp33_ASAP7_75t_SL g149 ( .A(n_117), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_109), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_118), .B(n_0), .Y(n_152) );
BUFx12f_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_103), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_126), .B(n_2), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_107), .B(n_3), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_110), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_110), .B(n_3), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_121), .B(n_4), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_113), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_113), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_116), .B(n_45), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_116), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_127), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
OR2x6_ASAP7_75t_L g166 ( .A(n_152), .B(n_128), .Y(n_166) );
BUFx10_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_158), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_146), .B(n_152), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_146), .B(n_106), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_147), .B(n_108), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_150), .A2(n_135), .B1(n_137), .B2(n_139), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_141), .B(n_105), .C(n_112), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_145), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_155), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_147), .B(n_108), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx1_ASAP7_75t_SL g184 ( .A(n_149), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_146), .B(n_114), .Y(n_187) );
NAND2xp33_ASAP7_75t_L g188 ( .A(n_162), .B(n_114), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_154), .B(n_141), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_155), .B(n_115), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_154), .B(n_115), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_144), .B(n_119), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_153), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_152), .B(n_136), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_148), .B(n_122), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_148), .B(n_122), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_151), .B(n_123), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_143), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_155), .B(n_127), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_151), .B(n_123), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_158), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_160), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_157), .B(n_153), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_190), .B(n_153), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_167), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_181), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_183), .A2(n_156), .B(n_159), .C(n_164), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_190), .B(n_144), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_167), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_174), .B(n_144), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_185), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_184), .B(n_195), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_196), .B(n_157), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g223 ( .A(n_188), .B(n_150), .C(n_156), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_200), .B(n_157), .Y(n_225) );
BUFx8_ASAP7_75t_L g226 ( .A(n_182), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_181), .B(n_159), .Y(n_227) );
NAND2xp33_ASAP7_75t_L g228 ( .A(n_205), .B(n_162), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_204), .B(n_130), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_207), .B(n_130), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_170), .B(n_139), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_183), .B(n_120), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_182), .B(n_140), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g234 ( .A(n_179), .B(n_163), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_191), .B(n_140), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_166), .A2(n_136), .B1(n_162), .B2(n_160), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_206), .B(n_163), .Y(n_238) );
AO221x1_ASAP7_75t_L g239 ( .A1(n_177), .A2(n_163), .B1(n_164), .B2(n_160), .C(n_124), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_206), .B(n_163), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_206), .B(n_164), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_186), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_192), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_166), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_211), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_186), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_206), .B(n_164), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_183), .B(n_131), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_167), .B(n_165), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_165), .B(n_132), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_189), .B(n_164), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_193), .B(n_104), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_194), .B(n_162), .Y(n_253) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_172), .B(n_129), .C(n_134), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_166), .B(n_162), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_166), .B(n_162), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
BUFx12f_ASAP7_75t_L g258 ( .A(n_194), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_166), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_165), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_165), .B(n_162), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_259), .A2(n_195), .B1(n_208), .B2(n_168), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_259), .A2(n_195), .B1(n_208), .B2(n_168), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_215), .A2(n_168), .B(n_198), .C(n_201), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_227), .B(n_187), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_260), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_259), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_227), .B(n_195), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_258), .B(n_168), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_263), .A2(n_198), .B(n_201), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_228), .A2(n_198), .B(n_201), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_245), .B(n_198), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_215), .A2(n_201), .B(n_179), .C(n_210), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_228), .A2(n_176), .B(n_175), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_233), .B(n_203), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_203), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_244), .B(n_209), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_217), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_220), .B(n_202), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_218), .B(n_209), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_223), .B(n_202), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_255), .A2(n_180), .B(n_169), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_258), .B(n_202), .Y(n_286) );
AOI21xp33_ASAP7_75t_L g287 ( .A1(n_216), .A2(n_205), .B(n_199), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_250), .A2(n_205), .B(n_143), .Y(n_288) );
OAI321xp33_ASAP7_75t_L g289 ( .A1(n_237), .A2(n_133), .A3(n_134), .B1(n_199), .B2(n_197), .C(n_205), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_249), .A2(n_205), .B(n_143), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_212), .B(n_197), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_236), .B(n_162), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_241), .A2(n_133), .B(n_178), .C(n_176), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_250), .A2(n_256), .B(n_249), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_221), .A2(n_143), .B(n_178), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_225), .A2(n_143), .B(n_175), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_229), .B(n_162), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_226), .B(n_180), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_247), .A2(n_173), .B(n_180), .C(n_171), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_230), .B(n_173), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_262), .A2(n_171), .B(n_169), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_232), .A2(n_46), .B(n_97), .Y(n_304) );
BUFx4f_ASAP7_75t_SL g305 ( .A(n_269), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_270), .B(n_226), .Y(n_307) );
AOI21x1_ASAP7_75t_SL g308 ( .A1(n_292), .A2(n_240), .B(n_251), .Y(n_308) );
OAI21x1_ASAP7_75t_SL g309 ( .A1(n_304), .A2(n_257), .B(n_243), .Y(n_309) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_295), .A2(n_239), .B(n_232), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_290), .A2(n_248), .B(n_235), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_271), .Y(n_312) );
BUFx12f_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_270), .B(n_226), .Y(n_314) );
CKINVDCx14_ASAP7_75t_R g315 ( .A(n_271), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_SL g316 ( .A1(n_266), .A2(n_248), .B(n_213), .C(n_235), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_282), .B(n_261), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_285), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_267), .B(n_254), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_298), .B(n_213), .Y(n_320) );
O2A1O1Ixp5_ASAP7_75t_L g321 ( .A1(n_287), .A2(n_252), .B(n_231), .C(n_219), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_275), .A2(n_219), .B(n_222), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_297), .A2(n_224), .B(n_217), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_288), .A2(n_222), .B(n_246), .Y(n_324) );
AO21x1_ASAP7_75t_L g325 ( .A1(n_295), .A2(n_253), .B(n_246), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_273), .A2(n_224), .B(n_217), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_288), .A2(n_242), .B(n_224), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_272), .A2(n_242), .B(n_234), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_301), .B(n_4), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_276), .A2(n_44), .B(n_96), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_286), .B(n_5), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_327), .A2(n_296), .B(n_304), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_322), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_321), .A2(n_289), .B(n_294), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_315), .A2(n_264), .B1(n_265), .B2(n_274), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_306), .B(n_280), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_306), .B(n_280), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_327), .A2(n_296), .B(n_303), .Y(n_339) );
AOI21x1_ASAP7_75t_L g340 ( .A1(n_325), .A2(n_284), .B(n_303), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_309), .A2(n_300), .B(n_293), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_309), .A2(n_294), .B(n_302), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_324), .A2(n_278), .B(n_277), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_324), .A2(n_299), .B(n_281), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_322), .Y(n_345) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_325), .A2(n_283), .B(n_291), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_318), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_318), .A2(n_268), .B(n_50), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_311), .A2(n_308), .B(n_330), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_326), .A2(n_5), .A3(n_6), .B(n_7), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_279), .B(n_51), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_317), .B(n_279), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_319), .B(n_6), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_311), .A2(n_42), .B(n_95), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_328), .A2(n_41), .B(n_93), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
AOI21x1_ASAP7_75t_L g359 ( .A1(n_310), .A2(n_323), .B(n_320), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_347), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_357), .B(n_310), .Y(n_362) );
AO21x1_ASAP7_75t_SL g363 ( .A1(n_360), .A2(n_314), .B(n_307), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_350), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
NAND2x1_ASAP7_75t_L g367 ( .A(n_333), .B(n_310), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_337), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_350), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_334), .A2(n_331), .B(n_310), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_360), .B(n_312), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_312), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_335), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_358), .B(n_7), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_338), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_352), .B(n_9), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_333), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_356), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_332), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_352), .B(n_9), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_338), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_356), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_336), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_340), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_343), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_348), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_346), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_382), .B(n_359), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_387), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_398), .B(n_353), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_398), .B(n_343), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_361), .B(n_349), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_361), .B(n_349), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_401), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_365), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_365), .B(n_341), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_365), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_364), .B(n_341), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_364), .B(n_355), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_368), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_384), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_368), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_362), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_368), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_370), .B(n_355), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_370), .B(n_354), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_366), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_362), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_371), .B(n_354), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_371), .B(n_10), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_366), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_378), .B(n_11), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_378), .B(n_11), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_379), .B(n_13), .Y(n_451) );
OAI21x1_ASAP7_75t_L g452 ( .A1(n_403), .A2(n_351), .B(n_305), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_389), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_379), .B(n_14), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_403), .A2(n_55), .B(n_92), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_369), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_369), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_389), .B(n_15), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_393), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_381), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_393), .B(n_17), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_405), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_380), .B(n_17), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_369), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_405), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_405), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_406), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_380), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_396), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_383), .B(n_18), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_396), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_406), .B(n_22), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_374), .B(n_23), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_366), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_406), .B(n_408), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_408), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_374), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_383), .B(n_24), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_395), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_408), .B(n_25), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_399), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_399), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_386), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_376), .B(n_100), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_375), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_410), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_459), .B(n_394), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_424), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_412), .B(n_372), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_458), .B(n_394), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_412), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_413), .B(n_372), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_458), .B(n_394), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_468), .B(n_394), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_413), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_410), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_411), .B(n_385), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_415), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_410), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_460), .Y(n_507) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_426), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_478), .Y(n_509) );
INVx4_ASAP7_75t_L g510 ( .A(n_439), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
BUFx8_ASAP7_75t_L g512 ( .A(n_461), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_415), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_420), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_461), .B(n_385), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_428), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_446), .B(n_385), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_446), .B(n_385), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_428), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_430), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_376), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_449), .B(n_376), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_414), .A2(n_376), .B1(n_366), .B2(n_373), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_420), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_421), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_421), .B(n_372), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_425), .B(n_372), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_425), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_450), .B(n_373), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_439), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_435), .B(n_367), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_448), .B(n_373), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_435), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_436), .B(n_367), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_436), .B(n_402), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_478), .Y(n_536) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_417), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_450), .B(n_373), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_438), .B(n_374), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_451), .Y(n_540) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_433), .B(n_363), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_438), .B(n_392), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_454), .B(n_363), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_430), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_480), .B(n_392), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_433), .B(n_392), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_444), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_448), .B(n_386), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_443), .B(n_386), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_475), .Y(n_552) );
INVx4_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_443), .B(n_407), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_444), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_414), .B(n_377), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_463), .B(n_407), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_479), .B(n_407), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_470), .B(n_407), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_447), .B(n_377), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_429), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_429), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_447), .B(n_377), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_475), .B(n_375), .Y(n_564) );
INVx5_ASAP7_75t_L g565 ( .A(n_473), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_430), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_375), .Y(n_567) );
BUFx3_ASAP7_75t_L g568 ( .A(n_474), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_431), .B(n_407), .Y(n_569) );
AND2x4_ASAP7_75t_SL g570 ( .A(n_473), .B(n_407), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_469), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_473), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_431), .B(n_404), .Y(n_573) );
BUFx2_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_472), .B(n_404), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_427), .B(n_26), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_462), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_472), .B(n_27), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_416), .B(n_29), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_469), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_462), .B(n_30), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_434), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_465), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_416), .B(n_32), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_465), .B(n_34), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_434), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_466), .B(n_35), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_481), .B(n_37), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_418), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_481), .B(n_38), .Y(n_590) );
INVx5_ASAP7_75t_L g591 ( .A(n_417), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_471), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_427), .B(n_39), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_471), .Y(n_594) );
NAND2x1_ASAP7_75t_L g595 ( .A(n_510), .B(n_455), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_491), .B(n_434), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_544), .B(n_441), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_496), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_493), .B(n_466), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_495), .B(n_441), .Y(n_600) );
AND3x1_ASAP7_75t_L g601 ( .A(n_512), .B(n_453), .C(n_487), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_499), .B(n_445), .Y(n_602) );
AND2x4_ASAP7_75t_SL g603 ( .A(n_510), .B(n_482), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_541), .B(n_418), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_515), .B(n_445), .Y(n_605) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_507), .B(n_455), .Y(n_606) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_541), .A2(n_440), .B(n_432), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_501), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_540), .B(n_467), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_542), .B(n_467), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_521), .B(n_440), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_504), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_511), .Y(n_613) );
OR2x6_ASAP7_75t_L g614 ( .A(n_553), .B(n_455), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_552), .B(n_476), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_512), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_522), .B(n_432), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_513), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_556), .B(n_476), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_509), .A2(n_409), .B(n_482), .Y(n_620) );
AND2x4_ASAP7_75t_SL g621 ( .A(n_553), .B(n_483), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_556), .B(n_485), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_500), .B(n_485), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_514), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_545), .B(n_483), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_511), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_498), .B(n_418), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_498), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_530), .B(n_484), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_490), .B(n_422), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_528), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_524), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_525), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_506), .Y(n_634) );
NAND2x1_ASAP7_75t_L g635 ( .A(n_494), .B(n_455), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_549), .B(n_555), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_533), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_577), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_503), .B(n_40), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_577), .B(n_484), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_583), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_583), .B(n_457), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_562), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_517), .B(n_422), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_564), .B(n_486), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_573), .B(n_419), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_566), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_502), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_565), .B(n_536), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_518), .B(n_419), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_529), .B(n_418), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_573), .B(n_456), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_494), .B(n_409), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_586), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_568), .B(n_456), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_569), .B(n_409), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_532), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_564), .B(n_457), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_543), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_543), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_557), .B(n_409), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_538), .B(n_457), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_557), .B(n_486), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_532), .B(n_486), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_523), .B(n_464), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_535), .B(n_464), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_558), .A2(n_464), .B1(n_488), .B2(n_477), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_508), .B(n_488), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_520), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_535), .B(n_477), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_508), .B(n_477), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_558), .B(n_423), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_520), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_509), .B(n_423), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_489), .B(n_477), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_548), .B(n_423), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_568), .B(n_423), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_536), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_489), .B(n_477), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_547), .B(n_575), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_539), .B(n_477), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_546), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_550), .B(n_423), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_551), .B(n_423), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_546), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_505), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_492), .B(n_417), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_560), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_539), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_531), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_531), .Y(n_693) );
INVx4_ASAP7_75t_L g694 ( .A(n_565), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_516), .B(n_417), .Y(n_695) );
NAND2x1p5_ASAP7_75t_L g696 ( .A(n_578), .B(n_452), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_571), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_616), .Y(n_698) );
AND2x2_ASAP7_75t_SL g699 ( .A(n_603), .B(n_572), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_638), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_692), .B(n_527), .Y(n_701) );
OAI21xp33_ASAP7_75t_SL g702 ( .A1(n_604), .A2(n_590), .B(n_579), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_597), .B(n_574), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_634), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_693), .B(n_497), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_600), .B(n_589), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_661), .B(n_497), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_598), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_598), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_662), .B(n_527), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_602), .B(n_589), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_655), .B(n_534), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_599), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_690), .B(n_492), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_638), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_655), .B(n_534), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_641), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_680), .B(n_526), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_682), .B(n_526), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_642), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_647), .B(n_519), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_614), .B(n_590), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_694), .B(n_565), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_605), .B(n_554), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_659), .B(n_576), .Y(n_726) );
NAND2x2_ASAP7_75t_L g727 ( .A(n_601), .B(n_588), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_630), .B(n_658), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_619), .B(n_594), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_663), .B(n_563), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_641), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_623), .B(n_592), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_611), .B(n_563), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_608), .Y(n_734) );
INVx2_ASAP7_75t_SL g735 ( .A(n_621), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_612), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_617), .B(n_580), .Y(n_737) );
OAI21xp33_ASAP7_75t_L g738 ( .A1(n_607), .A2(n_559), .B(n_576), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_640), .B(n_567), .Y(n_739) );
INVx2_ASAP7_75t_SL g740 ( .A(n_628), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_622), .B(n_584), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_646), .B(n_593), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_618), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g744 ( .A(n_694), .B(n_565), .Y(n_744) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_613), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_624), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_645), .B(n_559), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_652), .B(n_570), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_615), .Y(n_749) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_639), .B(n_587), .C(n_585), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_631), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_637), .Y(n_752) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_614), .B(n_587), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_596), .B(n_585), .Y(n_754) );
AO21x1_ASAP7_75t_L g755 ( .A1(n_595), .A2(n_581), .B(n_570), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_653), .B(n_591), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_660), .B(n_581), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_637), .Y(n_758) );
INVxp33_ASAP7_75t_SL g759 ( .A(n_657), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_651), .B(n_591), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_629), .B(n_664), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_674), .B(n_591), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_691), .B(n_591), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_671), .Y(n_764) );
NAND2x1_ASAP7_75t_L g765 ( .A(n_606), .B(n_537), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_626), .Y(n_766) );
AOI322xp5_ASAP7_75t_L g767 ( .A1(n_620), .A2(n_537), .A3(n_417), .B1(n_452), .B2(n_60), .C1(n_61), .C2(n_62), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_671), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_727), .A2(n_667), .B1(n_665), .B2(n_666), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_720), .B(n_654), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_714), .B(n_632), .Y(n_771) );
O2A1O1Ixp5_ASAP7_75t_L g772 ( .A1(n_755), .A2(n_635), .B(n_609), .C(n_610), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_764), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_700), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_764), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_759), .A2(n_678), .B1(n_686), .B2(n_685), .Y(n_776) );
OR4x1_ASAP7_75t_L g777 ( .A(n_735), .B(n_644), .C(n_643), .D(n_633), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_768), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_749), .B(n_643), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_699), .Y(n_780) );
AOI222xp33_ASAP7_75t_L g781 ( .A1(n_698), .A2(n_636), .B1(n_625), .B2(n_644), .C1(n_656), .C2(n_648), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_704), .B(n_648), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_700), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_733), .B(n_627), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_716), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_740), .A2(n_696), .B1(n_669), .B2(n_627), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_716), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_718), .Y(n_788) );
AOI22x1_ASAP7_75t_L g789 ( .A1(n_744), .A2(n_679), .B1(n_677), .B2(n_681), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_718), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_725), .B(n_676), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_760), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_768), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_745), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_715), .B(n_668), .Y(n_795) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_724), .A2(n_649), .B1(n_656), .B2(n_673), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_706), .B(n_697), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_731), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_731), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_752), .Y(n_800) );
OAI21xp33_ASAP7_75t_L g801 ( .A1(n_738), .A2(n_672), .B(n_649), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_761), .B(n_689), .Y(n_802) );
OAI322xp33_ASAP7_75t_L g803 ( .A1(n_739), .A2(n_741), .A3(n_719), .B1(n_722), .B2(n_757), .C1(n_734), .C2(n_736), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_710), .B(n_688), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_708), .Y(n_805) );
OAI32xp33_ASAP7_75t_L g806 ( .A1(n_702), .A2(n_675), .A3(n_687), .B1(n_684), .B2(n_650), .Y(n_806) );
AOI322xp5_ASAP7_75t_L g807 ( .A1(n_723), .A2(n_687), .A3(n_675), .B1(n_537), .B2(n_417), .C1(n_683), .C2(n_695), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_701), .B(n_537), .Y(n_808) );
OAI21xp5_ASAP7_75t_SL g809 ( .A1(n_780), .A2(n_753), .B(n_760), .Y(n_809) );
OAI21xp33_ASAP7_75t_SL g810 ( .A1(n_780), .A2(n_728), .B(n_703), .Y(n_810) );
AOI21xp33_ASAP7_75t_SL g811 ( .A1(n_794), .A2(n_726), .B(n_750), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g812 ( .A1(n_769), .A2(n_747), .B(n_763), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_769), .A2(n_742), .B1(n_737), .B2(n_713), .Y(n_813) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_806), .A2(n_765), .B(n_754), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_792), .B(n_794), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_781), .B(n_705), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_774), .Y(n_817) );
AOI32xp33_ASAP7_75t_L g818 ( .A1(n_792), .A2(n_712), .A3(n_717), .B1(n_713), .B2(n_756), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_789), .A2(n_717), .B1(n_732), .B2(n_729), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_801), .A2(n_730), .B1(n_746), .B2(n_743), .Y(n_820) );
INVx1_ASAP7_75t_SL g821 ( .A(n_804), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_803), .B(n_751), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_777), .A2(n_709), .B1(n_707), .B2(n_711), .C(n_721), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_777), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_783), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_786), .A2(n_762), .B1(n_748), .B2(n_758), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_796), .A2(n_758), .B(n_752), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g828 ( .A1(n_776), .A2(n_766), .B1(n_767), .B2(n_54), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_807), .B(n_52), .C(n_53), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_796), .A2(n_66), .B(n_67), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_822), .A2(n_782), .B1(n_771), .B2(n_772), .C(n_779), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_817), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_810), .A2(n_772), .B(n_782), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_SL g834 ( .A1(n_809), .A2(n_770), .B(n_802), .C(n_795), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_816), .B(n_805), .Y(n_835) );
AO22x1_ASAP7_75t_L g836 ( .A1(n_824), .A2(n_784), .B1(n_797), .B2(n_791), .Y(n_836) );
AOI211xp5_ASAP7_75t_L g837 ( .A1(n_828), .A2(n_808), .B(n_788), .C(n_799), .Y(n_837) );
AOI211xp5_ASAP7_75t_SL g838 ( .A1(n_830), .A2(n_787), .B(n_785), .C(n_790), .Y(n_838) );
AOI211xp5_ASAP7_75t_L g839 ( .A1(n_811), .A2(n_798), .B(n_800), .C(n_793), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_819), .A2(n_829), .B(n_813), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_823), .B(n_798), .C(n_800), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_832), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_840), .B(n_815), .Y(n_843) );
NAND3xp33_ASAP7_75t_L g844 ( .A(n_837), .B(n_818), .C(n_814), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_833), .A2(n_812), .B(n_827), .Y(n_845) );
NOR3xp33_ASAP7_75t_L g846 ( .A(n_835), .B(n_821), .C(n_820), .Y(n_846) );
NAND4xp25_ASAP7_75t_SL g847 ( .A(n_831), .B(n_826), .C(n_821), .D(n_825), .Y(n_847) );
NAND2x1p5_ASAP7_75t_SL g848 ( .A(n_843), .B(n_834), .Y(n_848) );
NOR3xp33_ASAP7_75t_SL g849 ( .A(n_847), .B(n_841), .C(n_838), .Y(n_849) );
NAND4xp25_ASAP7_75t_L g850 ( .A(n_844), .B(n_839), .C(n_836), .D(n_793), .Y(n_850) );
NOR3x1_ASAP7_75t_L g851 ( .A(n_845), .B(n_778), .C(n_775), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_851), .Y(n_852) );
OAI222xp33_ASAP7_75t_L g853 ( .A1(n_848), .A2(n_842), .B1(n_846), .B2(n_778), .C1(n_775), .C2(n_773), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_849), .B(n_773), .Y(n_854) );
XNOR2x1_ASAP7_75t_L g855 ( .A(n_854), .B(n_850), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_852), .B(n_68), .Y(n_856) );
AOI311xp33_ASAP7_75t_L g857 ( .A1(n_855), .A2(n_853), .A3(n_854), .B(n_72), .C(n_73), .Y(n_857) );
OAI22x1_ASAP7_75t_L g858 ( .A1(n_856), .A2(n_69), .B1(n_71), .B2(n_75), .Y(n_858) );
INVx4_ASAP7_75t_L g859 ( .A(n_857), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_859), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_860), .A2(n_858), .B(n_79), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_861), .A2(n_76), .B(n_82), .Y(n_862) );
OR2x6_ASAP7_75t_L g863 ( .A(n_862), .B(n_83), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_863), .A2(n_84), .B1(n_87), .B2(n_90), .Y(n_864) );
endmodule