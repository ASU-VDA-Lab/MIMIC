module fake_jpeg_12744_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_14),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_2),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_31),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_69),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_58),
.B1(n_74),
.B2(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_23),
.B1(n_16),
.B2(n_20),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_65),
.B1(n_24),
.B2(n_22),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_46),
.Y(n_82)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_23),
.B1(n_19),
.B2(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_20),
.B1(n_26),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_44),
.B1(n_33),
.B2(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_42),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_73),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_26),
.B1(n_19),
.B2(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_80),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_103),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_43),
.B1(n_39),
.B2(n_44),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_17),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_68),
.B1(n_56),
.B2(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_100),
.B1(n_42),
.B2(n_57),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_46),
.B1(n_42),
.B2(n_43),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_105),
.B(n_52),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_99),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_17),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_32),
.C(n_30),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_46),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_30),
.B1(n_34),
.B2(n_33),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_42),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_67),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_24),
.B(n_22),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_84),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_113),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_80),
.B1(n_95),
.B2(n_64),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_52),
.B1(n_44),
.B2(n_49),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_134),
.B1(n_138),
.B2(n_85),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_78),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_127),
.B(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_78),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_59),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_133),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_49),
.B1(n_59),
.B2(n_67),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_29),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_51),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_96),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_64),
.B1(n_51),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_88),
.B1(n_75),
.B2(n_84),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_140),
.A2(n_153),
.B1(n_167),
.B2(n_29),
.Y(n_195)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_149),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_75),
.B(n_98),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_144),
.A2(n_11),
.B(n_15),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_87),
.B(n_85),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_144),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_162),
.B1(n_129),
.B2(n_123),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_105),
.C(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_111),
.C(n_133),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_113),
.A2(n_102),
.B1(n_105),
.B2(n_95),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_81),
.B1(n_109),
.B2(n_101),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_99),
.B(n_109),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_104),
.B(n_77),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_112),
.A2(n_22),
.B(n_33),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_51),
.A3(n_86),
.B1(n_34),
.B2(n_72),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_29),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_86),
.B1(n_34),
.B2(n_72),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_0),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_1),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_127),
.B1(n_118),
.B2(n_138),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_127),
.B1(n_118),
.B2(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_177),
.B(n_179),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_121),
.B1(n_134),
.B2(n_117),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_168),
.B1(n_159),
.B2(n_169),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_111),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_111),
.C(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_111),
.C(n_119),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_164),
.C(n_147),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_119),
.B(n_128),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_201),
.B(n_1),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_128),
.B1(n_86),
.B2(n_72),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_203),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_194),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_198),
.B1(n_167),
.B2(n_142),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_161),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_11),
.B(n_15),
.C(n_14),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_154),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_10),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_172),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_140),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_218),
.C(n_222),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_216),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_219),
.B1(n_221),
.B2(n_225),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_217),
.B(n_194),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_145),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_153),
.B1(n_142),
.B2(n_147),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_142),
.B1(n_165),
.B2(n_154),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_166),
.B1(n_156),
.B2(n_141),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_175),
.B1(n_197),
.B2(n_191),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_148),
.C(n_146),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_226),
.C(n_200),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_25),
.C(n_18),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_174),
.A2(n_25),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_200),
.B(n_186),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_25),
.B1(n_14),
.B2(n_13),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_201),
.B(n_173),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_196),
.A2(n_12),
.B1(n_13),
.B2(n_5),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_245),
.B1(n_248),
.B2(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_202),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_246),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_218),
.B(n_202),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_221),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_251),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_199),
.B1(n_205),
.B2(n_198),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_185),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_176),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_252),
.C(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_199),
.B1(n_187),
.B2(n_186),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_230),
.B1(n_231),
.B2(n_212),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_204),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_211),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_204),
.C(n_12),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_256),
.C(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_12),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_248),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_255),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_226),
.C(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_272),
.C(n_274),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_223),
.C(n_211),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_253),
.C(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_236),
.C(n_241),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_286),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_256),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_249),
.B1(n_245),
.B2(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_290),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_244),
.C(n_223),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_223),
.C(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_4),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_262),
.B1(n_272),
.B2(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_268),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_277),
.B(n_267),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_303),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_277),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_292),
.B1(n_283),
.B2(n_7),
.Y(n_307)
);

AOI211xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_7),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_5),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_6),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_281),
.C(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_6),
.B1(n_7),
.B2(n_293),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_315),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_7),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_299),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_300),
.C(n_305),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_306),
.A2(n_301),
.B(n_310),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_307),
.C(n_312),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_315),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_327),
.A2(n_325),
.B(n_326),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B(n_319),
.C(n_320),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_331),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_324),
.Y(n_333)
);


endmodule