module fake_jpeg_7122_n_100 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_0),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_60),
.C(n_59),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_0),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_55),
.C(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_77),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_53),
.B1(n_48),
.B2(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_74),
.B1(n_45),
.B2(n_5),
.Y(n_84)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_51),
.B1(n_50),
.B2(n_49),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_82),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_44),
.B1(n_43),
.B2(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_6),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_85),
.B1(n_89),
.B2(n_21),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_18),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_27),
.C(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_30),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_31),
.C(n_32),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_33),
.B(n_34),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_38),
.Y(n_100)
);


endmodule