module fake_jpeg_78_n_691 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_553;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g169 ( 
.A(n_61),
.Y(n_169)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_64),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_66),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_68),
.Y(n_190)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_72),
.B(n_74),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_83),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_89),
.B(n_95),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_17),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx2_ASAP7_75t_SL g149 ( 
.A(n_101),
.Y(n_149)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_107),
.B(n_112),
.Y(n_216)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_117),
.B(n_12),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_44),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_130),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_127),
.Y(n_139)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_26),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_43),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_46),
.B1(n_21),
.B2(n_50),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_136),
.A2(n_138),
.B1(n_140),
.B2(n_145),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_46),
.B1(n_21),
.B2(n_50),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_46),
.B1(n_21),
.B2(n_50),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_83),
.A2(n_52),
.B1(n_51),
.B2(n_22),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_142),
.A2(n_171),
.B1(n_214),
.B2(n_221),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_74),
.B1(n_113),
.B2(n_61),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_19),
.B1(n_51),
.B2(n_40),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_151),
.A2(n_187),
.B(n_23),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_63),
.A2(n_52),
.B1(n_51),
.B2(n_40),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_155),
.A2(n_176),
.B1(n_193),
.B2(n_0),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_158),
.B(n_164),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_43),
.C(n_56),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_163),
.B(n_0),
.C(n_1),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_43),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_22),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_167),
.B(n_174),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_84),
.A2(n_22),
.B1(n_52),
.B2(n_40),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_28),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_65),
.A2(n_28),
.B1(n_31),
.B2(n_53),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_66),
.B(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_185),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_67),
.B(n_31),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_86),
.A2(n_31),
.B1(n_55),
.B2(n_53),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_70),
.B(n_56),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_196),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_87),
.A2(n_56),
.B1(n_55),
.B2(n_53),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_71),
.B(n_55),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_88),
.B(n_41),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_204),
.B(n_206),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_76),
.B(n_41),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_97),
.B(n_49),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_34),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_104),
.A2(n_49),
.B1(n_39),
.B2(n_36),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_105),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_217),
.B(n_11),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_111),
.A2(n_49),
.B1(n_39),
.B2(n_36),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_80),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_171),
.B1(n_221),
.B2(n_214),
.Y(n_241)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g307 ( 
.A(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_226),
.Y(n_349)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_227),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_138),
.A2(n_82),
.B1(n_81),
.B2(n_34),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_228),
.A2(n_239),
.B1(n_241),
.B2(n_245),
.Y(n_320)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_229),
.Y(n_328)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_230),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_231),
.B(n_246),
.Y(n_310)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_236),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_142),
.A2(n_33),
.B1(n_23),
.B2(n_26),
.Y(n_239)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_244),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_200),
.A2(n_33),
.B1(n_23),
.B2(n_26),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_169),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_247),
.Y(n_323)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_248),
.B(n_250),
.Y(n_314)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_249),
.Y(n_352)
);

BUFx16f_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_251),
.B(n_252),
.Y(n_353)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_254),
.B(n_256),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_156),
.A2(n_33),
.B1(n_27),
.B2(n_15),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_255),
.A2(n_260),
.B1(n_266),
.B2(n_293),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_258),
.Y(n_361)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_161),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_259),
.B(n_264),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_151),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_133),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_261),
.B(n_275),
.Y(n_341)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_262),
.B(n_265),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_157),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_263),
.A2(n_272),
.B1(n_284),
.B2(n_287),
.Y(n_308)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_162),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_222),
.A2(n_187),
.B1(n_136),
.B2(n_210),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_184),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_267),
.B(n_269),
.Y(n_339)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_270),
.B(n_271),
.Y(n_347)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_216),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_276),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_139),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_183),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_278),
.B(n_281),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_180),
.Y(n_279)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_159),
.Y(n_280)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_132),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_190),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_285),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g351 ( 
.A1(n_283),
.A2(n_194),
.B1(n_186),
.B2(n_220),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_181),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_193),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_137),
.B1(n_150),
.B2(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_143),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_181),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_195),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_146),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_291),
.A2(n_179),
.B1(n_159),
.B2(n_169),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_145),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_208),
.A2(n_219),
.B1(n_210),
.B2(n_140),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_134),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_294),
.B(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_192),
.B(n_10),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_172),
.B(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_297),
.B(n_3),
.Y(n_336)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_175),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_194),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_166),
.A2(n_11),
.B1(n_10),
.B2(n_5),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_186),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_302),
.A2(n_303),
.B1(n_137),
.B2(n_195),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_134),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_304),
.A2(n_313),
.B1(n_317),
.B2(n_333),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_215),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_305),
.B(n_321),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_131),
.B1(n_147),
.B2(n_223),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_315),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_224),
.A2(n_147),
.B1(n_131),
.B2(n_198),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_292),
.A2(n_179),
.B(n_169),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_319),
.A2(n_325),
.B(n_349),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_234),
.B(n_268),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_170),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_329),
.B(n_330),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_231),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_332),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_182),
.B1(n_198),
.B2(n_150),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_240),
.B(n_274),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_334),
.B(n_338),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_336),
.B(n_355),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_228),
.B(n_170),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_266),
.B(n_223),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_340),
.B(n_344),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_244),
.A2(n_212),
.B1(n_207),
.B2(n_201),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_342),
.A2(n_351),
.B(n_280),
.Y(n_370)
);

OR2x2_ASAP7_75t_SL g343 ( 
.A(n_250),
.B(n_135),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_343),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_278),
.B(n_220),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_277),
.A2(n_212),
.B1(n_207),
.B2(n_201),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_359),
.B1(n_226),
.B2(n_237),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_277),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_301),
.B1(n_230),
.B2(n_254),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_277),
.B(n_4),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_239),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_280),
.B(n_4),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_263),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_272),
.B(n_238),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_313),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_368),
.B(n_374),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_370),
.A2(n_413),
.B1(n_335),
.B2(n_306),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_373),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_361),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_250),
.C(n_271),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_379),
.C(n_399),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_276),
.C(n_256),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_376),
.B(n_387),
.C(n_396),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_378),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_264),
.C(n_267),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_299),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_361),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_406),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_340),
.A2(n_251),
.B1(n_229),
.B2(n_300),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_382),
.A2(n_394),
.B1(n_414),
.B2(n_352),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_355),
.A2(n_249),
.B1(n_302),
.B2(n_289),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_320),
.A2(n_326),
.B1(n_323),
.B2(n_338),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_320),
.A2(n_284),
.B1(n_279),
.B2(n_243),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_386),
.A2(n_397),
.B1(n_405),
.B2(n_408),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_303),
.C(n_236),
.Y(n_387)
);

BUFx8_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_393),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_326),
.A2(n_235),
.B1(n_290),
.B2(n_225),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_323),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_395),
.A2(n_400),
.B(n_410),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_363),
.A2(n_8),
.B1(n_9),
.B2(n_329),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_305),
.B(n_8),
.C(n_9),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_365),
.A2(n_8),
.B1(n_345),
.B2(n_310),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_334),
.C(n_311),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_322),
.C(n_337),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_404),
.B(n_353),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_346),
.A2(n_351),
.B1(n_317),
.B2(n_319),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_316),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_412),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_351),
.A2(n_348),
.B1(n_308),
.B2(n_324),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_333),
.A2(n_351),
.B1(n_304),
.B2(n_348),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_409),
.A2(n_361),
.B1(n_306),
.B2(n_357),
.Y(n_447)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_352),
.A2(n_349),
.B1(n_356),
.B2(n_353),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_336),
.B1(n_348),
.B2(n_312),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_312),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_428),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_377),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_424),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_401),
.B(n_314),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_423),
.B(n_452),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_377),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_403),
.A2(n_389),
.B1(n_394),
.B2(n_369),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_426),
.B1(n_442),
.B2(n_409),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_378),
.A2(n_362),
.B1(n_328),
.B2(n_358),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_402),
.Y(n_428)
);

AOI21xp33_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_350),
.B(n_347),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_429),
.A2(n_373),
.B(n_395),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_372),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_435),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_376),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_390),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_339),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_441),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_367),
.B(n_322),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_369),
.A2(n_353),
.B1(n_331),
.B2(n_328),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_356),
.B(n_307),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_444),
.A2(n_451),
.B(n_440),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_447),
.A2(n_418),
.B1(n_433),
.B2(n_382),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_375),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_453),
.C(n_398),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_451),
.A2(n_396),
.B(n_371),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_411),
.B(n_327),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_379),
.B(n_327),
.C(n_335),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_307),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_456),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_436),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_463),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_458),
.A2(n_470),
.B(n_477),
.Y(n_498)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_417),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_462),
.A2(n_447),
.B1(n_419),
.B2(n_422),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_455),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_430),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_465),
.B(n_471),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_467),
.A2(n_426),
.B1(n_442),
.B2(n_386),
.Y(n_518)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_433),
.A2(n_385),
.B1(n_400),
.B2(n_392),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_469),
.A2(n_481),
.B1(n_425),
.B2(n_437),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_444),
.A2(n_388),
.B(n_408),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_430),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_434),
.B(n_412),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_472),
.B(n_479),
.Y(n_515)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_473),
.Y(n_509)
);

AO22x1_ASAP7_75t_L g475 ( 
.A1(n_421),
.A2(n_405),
.B1(n_384),
.B2(n_388),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_SL g513 ( 
.A1(n_475),
.A2(n_481),
.B(n_467),
.C(n_469),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_406),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_397),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_489),
.C(n_449),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_418),
.A2(n_392),
.B1(n_374),
.B2(n_404),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_482),
.Y(n_508)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_454),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_420),
.B(n_399),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g524 ( 
.A(n_487),
.Y(n_524)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_416),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_490),
.Y(n_525)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_491),
.B(n_440),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_424),
.B(n_391),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_492),
.B(n_435),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_444),
.A2(n_388),
.B(n_383),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_493),
.A2(n_415),
.B(n_448),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_428),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_495),
.B(n_522),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_520),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_497),
.B(n_504),
.C(n_519),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_466),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_499),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_438),
.B(n_439),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_501),
.A2(n_502),
.B(n_526),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_477),
.A2(n_415),
.B(n_422),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_432),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_503),
.B(n_505),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_461),
.B(n_443),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_511),
.A2(n_512),
.B1(n_518),
.B2(n_523),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_514),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_466),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_462),
.A2(n_476),
.B1(n_493),
.B2(n_474),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_516),
.A2(n_476),
.B1(n_475),
.B2(n_477),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_417),
.C(n_432),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_468),
.Y(n_521)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_521),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_474),
.B(n_450),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_476),
.A2(n_431),
.B1(n_452),
.B2(n_441),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_486),
.B(n_446),
.Y(n_527)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_527),
.B(n_529),
.C(n_478),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_486),
.B(n_446),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_443),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_484),
.C(n_464),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_459),
.Y(n_533)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_533),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_417),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_534),
.B(n_545),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_536),
.A2(n_506),
.B1(n_518),
.B2(n_523),
.Y(n_568)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_525),
.Y(n_539)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_539),
.Y(n_574)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_525),
.Y(n_540)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_459),
.Y(n_541)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_541),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_524),
.B(n_471),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_542),
.B(n_560),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_511),
.A2(n_465),
.B1(n_478),
.B2(n_463),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_543),
.A2(n_563),
.B1(n_514),
.B2(n_521),
.Y(n_565)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_544),
.Y(n_566)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_550),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_507),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_507),
.B(n_457),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_553),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_519),
.B(n_453),
.C(n_480),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_559),
.C(n_503),
.Y(n_567)
);

BUFx12f_ASAP7_75t_SL g554 ( 
.A(n_498),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_554),
.A2(n_458),
.B(n_513),
.Y(n_588)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_494),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_556),
.B(n_557),
.Y(n_587)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_494),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_558),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_497),
.B(n_453),
.C(n_480),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_515),
.B(n_472),
.Y(n_560)
);

NAND2x1_ASAP7_75t_L g561 ( 
.A(n_498),
.B(n_492),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_561),
.B(n_562),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_499),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_515),
.B(n_487),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_564),
.B(n_491),
.Y(n_578)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_567),
.B(n_588),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_568),
.A2(n_569),
.B1(n_581),
.B2(n_544),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_536),
.A2(n_506),
.B1(n_502),
.B2(n_501),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_562),
.A2(n_516),
.B(n_512),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_570),
.A2(n_532),
.B(n_547),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_537),
.B(n_530),
.C(n_505),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_572),
.B(n_575),
.C(n_577),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_456),
.C(n_508),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_508),
.C(n_490),
.Y(n_577)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_578),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_559),
.B(n_427),
.C(n_488),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_580),
.B(n_583),
.C(n_555),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_550),
.A2(n_513),
.B1(n_475),
.B2(n_528),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_427),
.C(n_485),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_538),
.A2(n_475),
.B1(n_513),
.B2(n_509),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_592),
.B1(n_565),
.B2(n_566),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_555),
.B(n_545),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_590),
.B(n_549),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_543),
.A2(n_546),
.B1(n_532),
.B2(n_551),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_591),
.B(n_582),
.Y(n_594)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_594),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_595),
.B(n_605),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_587),
.B(n_533),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_596),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_548),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g623 ( 
.A(n_599),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_577),
.B(n_582),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_600),
.Y(n_628)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_601),
.Y(n_617)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_602),
.Y(n_629)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_604),
.B(n_616),
.Y(n_634)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_608),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_580),
.B(n_563),
.Y(n_607)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_607),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_549),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_539),
.C(n_540),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_613),
.C(n_614),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_610),
.B(n_611),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_569),
.B(n_561),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_568),
.A2(n_547),
.B1(n_541),
.B2(n_535),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_612),
.A2(n_557),
.B1(n_510),
.B2(n_509),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_561),
.C(n_535),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_585),
.B(n_558),
.C(n_556),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_554),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_615),
.B(n_588),
.C(n_566),
.Y(n_625)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_612),
.A2(n_592),
.B(n_579),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_618),
.A2(n_614),
.B(n_613),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_597),
.A2(n_589),
.B1(n_581),
.B2(n_574),
.Y(n_619)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_619),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_610),
.A2(n_576),
.B1(n_570),
.B2(n_579),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_620),
.B(n_626),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_625),
.B(n_429),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_596),
.A2(n_586),
.B1(n_571),
.B2(n_531),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_611),
.A2(n_571),
.B1(n_531),
.B2(n_513),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_630),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_572),
.C(n_571),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_510),
.Y(n_646)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_637),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_609),
.Y(n_638)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_638),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_626),
.A2(n_598),
.B(n_603),
.Y(n_639)
);

AO21x1_ASAP7_75t_L g661 ( 
.A1(n_639),
.A2(n_641),
.B(n_651),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_631),
.B(n_608),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_640),
.B(n_648),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_627),
.A2(n_603),
.B(n_615),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_624),
.B(n_593),
.C(n_606),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_642),
.B(n_644),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_624),
.B(n_593),
.C(n_578),
.Y(n_644)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_646),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_647),
.B(n_649),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_628),
.B(n_500),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_623),
.B(n_500),
.Y(n_649)
);

AOI211xp5_ASAP7_75t_L g651 ( 
.A1(n_617),
.A2(n_483),
.B(n_473),
.C(n_460),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_633),
.B(n_482),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_652),
.B(n_625),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_633),
.B(n_407),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_653),
.A2(n_620),
.B1(n_629),
.B2(n_619),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_643),
.B(n_630),
.C(n_621),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_656),
.B(n_659),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_657),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_650),
.A2(n_617),
.B1(n_622),
.B2(n_629),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g671 ( 
.A1(n_658),
.A2(n_651),
.B1(n_634),
.B2(n_647),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_637),
.B(n_635),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_663),
.B(n_665),
.Y(n_674)
);

OAI322xp33_ASAP7_75t_L g665 ( 
.A1(n_650),
.A2(n_621),
.A3(n_618),
.B1(n_635),
.B2(n_634),
.C1(n_427),
.C2(n_360),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_662),
.B(n_642),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_667),
.B(n_671),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g668 ( 
.A1(n_654),
.A2(n_644),
.B(n_639),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_668),
.A2(n_669),
.B(n_661),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_655),
.A2(n_641),
.B(n_645),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_664),
.B(n_652),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_672),
.B(n_675),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_660),
.B(n_357),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_678),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_671),
.B(n_654),
.Y(n_678)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_673),
.B(n_656),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_681),
.C(n_670),
.Y(n_682)
);

AOI21xp33_ASAP7_75t_L g681 ( 
.A1(n_674),
.A2(n_666),
.B(n_661),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_682),
.B(n_683),
.C(n_657),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_677),
.B(n_670),
.C(n_663),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_684),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_685),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_686),
.B(n_658),
.Y(n_688)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_688),
.B(n_679),
.C(n_357),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_689),
.A2(n_307),
.B(n_360),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_364),
.B(n_681),
.Y(n_691)
);


endmodule