module real_jpeg_16718_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_536),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_0),
.B(n_537),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_1),
.B(n_61),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_1),
.B(n_290),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_1),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_1),
.B(n_439),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g476 ( 
.A(n_1),
.B(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_1),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_1),
.B(n_509),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

NAND2x1p5_ASAP7_75t_L g35 ( 
.A(n_2),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_2),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_2),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_3),
.Y(n_351)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_3),
.Y(n_443)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g480 ( 
.A(n_4),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_5),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_5),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_5),
.A2(n_11),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_6),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_6),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_6),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_6),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_6),
.B(n_253),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_7),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_7),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_8),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_9),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_9),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_9),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_9),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_9),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_9),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_9),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_10),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_10),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_10),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_10),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_10),
.B(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_10),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_10),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_10),
.B(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_11),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_11),
.B(n_85),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_11),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_11),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_11),
.B(n_495),
.Y(n_494)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_85),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_13),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_13),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_13),
.B(n_297),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

BUFx4f_ASAP7_75t_L g249 ( 
.A(n_15),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_15),
.Y(n_422)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_16),
.Y(n_537)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_17),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_110),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_72),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_72),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_23),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_40),
.CI(n_55),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.C(n_33),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_25),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_25),
.A2(n_26),
.B1(n_63),
.B2(n_64),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_25),
.B(n_162),
.C(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_25),
.A2(n_26),
.B1(n_232),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_63),
.C(n_68),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_30),
.B(n_125),
.C(n_130),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_30),
.B(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx2_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_34),
.B(n_245),
.C(n_255),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_34),
.A2(n_35),
.B1(n_255),
.B2(n_256),
.Y(n_374)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_39),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_79),
.C(n_84),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_41),
.A2(n_53),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_45),
.Y(n_212)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_47),
.B(n_134),
.C(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_47),
.B(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.C(n_62),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_63),
.A2(n_64),
.B1(n_101),
.B2(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_63),
.A2(n_64),
.B1(n_155),
.B2(n_156),
.Y(n_320)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_101),
.C(n_105),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_64),
.B(n_156),
.C(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.C(n_95),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.C(n_90),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_83),
.Y(n_317)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_84),
.B(n_205),
.C(n_208),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_84),
.B(n_208),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_90),
.B(n_204),
.C(n_210),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_90),
.A2(n_91),
.B1(n_210),
.B2(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_168),
.C(n_173),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_91),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_94),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_108),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_97),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_102),
.B1(n_133),
.B2(n_134),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_101),
.A2(n_102),
.B1(n_299),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_133),
.C(n_138),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_102),
.B(n_299),
.C(n_300),
.Y(n_298)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_104),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21x1_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_177),
.B(n_534),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_114),
.B(n_117),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_143),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.C(n_132),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_124),
.B(n_132),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_130),
.A2(n_162),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_133),
.A2(n_134),
.B1(n_170),
.B2(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_134),
.B(n_252),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_SL g410 ( 
.A(n_134),
.B(n_308),
.Y(n_410)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_136),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_137),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_163),
.C(n_167),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_160),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_145),
.B(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_147),
.B(n_160),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.C(n_155),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_159),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_169),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_195),
.C(n_198),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_170),
.A2(n_171),
.B1(n_198),
.B2(n_199),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_170),
.B(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_171),
.B(n_418),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_172),
.Y(n_327)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_258),
.B(n_531),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_216),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_181),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_182),
.B(n_184),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_187),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_203),
.C(n_213),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_191),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_201),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_192),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_194),
.B(n_201),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_196),
.B(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_196),
.B(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_198),
.A2(n_199),
.B1(n_295),
.B2(n_296),
.Y(n_346)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_199),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_213),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_207),
.Y(n_301)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

OR2x2_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_217),
.B(n_219),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.C(n_226),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_220),
.B(n_224),
.Y(n_395)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_226),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_239),
.C(n_243),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_227),
.A2(n_228),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_236),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_229),
.B(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_231),
.B(n_237),
.Y(n_381)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_245),
.A2(n_246),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.C(n_252),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_247),
.A2(n_252),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_252),
.Y(n_308)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2x1_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_525),
.Y(n_258)
);

NAND4xp25_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_382),
.C(n_396),
.D(n_401),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_359),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_335),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_262),
.B(n_335),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_302),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_263),
.B(n_303),
.C(n_318),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_280),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_278),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_277),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_271),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_271),
.A2(n_274),
.B(n_278),
.C(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_273),
.B(n_277),
.Y(n_376)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_276),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_280),
.B(n_363),
.C(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_293),
.C(n_298),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_281),
.B(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_285),
.C(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_293),
.A2(n_294),
.B1(n_298),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_297),
.Y(n_518)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_299),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_300),
.B(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_318),
.Y(n_302)
);

XOR2x2_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_310),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_369),
.C(n_370),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_322),
.B(n_324),
.Y(n_321)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_SL g496 ( 
.A(n_313),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.C(n_328),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_321),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_328),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.C(n_333),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_329),
.B(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_330),
.A2(n_331),
.B1(n_333),
.B2(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.C(n_342),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_336),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_338),
.A2(n_339),
.B1(n_342),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.C(n_347),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_343),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_347),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_352),
.C(n_355),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_348),
.B(n_355),
.Y(n_448)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_352),
.B(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

OAI21x1_ASAP7_75t_SL g526 ( 
.A1(n_359),
.A2(n_527),
.B(n_528),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_360),
.B(n_361),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_366),
.C(n_380),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_379),
.B2(n_380),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_375),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_390),
.C(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

A2O1A1O1Ixp25_ASAP7_75t_L g525 ( 
.A1(n_382),
.A2(n_396),
.B(n_526),
.C(n_529),
.D(n_530),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_394),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_383),
.B(n_394),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.C(n_392),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_384),
.A2(n_385),
.B1(n_392),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_386),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_397),
.B(n_398),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_426),
.B(n_524),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_423),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_403),
.B(n_423),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.C(n_409),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_404),
.A2(n_405),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_407),
.B(n_409),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.C(n_417),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_417),
.B(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_422),
.Y(n_493)
);

AOI21x1_ASAP7_75t_SL g426 ( 
.A1(n_427),
.A2(n_452),
.B(n_523),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_449),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_428),
.B(n_449),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.C(n_447),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_447),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_438),
.C(n_444),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_457),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_444),
.Y(n_457)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_471),
.B(n_522),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_469),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_454),
.B(n_469),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.C(n_467),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_455),
.A2(n_456),
.B1(n_482),
.B2(n_484),
.Y(n_481)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_467),
.B1(n_468),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_464),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_459),
.A2(n_460),
.B1(n_464),
.B2(n_465),
.Y(n_474)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_485),
.B(n_521),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_481),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_473),
.B(n_481),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.C(n_479),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_498),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_476),
.B1(n_479),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_479),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_482),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_486),
.A2(n_500),
.B(n_520),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_497),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_487),
.B(n_497),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_494),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_494),
.Y(n_506)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_507),
.B(n_519),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_506),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_502),
.B(n_506),
.Y(n_519)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_515),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);


endmodule