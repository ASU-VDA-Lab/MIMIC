module fake_jpeg_17985_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_39),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_76),
.Y(n_90)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_44),
.B1(n_46),
.B2(n_55),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_43),
.B1(n_52),
.B2(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_98),
.Y(n_107)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_95),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_54),
.B1(n_48),
.B2(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_103),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_0),
.C(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_100),
.B1(n_87),
.B2(n_92),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_119),
.B1(n_110),
.B2(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_96),
.B1(n_85),
.B2(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_109),
.B1(n_104),
.B2(n_48),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_131),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_118),
.B(n_22),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_133),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_21),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_2),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_130),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_137),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_23),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_20),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_24),
.B(n_37),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_19),
.Y(n_145)
);

NAND4xp25_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_38),
.C(n_16),
.D(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_26),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_14),
.B(n_30),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_13),
.CI(n_28),
.CON(n_149),
.SN(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_32),
.B(n_11),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);


endmodule