module fake_jpeg_31851_n_439 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_439);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_71),
.Y(n_99)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_34),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_19),
.B1(n_21),
.B2(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_87),
.A2(n_104),
.B1(n_107),
.B2(n_42),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_35),
.B1(n_41),
.B2(n_23),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_88),
.B(n_93),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_25),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_106),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_59),
.B1(n_60),
.B2(n_41),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_25),
.B(n_40),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_35),
.B1(n_41),
.B2(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_20),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_20),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_36),
.Y(n_164)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_133),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_58),
.B1(n_51),
.B2(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_149),
.B1(n_162),
.B2(n_79),
.Y(n_182)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_144),
.Y(n_169)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_34),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_147),
.Y(n_193)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_20),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_23),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_157),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_50),
.B1(n_78),
.B2(n_55),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_71),
.B1(n_65),
.B2(n_72),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

CKINVDCx12_ASAP7_75t_R g155 ( 
.A(n_85),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_87),
.A2(n_45),
.B1(n_67),
.B2(n_73),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_35),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_34),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_111),
.B1(n_115),
.B2(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_183),
.B1(n_187),
.B2(n_113),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_65),
.B(n_71),
.C(n_72),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_182),
.B1(n_96),
.B2(n_122),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_40),
.B(n_38),
.C(n_42),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_36),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_117),
.B1(n_115),
.B2(n_112),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_61),
.C(n_90),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_63),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_100),
.B1(n_121),
.B2(n_117),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_142),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_201),
.Y(n_225)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_209),
.B1(n_215),
.B2(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_203),
.B(n_171),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_204),
.Y(n_236)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_169),
.C(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_211),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_146),
.B1(n_143),
.B2(n_98),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_214),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_114),
.B1(n_161),
.B2(n_152),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_114),
.B1(n_161),
.B2(n_148),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_175),
.A2(n_161),
.B1(n_160),
.B2(n_154),
.Y(n_216)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_181),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_170),
.B(n_179),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_194),
.C(n_200),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_172),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_182),
.B1(n_169),
.B2(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_214),
.B1(n_208),
.B2(n_129),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_238),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_192),
.B(n_177),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_193),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_194),
.B(n_203),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_195),
.B(n_192),
.C(n_201),
.D(n_198),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_242),
.B(n_247),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_209),
.B1(n_199),
.B2(n_206),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_243),
.A2(n_219),
.B1(n_240),
.B2(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_172),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_245),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_266),
.C(n_268),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_237),
.B1(n_219),
.B2(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_222),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_205),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_262),
.B1(n_242),
.B2(n_250),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_228),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_248),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_186),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_208),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_227),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_186),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_269),
.B(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_222),
.C(n_225),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_297),
.C(n_254),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_293),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_261),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_166),
.B1(n_176),
.B2(n_190),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_240),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_248),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_286),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_264),
.B1(n_252),
.B2(n_265),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_285),
.B(n_256),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_239),
.B(n_235),
.C(n_232),
.D(n_219),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_239),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_295),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_253),
.B(n_235),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_234),
.C(n_236),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_299),
.A2(n_310),
.B1(n_312),
.B2(n_318),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_245),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_303),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_267),
.B1(n_257),
.B2(n_262),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_304),
.A2(n_320),
.B1(n_284),
.B2(n_276),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_271),
.C(n_279),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_244),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_309),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_285),
.A2(n_252),
.B1(n_243),
.B2(n_249),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_257),
.C(n_251),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_269),
.C(n_280),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_249),
.B1(n_255),
.B2(n_234),
.Y(n_312)
);

AND3x1_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_308),
.C(n_314),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_256),
.B(n_236),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_191),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_315),
.B(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_181),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_165),
.B1(n_185),
.B2(n_191),
.Y(n_318)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_176),
.B1(n_190),
.B2(n_189),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_134),
.B1(n_132),
.B2(n_135),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_217),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_289),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_282),
.B1(n_277),
.B2(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_287),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_329),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_293),
.C(n_298),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_336),
.C(n_337),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_286),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_332),
.B(n_339),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_334),
.A2(n_299),
.B1(n_310),
.B2(n_308),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_274),
.C(n_189),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_178),
.C(n_153),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_102),
.B(n_122),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_196),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_36),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_344),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_217),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_348),
.C(n_330),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_196),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g347 ( 
.A(n_300),
.B(n_39),
.CI(n_38),
.CON(n_347),
.SN(n_347)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_39),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_163),
.C(n_136),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_351),
.A2(n_90),
.B1(n_32),
.B2(n_54),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_304),
.B(n_318),
.Y(n_352)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_346),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g373 ( 
.A(n_353),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_319),
.C(n_321),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_361),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_140),
.B(n_39),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_356),
.A2(n_357),
.B(n_362),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_14),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_358),
.Y(n_379)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_338),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_102),
.Y(n_380)
);

A2O1A1O1Ixp25_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_40),
.B(n_137),
.C(n_16),
.D(n_18),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_353),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_340),
.B1(n_331),
.B2(n_343),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_365),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_336),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_337),
.A2(n_105),
.B1(n_98),
.B2(n_84),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_368),
.A2(n_84),
.B1(n_128),
.B2(n_44),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_342),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_369),
.B(n_329),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_375),
.Y(n_389)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_328),
.C(n_339),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_387),
.C(n_361),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_350),
.A2(n_348),
.B1(n_347),
.B2(n_105),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_383),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_381),
.A2(n_355),
.B1(n_368),
.B2(n_358),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_382),
.A2(n_102),
.B1(n_47),
.B2(n_28),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_351),
.A2(n_128),
.B1(n_32),
.B2(n_54),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_357),
.B(n_16),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_385),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_356),
.A2(n_370),
.B1(n_360),
.B2(n_362),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_75),
.C(n_70),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_367),
.B(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_394),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_363),
.B(n_366),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_372),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_396),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_367),
.B1(n_32),
.B2(n_48),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_68),
.C(n_64),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_373),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_10),
.B(n_17),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_399),
.B(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_398),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_403),
.B(n_410),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_408),
.B1(n_400),
.B2(n_46),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_379),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_404),
.B(n_409),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_372),
.B1(n_382),
.B2(n_381),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_387),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_383),
.B(n_10),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_13),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_397),
.B(n_8),
.Y(n_412)
);

NOR4xp25_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_11),
.C(n_13),
.D(n_12),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_416),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_391),
.B(n_395),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_415),
.A2(n_0),
.B(n_1),
.Y(n_424)
);

AOI322xp5_ASAP7_75t_L g417 ( 
.A1(n_402),
.A2(n_47),
.A3(n_21),
.B1(n_13),
.B2(n_11),
.C1(n_8),
.C2(n_28),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_418),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_8),
.C(n_21),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_419),
.A2(n_421),
.B(n_409),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_0),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_1),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_428),
.Y(n_430)
);

AOI322xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_425),
.A3(n_429),
.B1(n_417),
.B2(n_418),
.C1(n_21),
.C2(n_5),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_422),
.A2(n_1),
.B(n_2),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_432),
.C(n_433),
.Y(n_434)
);

AOI322xp5_ASAP7_75t_L g432 ( 
.A1(n_427),
.A2(n_21),
.A3(n_28),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_7),
.Y(n_432)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_21),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_433)
);

AOI321xp33_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_21),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_435),
.B(n_2),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_436),
.B(n_434),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_3),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_6),
.B(n_7),
.Y(n_439)
);


endmodule