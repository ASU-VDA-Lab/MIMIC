module fake_jpeg_5499_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_16),
.B1(n_27),
.B2(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_54),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_26),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_75),
.B1(n_89),
.B2(n_99),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_34),
.C(n_33),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_18),
.Y(n_116)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_25),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_25),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_76),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_32),
.B(n_28),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_80),
.Y(n_126)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_34),
.B1(n_33),
.B2(n_16),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_22),
.B1(n_19),
.B2(n_31),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_88),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_16),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_40),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_97),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_17),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_17),
.B1(n_31),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_66),
.B1(n_86),
.B2(n_53),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_21),
.B1(n_27),
.B2(n_24),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_54),
.B1(n_83),
.B2(n_79),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_21),
.B1(n_27),
.B2(n_19),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_122),
.B1(n_130),
.B2(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_89),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_17),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_125),
.B(n_106),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_69),
.B(n_62),
.C(n_57),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_135),
.B1(n_138),
.B2(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_70),
.B1(n_66),
.B2(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_146),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_140),
.B1(n_143),
.B2(n_107),
.Y(n_183)
);

OAI22x1_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_86),
.B1(n_91),
.B2(n_81),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_147),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_65),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_151),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_62),
.B1(n_100),
.B2(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_17),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_154),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_129),
.B(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_84),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_10),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_85),
.C(n_87),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.C(n_128),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_101),
.A3(n_126),
.B1(n_109),
.B2(n_127),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_101),
.B(n_85),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_128),
.B1(n_107),
.B2(n_102),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_57),
.B1(n_61),
.B2(n_87),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_165),
.B1(n_111),
.B2(n_103),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_101),
.A2(n_31),
.B1(n_61),
.B2(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_0),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_116),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_154),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_178),
.Y(n_202)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_181),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_200),
.B1(n_194),
.B2(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_103),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_116),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_31),
.B1(n_117),
.B2(n_118),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_163),
.B1(n_160),
.B2(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_0),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_195),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_0),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_138),
.A2(n_117),
.B1(n_115),
.B2(n_10),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_166),
.B(n_136),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_117),
.C(n_115),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_144),
.C(n_132),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_12),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_204),
.C(n_215),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_157),
.C(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_225),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_211),
.B(n_193),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_142),
.B(n_147),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_214),
.B1(n_221),
.B2(n_187),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_152),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_218),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_179),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_137),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_188),
.A2(n_165),
.B1(n_152),
.B2(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_233),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_231),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_167),
.B1(n_173),
.B2(n_168),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_232),
.A2(n_242),
.B1(n_201),
.B2(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_171),
.B1(n_167),
.B2(n_184),
.C(n_189),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_241),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_239),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_198),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_211),
.B1(n_221),
.B2(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_178),
.C(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_195),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_202),
.B(n_170),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_197),
.C(n_204),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_208),
.B1(n_209),
.B2(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_246),
.C(n_247),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_241),
.B(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_229),
.A2(n_223),
.B1(n_210),
.B2(n_217),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_274),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_229),
.B1(n_227),
.B2(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_248),
.C(n_238),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_232),
.B(n_239),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_246),
.C(n_238),
.Y(n_274)
);

NAND4xp25_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_176),
.C(n_207),
.D(n_225),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_252),
.C(n_248),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_249),
.B1(n_257),
.B2(n_251),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_277),
.A2(n_284),
.B(n_285),
.C(n_261),
.Y(n_292)
);

NAND4xp25_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_250),
.C(n_262),
.D(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_287),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_227),
.B1(n_254),
.B2(n_230),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_272),
.B(n_273),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_291),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_210),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_185),
.B(n_237),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_276),
.C(n_274),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_278),
.B1(n_264),
.B2(n_287),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_271),
.B(n_214),
.C(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_268),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_296),
.B(n_228),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_254),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.C(n_301),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_180),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_295),
.B(n_279),
.C(n_228),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_180),
.A3(n_168),
.B1(n_175),
.B2(n_279),
.C1(n_267),
.C2(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_175),
.C(n_9),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_304),
.Y(n_309)
);


endmodule