module fake_jpeg_2951_n_211 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_211);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_82),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_58),
.B1(n_74),
.B2(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_52),
.B1(n_55),
.B2(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_88),
.B1(n_55),
.B2(n_61),
.Y(n_101)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_103),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_57),
.B(n_63),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_112),
.C(n_80),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_73),
.B(n_64),
.C(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_59),
.B1(n_27),
.B2(n_28),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_114),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_82),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_82),
.B(n_76),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_30),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_130),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_74),
.B1(n_77),
.B2(n_94),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_135),
.B1(n_48),
.B2(n_29),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_70),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.C(n_5),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_70),
.C(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_4),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_72),
.B1(n_69),
.B2(n_82),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_113),
.B(n_96),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_59),
.B(n_24),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_133),
.B(n_104),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_22),
.B1(n_47),
.B2(n_46),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_5),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_141),
.Y(n_164)
);

AOI21x1_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_13),
.B(n_14),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_151),
.C(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_149),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_162)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_156),
.C(n_157),
.Y(n_167)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g166 ( 
.A(n_147),
.Y(n_166)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_21),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_116),
.B(n_133),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_31),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_6),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_15),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_149),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_37),
.C(n_45),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_167),
.C(n_153),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_173),
.B(n_151),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_13),
.B(n_15),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_181),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_172),
.B(n_157),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_187),
.C(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_188),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_151),
.B(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_148),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_175),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_192),
.C(n_193),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_169),
.C(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_163),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_177),
.B(n_163),
.Y(n_199)
);

AOI31xp67_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_171),
.A3(n_166),
.B(n_162),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_201),
.B1(n_16),
.B2(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_190),
.C(n_32),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.C(n_198),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_202),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_35),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_39),
.B(n_40),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_42),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_43),
.Y(n_211)
);


endmodule