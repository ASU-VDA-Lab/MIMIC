module fake_jpeg_16273_n_90 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx13_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_2),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_1),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_51),
.B1(n_5),
.B2(n_6),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_35),
.B1(n_38),
.B2(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_54),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_2),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_3),
.B(n_4),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_65),
.B(n_19),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_63),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_68),
.B1(n_52),
.B2(n_15),
.Y(n_70)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_12),
.B1(n_16),
.B2(n_18),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.C(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_77),
.B1(n_65),
.B2(n_24),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_22),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_83),
.B1(n_80),
.B2(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_74),
.C(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_23),
.B(n_25),
.Y(n_88)
);

OAI211xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_61),
.Y(n_90)
);


endmodule