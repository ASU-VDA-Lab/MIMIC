module real_jpeg_2515_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_244;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_1),
.A2(n_57),
.B1(n_71),
.B2(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_57),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_57),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_2),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_71),
.B(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_61),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_2),
.A2(n_59),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_29),
.C(n_48),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_171),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_2),
.B(n_31),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_53),
.Y(n_226)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_71),
.B1(n_72),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_4),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_145),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_145),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_145),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_45),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_5),
.A2(n_45),
.B1(n_71),
.B2(n_72),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_7),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_277)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_9),
.A2(n_71),
.B1(n_72),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_80),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_80),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_10),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_13),
.A2(n_71),
.B1(n_72),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_13),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_82),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_82),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_82),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_14),
.A2(n_71),
.B1(n_72),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_14),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_125),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_125),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_14),
.A2(n_29),
.B1(n_35),
.B2(n_125),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_16),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_261),
.B1(n_283),
.B2(n_284),
.Y(n_19)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_127),
.B(n_260),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_109),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_22),
.B(n_109),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_23),
.B(n_93),
.C(n_108),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_54),
.C(n_67),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_24),
.A2(n_25),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_28),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_28),
.A2(n_31),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_31),
.B1(n_138),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_28),
.A2(n_31),
.B1(n_175),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_28),
.A2(n_31),
.B1(n_171),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_28),
.A2(n_31),
.B1(n_224),
.B2(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_29),
.B(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_30),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_30),
.A2(n_34),
.B1(n_97),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_30),
.A2(n_97),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_30),
.A2(n_97),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_42),
.A2(n_50),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AO22x2_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_44),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_43),
.B(n_63),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_44),
.A2(n_59),
.A3(n_62),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_44),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_53),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_46),
.A2(n_53),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_46),
.A2(n_53),
.B1(n_167),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_46),
.A2(n_53),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_46),
.A2(n_53),
.B1(n_194),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_46),
.A2(n_53),
.B(n_91),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_50),
.A2(n_118),
.B1(n_166),
.B2(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_61),
.B1(n_87),
.B2(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_59),
.B1(n_74),
.B2(n_76),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_58),
.B(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_58),
.B(n_171),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_72),
.A3(n_76),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_66),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_60),
.A2(n_66),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_60),
.A2(n_66),
.B1(n_141),
.B2(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_60),
.A2(n_66),
.B1(n_156),
.B2(n_203),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_61),
.A2(n_87),
.B1(n_88),
.B2(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_77),
.B1(n_81),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_68),
.A2(n_77),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_68),
.A2(n_77),
.B1(n_144),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_68),
.A2(n_77),
.B1(n_106),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_79),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_108),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_92),
.A2(n_267),
.B1(n_279),
.B2(n_280),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_92),
.Y(n_279)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_103),
.A2(n_105),
.B(n_107),
.Y(n_265)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_114),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.C(n_123),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_116),
.B(n_119),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_150),
.B(n_259),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_148),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_129),
.B(n_148),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_147),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_130),
.B(n_147),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_132),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.C(n_143),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_133),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_137),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_140),
.B(n_143),
.Y(n_250)
);

AOI31xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_244),
.A3(n_253),
.B(n_256),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_189),
.B(n_243),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_177),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_153),
.B(n_177),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.C(n_168),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_154),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_159),
.C(n_163),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_164),
.B(n_168),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_177),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_254),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.CI(n_180),
.CON(n_177),
.SN(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_181),
.B(n_184),
.C(n_188),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_238),
.B(n_242),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_207),
.B(n_237),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_196),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_202),
.C(n_205),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_218),
.B(n_236),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_230),
.B(n_235),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_225),
.B(n_229),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.C(n_252),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_282),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_281),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_278),
.Y(n_272)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);


endmodule