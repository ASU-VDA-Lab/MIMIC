module fake_netlist_6_1276_n_1733 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1733);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1733;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_20),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g154 ( 
.A(n_45),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_54),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_79),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_45),
.Y(n_164)
);

BUFx8_ASAP7_75t_SL g165 ( 
.A(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_81),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_26),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_34),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_53),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_82),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_27),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_90),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_44),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_41),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_25),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_101),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_83),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_22),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_149),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_96),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_5),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_103),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_57),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_110),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_92),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_99),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_18),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_69),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_18),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_42),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_105),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_93),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_41),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_49),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_44),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_84),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_32),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_10),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_107),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_51),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_50),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_61),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_7),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_108),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_9),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_97),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_59),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_42),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_31),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_78),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_94),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_9),
.Y(n_258)
);

INVx4_ASAP7_75t_R g259 ( 
.A(n_63),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_71),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_60),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_77),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_38),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_118),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_74),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_33),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_26),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_111),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_13),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_40),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_114),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_80),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_65),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_134),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_15),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_43),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_116),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_137),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_23),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_48),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_148),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_12),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_151),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_30),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_39),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_147),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_112),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_117),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_48),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_100),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_121),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_88),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_139),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_165),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_157),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_181),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_162),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_217),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_189),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_167),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_167),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_189),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_208),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_167),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_167),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_277),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_164),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_197),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_183),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_164),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_220),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_228),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_202),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_203),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_217),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_231),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_160),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_231),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_283),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_161),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_166),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_190),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_195),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_219),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_235),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_238),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_243),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_208),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_282),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_247),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_211),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_250),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_205),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_227),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_280),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_207),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_226),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_214),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_226),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_215),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_277),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_304),
.A2(n_274),
.B1(n_253),
.B2(n_258),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_364),
.B(n_267),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_303),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_179),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_316),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_248),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_313),
.A2(n_274),
.B1(n_253),
.B2(n_258),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_306),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_309),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_307),
.B(n_248),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_310),
.Y(n_404)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_302),
.B(n_156),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_307),
.B(n_172),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_311),
.B(n_172),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_159),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_333),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_330),
.A2(n_267),
.B1(n_292),
.B2(n_282),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_302),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_175),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_314),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_367),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_314),
.B(n_175),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_185),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_336),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g422 ( 
.A(n_337),
.B(n_286),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_155),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_342),
.A2(n_293),
.B1(n_290),
.B2(n_286),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_344),
.B(n_284),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_338),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_346),
.B(n_284),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_343),
.B(n_185),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_366),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_326),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_372),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_326),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_327),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_320),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_327),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_328),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_328),
.A2(n_163),
.B(n_158),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_380),
.B(n_349),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_387),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_390),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_430),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_374),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_442),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_406),
.B(n_178),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_389),
.B(n_308),
.Y(n_462)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_360),
.C(n_355),
.Y(n_463)
);

NOR2x1p5_ASAP7_75t_L g464 ( 
.A(n_402),
.B(n_289),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_321),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_430),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_381),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_398),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_428),
.A2(n_255),
.B1(n_252),
.B2(n_270),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_398),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_425),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_404),
.B(n_185),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_406),
.B(n_407),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

AND3x2_ASAP7_75t_L g494 ( 
.A(n_418),
.B(n_362),
.C(n_169),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_395),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_380),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_407),
.B(n_176),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_410),
.B(n_359),
.Y(n_501)
);

NOR2x1p5_ASAP7_75t_L g502 ( 
.A(n_421),
.B(n_289),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_391),
.B(n_346),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_432),
.B(n_288),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_436),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_391),
.B(n_331),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_391),
.B(n_331),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_438),
.B(n_361),
.Y(n_511)
);

BUFx4f_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_415),
.B(n_237),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_380),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_435),
.B(n_288),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_416),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_411),
.A2(n_245),
.B1(n_269),
.B2(n_273),
.Y(n_519)
);

BUFx6f_ASAP7_75t_SL g520 ( 
.A(n_427),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_392),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

AO21x1_ASAP7_75t_L g524 ( 
.A1(n_415),
.A2(n_173),
.B(n_168),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_419),
.B(n_216),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_422),
.B(n_419),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_386),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_378),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_378),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_431),
.B(n_182),
.C(n_153),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_409),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_386),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_444),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_380),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_444),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_379),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_379),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_403),
.B(n_218),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_444),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_418),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_409),
.B(n_154),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_428),
.B(n_291),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_383),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g549 ( 
.A1(n_403),
.A2(n_177),
.B(n_174),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_403),
.B(n_223),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_420),
.B(n_291),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_383),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_403),
.B(n_224),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_386),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_411),
.A2(n_412),
.B1(n_423),
.B2(n_434),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_445),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_445),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_382),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_393),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_393),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_434),
.B(n_221),
.C(n_184),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_420),
.B(n_296),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_423),
.B(n_376),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_396),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_396),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_409),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_400),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_400),
.B(n_225),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_382),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_427),
.B(n_296),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_386),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_427),
.B(n_229),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_399),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_399),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_399),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_405),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_409),
.A2(n_212),
.B1(n_234),
.B2(n_236),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_427),
.B(n_297),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_399),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_414),
.B(n_349),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_399),
.Y(n_585)
);

INVx4_ASAP7_75t_SL g586 ( 
.A(n_399),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_440),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_414),
.B(n_209),
.C(n_233),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_429),
.A2(n_206),
.B1(n_204),
.B2(n_201),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_414),
.B(n_232),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_424),
.B(n_244),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_429),
.A2(n_239),
.B1(n_222),
.B2(n_210),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_440),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_440),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_492),
.B(n_249),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_476),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_526),
.B(n_500),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_514),
.B(n_440),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_563),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_563),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_564),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g603 ( 
.A(n_567),
.B(n_433),
.C(n_443),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_564),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_573),
.A2(n_377),
.B1(n_279),
.B2(n_227),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_512),
.B(n_249),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_568),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_525),
.A2(n_241),
.B1(n_301),
.B2(n_300),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_458),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

AND2x6_ASAP7_75t_SL g614 ( 
.A(n_511),
.B(n_501),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_460),
.B(n_446),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_460),
.B(n_446),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_476),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_455),
.B(n_446),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_478),
.B(n_433),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_449),
.B(n_446),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_509),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_478),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_509),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_449),
.B(n_405),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_450),
.B(n_580),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_450),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_405),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_545),
.B(n_443),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_528),
.B(n_405),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_584),
.A2(n_199),
.B1(n_188),
.B2(n_193),
.Y(n_632)
);

O2A1O1Ixp5_ASAP7_75t_L g633 ( 
.A1(n_512),
.A2(n_299),
.B(n_213),
.C(n_256),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_479),
.Y(n_634)
);

INVx8_ASAP7_75t_L g635 ( 
.A(n_546),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_528),
.B(n_529),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_479),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_458),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_512),
.B(n_249),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_529),
.B(n_405),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_480),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_533),
.B(n_249),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_515),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_559),
.B(n_547),
.C(n_463),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

OR2x2_ASAP7_75t_SL g646 ( 
.A(n_530),
.B(n_194),
.Y(n_646)
);

NAND2x1_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_259),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_480),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_447),
.Y(n_649)
);

BUFx5_ASAP7_75t_L g650 ( 
.A(n_451),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_485),
.B(n_439),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_487),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_487),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_550),
.B(n_439),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_581),
.B(n_297),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_533),
.B(n_249),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_540),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_L g658 ( 
.A(n_448),
.B(n_506),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_540),
.B(n_424),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_541),
.B(n_426),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_520),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_447),
.B(n_261),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_447),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_541),
.B(n_426),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_548),
.B(n_275),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_548),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_553),
.B(n_294),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_553),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_533),
.B(n_254),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_569),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_571),
.B(n_437),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_484),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_571),
.B(n_437),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_590),
.B(n_437),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_503),
.B(n_591),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_448),
.B(n_227),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_587),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_588),
.B(n_186),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_503),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_481),
.B(n_350),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_441),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_587),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_584),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_593),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_542),
.B(n_441),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_593),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_519),
.A2(n_356),
.B(n_371),
.C(n_370),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_594),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_565),
.B(n_191),
.C(n_198),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_551),
.B(n_441),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_584),
.B(n_552),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_584),
.Y(n_694)
);

NOR3xp33_ASAP7_75t_L g695 ( 
.A(n_517),
.B(n_371),
.C(n_370),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_519),
.A2(n_369),
.B(n_368),
.C(n_365),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_524),
.A2(n_254),
.B1(n_170),
.B2(n_285),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_594),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_451),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_574),
.A2(n_369),
.B(n_368),
.C(n_365),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_554),
.B(n_246),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_457),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_452),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g704 ( 
.A(n_506),
.B(n_279),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_489),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_524),
.B(n_254),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_562),
.A2(n_254),
.B1(n_170),
.B2(n_285),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_454),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_452),
.Y(n_709)
);

INVx8_ASAP7_75t_L g710 ( 
.A(n_546),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_457),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_576),
.B(n_257),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_489),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_491),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_459),
.B(n_350),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_520),
.A2(n_265),
.B1(n_278),
.B2(n_260),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_484),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_566),
.B(n_464),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_490),
.B(n_262),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_484),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_490),
.B(n_263),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_469),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_491),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_493),
.B(n_454),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_495),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_546),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_462),
.B(n_187),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_493),
.B(n_268),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_484),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_493),
.B(n_272),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_454),
.B(n_276),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_470),
.B(n_254),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_504),
.B(n_200),
.Y(n_733)
);

BUFx8_ASAP7_75t_L g734 ( 
.A(n_520),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_494),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_465),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_470),
.B(n_170),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_470),
.B(n_170),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_531),
.B(n_170),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_531),
.A2(n_170),
.B1(n_285),
.B2(n_357),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_484),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_488),
.B(n_271),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_570),
.B(n_363),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_570),
.B(n_285),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_521),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_582),
.A2(n_295),
.B1(n_358),
.B2(n_357),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_464),
.B(n_279),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_589),
.B(n_363),
.C(n_358),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_523),
.B(n_285),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_469),
.B(n_285),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_592),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_523),
.B(n_285),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_471),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_471),
.B(n_356),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_495),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_472),
.B(n_295),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_498),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_472),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_562),
.A2(n_354),
.B1(n_353),
.B2(n_352),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_473),
.A2(n_354),
.B1(n_353),
.B2(n_352),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_473),
.B(n_351),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_477),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_477),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_612),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

BUFx4f_ASAP7_75t_L g766 ( 
.A(n_638),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_707),
.A2(n_521),
.B1(n_468),
.B2(n_505),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_679),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_639),
.B(n_486),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_649),
.B(n_453),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_628),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_630),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_598),
.B(n_482),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_677),
.B(n_482),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_651),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_686),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_703),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_502),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_715),
.B(n_468),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_654),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_615),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_R g785 ( 
.A(n_709),
.B(n_549),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_657),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_596),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_649),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_618),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_649),
.Y(n_790)
);

NOR2x1_ASAP7_75t_L g791 ( 
.A(n_658),
.B(n_496),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_667),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_649),
.B(n_643),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_672),
.B(n_483),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_669),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_685),
.B(n_575),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_674),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_639),
.B(n_486),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_751),
.B(n_483),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_599),
.B(n_497),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_682),
.B(n_332),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_669),
.Y(n_802)
);

AND2x4_ASAP7_75t_SL g803 ( 
.A(n_726),
.B(n_486),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_671),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_623),
.Y(n_805)
);

INVxp33_ASAP7_75t_L g806 ( 
.A(n_620),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_650),
.B(n_486),
.Y(n_807)
);

HAxp5_ASAP7_75t_L g808 ( 
.A(n_608),
.B(n_0),
.CON(n_808),
.SN(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_709),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_707),
.A2(n_522),
.B1(n_513),
.B2(n_497),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_697),
.A2(n_505),
.B1(n_522),
.B2(n_513),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_674),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_636),
.B(n_498),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_650),
.B(n_486),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_671),
.B(n_507),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_745),
.B(n_332),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_681),
.B(n_507),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_600),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_655),
.A2(n_518),
.B(n_516),
.C(n_508),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_635),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_674),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_622),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_676),
.B(n_508),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_624),
.B(n_516),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_600),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_496),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_745),
.Y(n_827)
);

INVx6_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_697),
.A2(n_475),
.B1(n_466),
.B2(n_465),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_644),
.A2(n_537),
.B1(n_544),
.B2(n_532),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_601),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_706),
.A2(n_475),
.B1(n_466),
.B2(n_558),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_614),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_655),
.B(n_532),
.Y(n_834)
);

NOR2x2_ASAP7_75t_L g835 ( 
.A(n_704),
.B(n_575),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_662),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_706),
.A2(n_539),
.B1(n_544),
.B2(n_543),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_662),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_693),
.B(n_453),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_733),
.B(n_549),
.C(n_339),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_694),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_602),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_643),
.Y(n_843)
);

AND3x1_ASAP7_75t_L g844 ( 
.A(n_678),
.B(n_335),
.C(n_339),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_595),
.A2(n_539),
.B(n_536),
.C(n_537),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_L g846 ( 
.A1(n_733),
.A2(n_335),
.B(n_340),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_626),
.A2(n_543),
.B1(n_557),
.B2(n_558),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_664),
.B(n_577),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_661),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_662),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_650),
.B(n_456),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_607),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_683),
.B(n_496),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_603),
.B(n_340),
.C(n_555),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_661),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_609),
.A2(n_555),
.B1(n_557),
.B2(n_560),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_L g857 ( 
.A(n_635),
.B(n_456),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_747),
.B(n_560),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_710),
.B(n_561),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_742),
.B(n_453),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_643),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_610),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_718),
.A2(n_536),
.B1(n_561),
.B2(n_535),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_659),
.B(n_535),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_735),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_613),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_734),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_613),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_734),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_734),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_691),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_650),
.B(n_456),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_660),
.B(n_535),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_727),
.B(n_577),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_634),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_597),
.B(n_585),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_604),
.B(n_585),
.Y(n_877)
);

AND2x6_ASAP7_75t_L g878 ( 
.A(n_629),
.B(n_583),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_684),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_634),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_665),
.B(n_534),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_687),
.B(n_534),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_666),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_688),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_609),
.A2(n_467),
.B(n_456),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_692),
.B(n_534),
.Y(n_886)
);

AO21x2_ASAP7_75t_L g887 ( 
.A1(n_619),
.A2(n_617),
.B(n_616),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_690),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_710),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_698),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_643),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_712),
.B(n_456),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_637),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_650),
.B(n_461),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_650),
.B(n_461),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_699),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_674),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_637),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_641),
.Y(n_899)
);

INVx3_ASAP7_75t_SL g900 ( 
.A(n_646),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_756),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_645),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_461),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_605),
.B(n_461),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_742),
.B(n_727),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_650),
.B(n_461),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_606),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_645),
.B(n_583),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_625),
.A2(n_467),
.B(n_578),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_645),
.B(n_579),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_702),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_680),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_680),
.B(n_467),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_748),
.B(n_579),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_627),
.B(n_578),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_711),
.Y(n_918)
);

AO21x2_ASAP7_75t_L g919 ( 
.A1(n_595),
.A2(n_586),
.B(n_578),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_556),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_722),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_717),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_763),
.B(n_556),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_717),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_641),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_753),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_762),
.B(n_556),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_627),
.B(n_556),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_631),
.A2(n_474),
.B(n_556),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_716),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_758),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_695),
.B(n_586),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_720),
.B(n_474),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_640),
.A2(n_474),
.B(n_527),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_668),
.B(n_586),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_689),
.B(n_586),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_717),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_705),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_717),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_713),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_611),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_713),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_741),
.B(n_474),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_729),
.B(n_474),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_788),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_906),
.A2(n_696),
.B(n_632),
.C(n_746),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_765),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_906),
.B(n_696),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_914),
.A2(n_621),
.B(n_656),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_773),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_827),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_929),
.A2(n_724),
.B(n_708),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_914),
.A2(n_642),
.B(n_656),
.Y(n_953)
);

OA22x2_ASAP7_75t_L g954 ( 
.A1(n_774),
.A2(n_740),
.B1(n_744),
.B2(n_739),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_788),
.B(n_720),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_781),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_892),
.A2(n_904),
.B(n_887),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_SL g958 ( 
.A1(n_771),
.A2(n_642),
.B(n_670),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_792),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_902),
.A2(n_700),
.B(n_754),
.C(n_761),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_887),
.A2(n_670),
.B(n_647),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_776),
.A2(n_720),
.B(n_731),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_939),
.A2(n_729),
.B(n_728),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_902),
.B(n_673),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_SL g965 ( 
.A1(n_771),
.A2(n_744),
.B(n_739),
.C(n_752),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_939),
.A2(n_821),
.B(n_797),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_764),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_816),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_920),
.A2(n_730),
.B(n_721),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_784),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_809),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_SL g972 ( 
.A1(n_795),
.A2(n_749),
.B(n_804),
.C(n_802),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_774),
.B(n_777),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_799),
.A2(n_633),
.B(n_675),
.C(n_737),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_807),
.A2(n_732),
.B(n_719),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_777),
.B(n_759),
.Y(n_976)
);

CKINVDCx14_ASAP7_75t_R g977 ( 
.A(n_828),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_779),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_798),
.A2(n_738),
.B(n_750),
.C(n_708),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_786),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_920),
.A2(n_729),
.B(n_708),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_782),
.B(n_725),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_775),
.A2(n_729),
.B(n_757),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_834),
.A2(n_736),
.B1(n_757),
.B2(n_755),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_714),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_860),
.A2(n_714),
.B(n_755),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_896),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_768),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_788),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_883),
.B(n_725),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_912),
.Y(n_991)
);

CKINVDCx8_ASAP7_75t_R g992 ( 
.A(n_833),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_788),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_860),
.A2(n_723),
.B(n_652),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_889),
.B(n_723),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_806),
.B(n_736),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_822),
.B(n_653),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_789),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_SL g999 ( 
.A1(n_840),
.A2(n_653),
.B(n_652),
.C(n_648),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_918),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_839),
.A2(n_760),
.B(n_474),
.C(n_527),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_798),
.A2(n_819),
.B(n_845),
.C(n_935),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_834),
.A2(n_760),
.B1(n_527),
.B2(n_62),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_806),
.B(n_527),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_783),
.B(n_6),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_828),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_797),
.A2(n_527),
.B(n_58),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_822),
.B(n_858),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_819),
.A2(n_72),
.B(n_146),
.C(n_145),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_930),
.B(n_138),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_797),
.A2(n_527),
.B(n_136),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_766),
.B(n_133),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_789),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_921),
.B(n_6),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_926),
.B(n_10),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_839),
.A2(n_128),
.B1(n_125),
.B2(n_124),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_767),
.A2(n_122),
.B1(n_109),
.B2(n_106),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_871),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_766),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_767),
.B(n_11),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_812),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_16),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_808),
.B(n_19),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_931),
.B(n_19),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_874),
.B(n_20),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_910),
.A2(n_87),
.B(n_102),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_823),
.A2(n_98),
.B(n_89),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_853),
.A2(n_76),
.B(n_73),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_769),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_801),
.B(n_817),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_800),
.A2(n_52),
.B(n_104),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_882),
.A2(n_21),
.B(n_24),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_886),
.A2(n_21),
.B(n_24),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_850),
.B(n_25),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_867),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_L g1036 ( 
.A(n_865),
.B(n_28),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_889),
.B(n_29),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_813),
.A2(n_32),
.B(n_35),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_808),
.B(n_35),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_941),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_812),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_770),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_828),
.Y(n_1043)
);

BUFx2_ASAP7_75t_SL g1044 ( 
.A(n_901),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_778),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_900),
.B(n_39),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_869),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_835),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_915),
.A2(n_43),
.B(n_46),
.C(n_47),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_836),
.A2(n_838),
.B1(n_863),
.B2(n_790),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_790),
.A2(n_793),
.B1(n_797),
.B2(n_924),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_807),
.A2(n_814),
.B(n_851),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_870),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_908),
.B(n_824),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_SL g1055 ( 
.A(n_846),
.B(n_854),
.C(n_879),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_841),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_841),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_787),
.B(n_805),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_844),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_901),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_917),
.B(n_796),
.Y(n_1061)
);

CKINVDCx8_ASAP7_75t_R g1062 ( 
.A(n_780),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_849),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_L g1064 ( 
.A(n_820),
.B(n_812),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_821),
.B(n_924),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_936),
.A2(n_917),
.B1(n_796),
.B2(n_830),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_821),
.B(n_924),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_814),
.A2(n_907),
.B(n_895),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_884),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_852),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_812),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_840),
.A2(n_888),
.B(n_890),
.C(n_826),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_875),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_872),
.A2(n_894),
.B(n_909),
.C(n_911),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_780),
.B(n_859),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_903),
.B(n_843),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_872),
.A2(n_894),
.B(n_873),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_803),
.B(n_848),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_862),
.B(n_868),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_897),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_SL g1081 ( 
.A1(n_855),
.A2(n_859),
.B1(n_793),
.B2(n_932),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_987),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_991),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_948),
.A2(n_949),
.B(n_958),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_952),
.A2(n_845),
.B(n_885),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1000),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_SL g1087 ( 
.A1(n_1031),
.A2(n_1027),
.B(n_1028),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_981),
.A2(n_856),
.B(n_934),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_964),
.B(n_794),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_988),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_957),
.A2(n_1066),
.A3(n_953),
.B(n_974),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_949),
.A2(n_881),
.B(n_864),
.Y(n_1092)
);

AO32x2_ASAP7_75t_L g1093 ( 
.A1(n_1081),
.A2(n_785),
.A3(n_878),
.B1(n_811),
.B2(n_810),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_946),
.B(n_791),
.C(n_857),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_989),
.B(n_937),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1003),
.A2(n_936),
.B(n_932),
.C(n_848),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1030),
.B(n_842),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_985),
.B(n_866),
.Y(n_1098)
);

NOR4xp25_ASAP7_75t_L g1099 ( 
.A(n_1049),
.B(n_938),
.C(n_942),
.D(n_940),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_970),
.B(n_968),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_SL g1101 ( 
.A1(n_1018),
.A2(n_810),
.B1(n_811),
.B2(n_847),
.C(n_815),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_969),
.A2(n_772),
.B(n_933),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_976),
.B(n_831),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_957),
.A2(n_772),
.B(n_933),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1001),
.A2(n_923),
.A3(n_927),
.B(n_905),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_981),
.A2(n_837),
.B(n_832),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_962),
.A2(n_943),
.B(n_897),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_975),
.A2(n_837),
.B(n_832),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_960),
.A2(n_903),
.B(n_877),
.C(n_876),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_967),
.B(n_785),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1054),
.B(n_825),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1055),
.A2(n_877),
.B(n_876),
.C(n_818),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1077),
.A2(n_847),
.B(n_916),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1077),
.A2(n_916),
.B(n_928),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1029),
.Y(n_1115)
);

OAI22x1_ASAP7_75t_L g1116 ( 
.A1(n_1020),
.A2(n_891),
.B1(n_861),
.B2(n_843),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1002),
.A2(n_829),
.B(n_899),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_973),
.B(n_803),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_1043),
.B(n_820),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_951),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_989),
.B(n_937),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1008),
.A2(n_829),
.B1(n_859),
.B2(n_922),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_961),
.A2(n_944),
.B(n_880),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1042),
.Y(n_1124)
);

NOR4xp25_ASAP7_75t_L g1125 ( 
.A(n_1023),
.B(n_925),
.C(n_898),
.D(n_893),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1070),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_998),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1045),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_1039),
.A2(n_861),
.B1(n_891),
.B2(n_878),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_SL g1130 ( 
.A(n_1010),
.B(n_878),
.C(n_919),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_955),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_961),
.A2(n_1072),
.A3(n_986),
.B(n_994),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1075),
.B(n_897),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_978),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1048),
.B(n_897),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_986),
.A2(n_994),
.B(n_962),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_878),
.B(n_922),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_SL g1139 ( 
.A1(n_1031),
.A2(n_922),
.B(n_1027),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1025),
.A2(n_922),
.B1(n_947),
.B2(n_950),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1073),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_997),
.B(n_996),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1040),
.A2(n_1059),
.B1(n_971),
.B2(n_1061),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_982),
.A2(n_1005),
.B(n_1046),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1063),
.Y(n_1145)
);

NOR4xp25_ASAP7_75t_L g1146 ( 
.A(n_1017),
.B(n_1014),
.C(n_1015),
.D(n_1024),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1052),
.A2(n_1068),
.B(n_983),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1021),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_956),
.B(n_959),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1056),
.B(n_1057),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_983),
.A2(n_963),
.B(n_972),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1058),
.B(n_1006),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1026),
.A2(n_954),
.B(n_984),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_954),
.A2(n_1026),
.B(n_999),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_990),
.B(n_980),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1069),
.B(n_1037),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1022),
.A2(n_1034),
.B(n_1038),
.C(n_1032),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1074),
.A2(n_979),
.B(n_965),
.Y(n_1158)
);

AOI31xp67_ASAP7_75t_L g1159 ( 
.A1(n_1004),
.A2(n_1079),
.A3(n_1012),
.B(n_1067),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1021),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_995),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1050),
.A2(n_966),
.B(n_955),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1051),
.A2(n_1011),
.B(n_1007),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1032),
.A2(n_1033),
.B(n_1076),
.C(n_1016),
.Y(n_1164)
);

NAND3x1_ASAP7_75t_L g1165 ( 
.A(n_1033),
.B(n_992),
.C(n_977),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1065),
.A2(n_1041),
.B(n_945),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_993),
.A2(n_1062),
.A3(n_1075),
.B1(n_1064),
.B2(n_989),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1065),
.A2(n_1041),
.B(n_1078),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1071),
.A2(n_989),
.B(n_993),
.Y(n_1169)
);

AOI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1037),
.A2(n_1071),
.B(n_1036),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1071),
.A2(n_1080),
.B(n_1021),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1080),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1080),
.B(n_1044),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1035),
.A2(n_1047),
.B(n_1053),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1023),
.A2(n_906),
.B(n_1039),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_957),
.A2(n_1066),
.A3(n_953),
.B(n_974),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_967),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_955),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_948),
.A2(n_906),
.B(n_949),
.Y(n_1180)
);

NAND3x1_ASAP7_75t_L g1181 ( 
.A(n_1023),
.B(n_392),
.C(n_562),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_948),
.B(n_598),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1043),
.B(n_820),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_948),
.A2(n_906),
.B(n_949),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_969),
.A2(n_957),
.B(n_906),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_R g1186 ( 
.A(n_1010),
.B(n_506),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_969),
.A2(n_957),
.B(n_906),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_948),
.B(n_598),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1019),
.B(n_658),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_970),
.B(n_906),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_SL g1191 ( 
.A(n_948),
.B(n_913),
.C(n_906),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_957),
.A2(n_961),
.B(n_953),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_948),
.A2(n_906),
.B(n_914),
.C(n_953),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_948),
.A2(n_906),
.B(n_949),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_967),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_987),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1021),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_957),
.A2(n_1002),
.B(n_961),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_970),
.B(n_906),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_948),
.B(n_598),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_987),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_987),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_967),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_968),
.B(n_906),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1075),
.B(n_889),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_969),
.A2(n_957),
.B(n_906),
.Y(n_1211)
);

NAND2x1_ASAP7_75t_L g1212 ( 
.A(n_993),
.B(n_788),
.Y(n_1212)
);

AOI31xp67_ASAP7_75t_L g1213 ( 
.A1(n_954),
.A2(n_706),
.A3(n_595),
.B(n_609),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_978),
.Y(n_1214)
);

O2A1O1Ixp5_ASAP7_75t_SL g1215 ( 
.A1(n_1017),
.A2(n_706),
.B(n_595),
.C(n_902),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_952),
.A2(n_981),
.B(n_975),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1100),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1191),
.A2(n_1184),
.B1(n_1195),
.B2(n_1180),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1180),
.A2(n_1184),
.B1(n_1195),
.B2(n_1188),
.Y(n_1219)
);

NOR3xp33_ASAP7_75t_SL g1220 ( 
.A(n_1186),
.B(n_1144),
.C(n_1175),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1190),
.A2(n_1202),
.B1(n_1182),
.B2(n_1203),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1135),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1086),
.Y(n_1224)
);

NAND2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_1172),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1194),
.A2(n_1188),
.B(n_1182),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1091),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1082),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1083),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1203),
.B(n_1089),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1146),
.A2(n_1157),
.B(n_1164),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_1208),
.B1(n_1089),
.B2(n_1094),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1193),
.A2(n_1216),
.B(n_1209),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1197),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1146),
.A2(n_1112),
.B(n_1211),
.Y(n_1235)
);

OR2x6_ASAP7_75t_L g1236 ( 
.A(n_1119),
.B(n_1183),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1181),
.A2(n_1175),
.B1(n_1156),
.B2(n_1129),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1145),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1204),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1142),
.A2(n_1110),
.B1(n_1097),
.B2(n_1103),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1120),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1137),
.A2(n_1187),
.B(n_1154),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1206),
.Y(n_1243)
);

INVx3_ASAP7_75t_SL g1244 ( 
.A(n_1214),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1149),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1111),
.B(n_1103),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1210),
.B(n_1134),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1137),
.A2(n_1151),
.B(n_1158),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1158),
.A2(n_1201),
.B(n_1205),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1200),
.A2(n_1107),
.B(n_1102),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1179),
.B(n_1152),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1149),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1109),
.A2(n_1140),
.B(n_1215),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1174),
.Y(n_1254)
);

OAI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1143),
.A2(n_1207),
.B1(n_1196),
.B2(n_1189),
.C(n_1099),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1119),
.B(n_1183),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1153),
.A2(n_1092),
.B(n_1088),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1168),
.B(n_1171),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1114),
.A2(n_1104),
.B(n_1123),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1196),
.A2(n_1177),
.B1(n_1136),
.B2(n_1118),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1111),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1096),
.A2(n_1150),
.B(n_1133),
.C(n_1127),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1092),
.A2(n_1099),
.B(n_1165),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1148),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1108),
.A2(n_1113),
.B(n_1106),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1125),
.A2(n_1159),
.B(n_1162),
.Y(n_1266)
);

INVx8_ASAP7_75t_L g1267 ( 
.A(n_1183),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1126),
.A2(n_1090),
.B1(n_1124),
.B2(n_1115),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1163),
.A2(n_1139),
.B(n_1138),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1155),
.Y(n_1270)
);

AO21x1_ASAP7_75t_L g1271 ( 
.A1(n_1122),
.A2(n_1098),
.B(n_1131),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1117),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1212),
.B(n_1166),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1117),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1101),
.A2(n_1098),
.B(n_1122),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1128),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1141),
.A2(n_1161),
.B1(n_1116),
.B2(n_1130),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1125),
.A2(n_1101),
.B(n_1213),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1138),
.A2(n_1199),
.B(n_1169),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1095),
.B(n_1121),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1173),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1199),
.A2(n_1170),
.B(n_1095),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1173),
.B(n_1160),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1192),
.A2(n_1091),
.B(n_1176),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1148),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1167),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1148),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1192),
.A2(n_1093),
.B1(n_1160),
.B2(n_1198),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1093),
.A2(n_1167),
.B(n_1105),
.C(n_1176),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1176),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1160),
.A2(n_1198),
.B1(n_1132),
.B2(n_1105),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1132),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1198),
.B(n_1105),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1132),
.B(n_1119),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1086),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1086),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1086),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1086),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1180),
.A2(n_906),
.B(n_948),
.C(n_1184),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1194),
.A2(n_906),
.B(n_1180),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1086),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1086),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1137),
.A2(n_1087),
.B(n_1185),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1135),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1194),
.A2(n_906),
.B(n_1180),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1191),
.A2(n_906),
.B1(n_913),
.B2(n_511),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1135),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1196),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1086),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1190),
.B(n_1202),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1086),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1100),
.Y(n_1316)
);

INVx8_ASAP7_75t_L g1317 ( 
.A(n_1119),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1086),
.Y(n_1318)
);

AO32x2_ASAP7_75t_L g1319 ( 
.A1(n_1140),
.A2(n_1125),
.A3(n_1122),
.B1(n_1081),
.B2(n_1017),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1186),
.A2(n_913),
.B(n_511),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_SL g1321 ( 
.A(n_1214),
.B(n_506),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1191),
.A2(n_906),
.B1(n_644),
.B2(n_1020),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1191),
.A2(n_906),
.B1(n_644),
.B2(n_1020),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1180),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1086),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1194),
.A2(n_906),
.B(n_1180),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1086),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1191),
.A2(n_906),
.B1(n_644),
.B2(n_1020),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1135),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1190),
.B(n_1202),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1180),
.A2(n_1195),
.B(n_1184),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1190),
.B(n_1202),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1137),
.A2(n_1087),
.B(n_1185),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1135),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1190),
.B(n_1202),
.Y(n_1335)
);

AND2x2_ASAP7_75t_SL g1336 ( 
.A(n_1146),
.B(n_906),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1191),
.A2(n_913),
.B1(n_906),
.B2(n_1175),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1180),
.A2(n_906),
.B(n_948),
.C(n_1184),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1100),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1147),
.A2(n_1085),
.B(n_1178),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1086),
.Y(n_1342)
);

AND2x2_ASAP7_75t_SL g1343 ( 
.A(n_1336),
.B(n_1218),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1310),
.A2(n_1322),
.B1(n_1323),
.B2(n_1328),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1223),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1322),
.A2(n_1323),
.B1(n_1328),
.B2(n_1314),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1222),
.B(n_1230),
.Y(n_1347)
);

AND2x2_ASAP7_75t_SL g1348 ( 
.A(n_1336),
.B(n_1218),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1301),
.A2(n_1338),
.B(n_1254),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1324),
.B(n_1219),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1324),
.B(n_1219),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1337),
.B(n_1335),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1220),
.A2(n_1217),
.B1(n_1339),
.B2(n_1316),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1302),
.B(n_1309),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1266),
.A2(n_1235),
.B(n_1231),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1337),
.A2(n_1301),
.B(n_1338),
.C(n_1255),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1281),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1220),
.A2(n_1260),
.B1(n_1232),
.B2(n_1237),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1326),
.B(n_1286),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1270),
.B(n_1240),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1331),
.B(n_1232),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1261),
.A2(n_1256),
.B(n_1236),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1238),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1330),
.A2(n_1332),
.B1(n_1240),
.B2(n_1320),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1241),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1312),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1263),
.A2(n_1253),
.B(n_1271),
.C(n_1226),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1319),
.B(n_1294),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1227),
.A2(n_1290),
.B(n_1246),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1262),
.A2(n_1251),
.B(n_1261),
.C(n_1236),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1245),
.B(n_1252),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1278),
.A2(n_1269),
.B(n_1279),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1236),
.A2(n_1256),
.B(n_1294),
.C(n_1239),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1250),
.A2(n_1259),
.B(n_1221),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1224),
.B(n_1297),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1280),
.A2(n_1294),
.B(n_1238),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1295),
.A2(n_1307),
.B(n_1341),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1319),
.B(n_1288),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1297),
.B(n_1313),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1340),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1287),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1313),
.B(n_1315),
.Y(n_1382)
);

OA22x2_ASAP7_75t_L g1383 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_1234),
.B2(n_1342),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1223),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1315),
.B(n_1283),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1296),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_SL g1387 ( 
.A(n_1329),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1298),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1319),
.B(n_1293),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1267),
.B(n_1317),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1293),
.B(n_1275),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1299),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1283),
.B(n_1276),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1303),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1304),
.B(n_1318),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_L g1396 ( 
.A(n_1325),
.B(n_1327),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1268),
.B(n_1275),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1275),
.B(n_1247),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1292),
.A2(n_1274),
.B(n_1272),
.C(n_1277),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1267),
.B(n_1317),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1233),
.A2(n_1274),
.B(n_1292),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_SL g1402 ( 
.A1(n_1311),
.A2(n_1267),
.B(n_1317),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1321),
.A2(n_1289),
.B(n_1244),
.C(n_1225),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1248),
.A2(n_1289),
.B(n_1242),
.C(n_1305),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1291),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1258),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1282),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1242),
.B(n_1244),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1287),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1311),
.A2(n_1334),
.B(n_1306),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_SL g1412 ( 
.A1(n_1306),
.A2(n_1334),
.B(n_1273),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1280),
.A2(n_1242),
.B(n_1333),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1285),
.A2(n_1264),
.B(n_1257),
.C(n_1284),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1273),
.A2(n_1265),
.B(n_1249),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1222),
.B(n_1230),
.Y(n_1417)
);

O2A1O1Ixp5_ASAP7_75t_L g1418 ( 
.A1(n_1231),
.A2(n_906),
.B(n_1235),
.C(n_1194),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1324),
.B(n_1175),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1301),
.A2(n_906),
.B(n_1180),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1301),
.A2(n_1338),
.B(n_906),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1222),
.B(n_1230),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1229),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1229),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1324),
.B(n_1175),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1415),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1383),
.Y(n_1429)
);

OAI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1344),
.A2(n_1346),
.B1(n_1418),
.B2(n_1420),
.C(n_1352),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1391),
.B(n_1389),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1383),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1387),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1414),
.A2(n_1416),
.B(n_1413),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1347),
.B(n_1417),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1414),
.A2(n_1407),
.B(n_1422),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1423),
.B(n_1354),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1401),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1362),
.B(n_1376),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1391),
.B(n_1389),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1409),
.B(n_1406),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1368),
.B(n_1378),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1398),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1361),
.A2(n_1354),
.B(n_1405),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1373),
.B(n_1406),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1355),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1355),
.B(n_1408),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1361),
.B(n_1350),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1356),
.A2(n_1349),
.B(n_1360),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1352),
.A2(n_1358),
.B1(n_1348),
.B2(n_1343),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1404),
.A2(n_1367),
.B(n_1399),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1372),
.A2(n_1374),
.B(n_1369),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1397),
.A2(n_1351),
.B(n_1424),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1425),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1355),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1421),
.B(n_1359),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1359),
.B(n_1343),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1419),
.B(n_1427),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1348),
.B(n_1372),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1388),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1386),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1394),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1375),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1371),
.B(n_1392),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1379),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1382),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1353),
.A2(n_1364),
.B1(n_1357),
.B2(n_1365),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1447),
.B(n_1454),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1437),
.B(n_1385),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1433),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1437),
.B(n_1448),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.B(n_1380),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1455),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1455),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1431),
.B(n_1374),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1431),
.B(n_1380),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1440),
.B(n_1380),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1455),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1453),
.A2(n_1396),
.B(n_1395),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1435),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1428),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1377),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1465),
.B(n_1461),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1462),
.B(n_1454),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1435),
.B(n_1393),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1458),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1430),
.B(n_1370),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1382),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1454),
.B(n_1377),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1492),
.A2(n_1430),
.B1(n_1450),
.B2(n_1471),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1493),
.B(n_1486),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1492),
.A2(n_1450),
.B1(n_1471),
.B2(n_1459),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1485),
.A2(n_1451),
.B1(n_1450),
.B2(n_1460),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1478),
.Y(n_1499)
);

AND2x4_ASAP7_75t_SL g1500 ( 
.A(n_1493),
.B(n_1439),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1490),
.A2(n_1451),
.B1(n_1439),
.B2(n_1459),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1489),
.A2(n_1459),
.B(n_1403),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1489),
.A2(n_1450),
.B(n_1456),
.C(n_1446),
.Y(n_1503)
);

AOI33xp33_ASAP7_75t_L g1504 ( 
.A1(n_1494),
.A2(n_1366),
.A3(n_1429),
.B1(n_1432),
.B2(n_1464),
.B3(n_1466),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1485),
.A2(n_1450),
.B1(n_1439),
.B2(n_1432),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

OAI211xp5_ASAP7_75t_L g1507 ( 
.A1(n_1490),
.A2(n_1456),
.B(n_1429),
.C(n_1468),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1474),
.A2(n_1439),
.B1(n_1390),
.B2(n_1476),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1493),
.B(n_1441),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1472),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_R g1511 ( 
.A(n_1475),
.B(n_1345),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

AOI33xp33_ASAP7_75t_L g1513 ( 
.A1(n_1494),
.A2(n_1466),
.A3(n_1464),
.B1(n_1467),
.B2(n_1469),
.B3(n_1457),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1476),
.A2(n_1439),
.B1(n_1460),
.B2(n_1445),
.Y(n_1514)
);

OAI31xp33_ASAP7_75t_L g1515 ( 
.A1(n_1489),
.A2(n_1460),
.A3(n_1468),
.B(n_1463),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1486),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1345),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1479),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1475),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1488),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1489),
.A2(n_1444),
.B1(n_1449),
.B2(n_1463),
.C(n_1443),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1493),
.A2(n_1439),
.B1(n_1444),
.B2(n_1445),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1472),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1473),
.A2(n_1384),
.B1(n_1400),
.B2(n_1445),
.C(n_1363),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1494),
.A2(n_1444),
.B1(n_1449),
.B2(n_1443),
.C(n_1470),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1493),
.B(n_1470),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1493),
.B(n_1467),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1483),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1473),
.B(n_1469),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1484),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1503),
.B(n_1445),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1511),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1496),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1499),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1500),
.B(n_1491),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1512),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1525),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1510),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1517),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1532),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1533),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_L g1550 ( 
.A(n_1495),
.B(n_1384),
.C(n_1473),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1526),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1500),
.B(n_1509),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1535),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1513),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1536),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1513),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1516),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1528),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1522),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1522),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1535),
.B(n_1440),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1536),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1524),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1534),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1540),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1554),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1550),
.A2(n_1497),
.B(n_1505),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1554),
.A2(n_1521),
.B1(n_1529),
.B2(n_1503),
.C(n_1498),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1539),
.B(n_1509),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1556),
.B(n_1482),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1546),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1546),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1539),
.B(n_1509),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1502),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1557),
.Y(n_1582)
);

INVx4_ASAP7_75t_L g1583 ( 
.A(n_1537),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1561),
.B(n_1504),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1562),
.Y(n_1586)
);

BUFx4f_ASAP7_75t_SL g1587 ( 
.A(n_1542),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1520),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1482),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1541),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1551),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1543),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1544),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1551),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1544),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1564),
.B(n_1481),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1545),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1545),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1548),
.B(n_1504),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1601),
.B(n_1566),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1578),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1578),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1581),
.B(n_1559),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1567),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1582),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1569),
.B(n_1560),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1537),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1569),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1586),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1573),
.B(n_1537),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1587),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1568),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1571),
.B(n_1537),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1590),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1549),
.Y(n_1623)
);

OAI31xp33_ASAP7_75t_L g1624 ( 
.A1(n_1570),
.A2(n_1501),
.A3(n_1507),
.B(n_1514),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1549),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1572),
.B(n_1576),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1590),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1574),
.B(n_1480),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1579),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1574),
.B(n_1480),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1577),
.B(n_1530),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1589),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1570),
.B(n_1530),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1584),
.B(n_1487),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1591),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1626),
.B(n_1572),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1626),
.B(n_1576),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1634),
.A2(n_1583),
.B1(n_1523),
.B2(n_1527),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1611),
.A2(n_1583),
.B1(n_1508),
.B2(n_1434),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1619),
.B(n_1580),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1580),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1624),
.A2(n_1583),
.B1(n_1434),
.B2(n_1589),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1624),
.A2(n_1583),
.B1(n_1434),
.B2(n_1594),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1588),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1604),
.A2(n_1434),
.B1(n_1436),
.B2(n_1452),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1612),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1608),
.B(n_1592),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1610),
.B(n_1588),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1612),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1598),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1633),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1614),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1615),
.B(n_1598),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1633),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1617),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1646),
.A2(n_1631),
.B(n_1629),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1659),
.Y(n_1664)
);

AOI32xp33_ASAP7_75t_L g1665 ( 
.A1(n_1645),
.A2(n_1635),
.A3(n_1606),
.B1(n_1615),
.B2(n_1618),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1662),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1662),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1656),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1639),
.A2(n_1623),
.B1(n_1602),
.B2(n_1609),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1657),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1647),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1657),
.Y(n_1672)
);

AOI322xp5_ASAP7_75t_L g1673 ( 
.A1(n_1640),
.A2(n_1632),
.A3(n_1621),
.B1(n_1618),
.B2(n_1628),
.C1(n_1627),
.C2(n_1620),
.Y(n_1673)
);

OAI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1640),
.A2(n_1602),
.B1(n_1623),
.B2(n_1625),
.C(n_1636),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1656),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1625),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1617),
.C(n_1620),
.Y(n_1678)
);

AOI221x1_ASAP7_75t_L g1679 ( 
.A1(n_1643),
.A2(n_1636),
.B1(n_1628),
.B2(n_1627),
.C(n_1630),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1661),
.B(n_1618),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1642),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1671),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1664),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1664),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1666),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1681),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1667),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1675),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1672),
.B(n_1637),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1642),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1683),
.Y(n_1692)
);

NAND4xp25_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1669),
.C(n_1663),
.D(n_1665),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_SL g1695 ( 
.A(n_1684),
.B(n_1680),
.Y(n_1695)
);

OAI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1689),
.A2(n_1669),
.B(n_1673),
.C(n_1680),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_SL g1697 ( 
.A(n_1691),
.B(n_1674),
.C(n_1678),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1685),
.A2(n_1677),
.B1(n_1648),
.B2(n_1654),
.C(n_1643),
.Y(n_1698)
);

NOR3x1_ASAP7_75t_L g1699 ( 
.A(n_1690),
.B(n_1650),
.C(n_1648),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1691),
.A2(n_1679),
.B(n_1684),
.Y(n_1700)
);

AOI322xp5_ASAP7_75t_L g1701 ( 
.A1(n_1697),
.A2(n_1687),
.A3(n_1688),
.B1(n_1668),
.B2(n_1676),
.C1(n_1683),
.C2(n_1650),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1694),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1696),
.A2(n_1654),
.B(n_1652),
.C(n_1651),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1695),
.B(n_1653),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1693),
.A2(n_1651),
.B1(n_1652),
.B2(n_1659),
.C(n_1658),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1702),
.B(n_1700),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1704),
.B(n_1692),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1703),
.A2(n_1698),
.B(n_1658),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1701),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1705),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.Y(n_1711)
);

NAND4xp75_ASAP7_75t_L g1712 ( 
.A(n_1706),
.B(n_1699),
.C(n_1653),
.D(n_1641),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1709),
.A2(n_1411),
.B(n_1519),
.C(n_1603),
.Y(n_1713)
);

OAI321xp33_ASAP7_75t_L g1714 ( 
.A1(n_1707),
.A2(n_1638),
.A3(n_1660),
.B1(n_1655),
.B2(n_1644),
.C(n_1649),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1711),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1710),
.B(n_1659),
.Y(n_1716)
);

NAND4xp25_ASAP7_75t_L g1717 ( 
.A(n_1713),
.B(n_1708),
.C(n_1659),
.D(n_1644),
.Y(n_1717)
);

NAND4xp75_ASAP7_75t_L g1718 ( 
.A(n_1716),
.B(n_1660),
.C(n_1655),
.D(n_1603),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1712),
.B(n_1605),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1717),
.B(n_1715),
.C(n_1714),
.Y(n_1720)
);

AOI322xp5_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1719),
.A3(n_1718),
.B1(n_1649),
.B2(n_1605),
.C1(n_1622),
.C2(n_1630),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1721),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1721),
.A2(n_1622),
.B1(n_1555),
.B2(n_1563),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_L g1724 ( 
.A(n_1722),
.B(n_1410),
.C(n_1381),
.D(n_1363),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1723),
.B(n_1593),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1725),
.Y(n_1726)
);

CKINVDCx20_ASAP7_75t_R g1727 ( 
.A(n_1724),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1593),
.B1(n_1596),
.B2(n_1579),
.Y(n_1728)
);

AOI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1727),
.B(n_1381),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1729),
.B(n_1596),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_R g1731 ( 
.A1(n_1730),
.A2(n_1412),
.B1(n_1579),
.B2(n_1402),
.C(n_1600),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1600),
.B1(n_1595),
.B2(n_1597),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1410),
.B(n_1599),
.C(n_1597),
.Y(n_1733)
);


endmodule