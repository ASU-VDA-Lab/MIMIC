module fake_jpeg_21864_n_271 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_53),
.B1(n_17),
.B2(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_15),
.B(n_27),
.C(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_72),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_27),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_0),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_27),
.B1(n_36),
.B2(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_70),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_38),
.B1(n_17),
.B2(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2x1_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_28),
.B1(n_25),
.B2(n_24),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_20),
.B1(n_28),
.B2(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_82),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_89),
.B1(n_78),
.B2(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_96),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_44),
.B1(n_55),
.B2(n_57),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_51),
.B1(n_40),
.B2(n_26),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_75),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_35),
.Y(n_96)
);

AO21x2_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_54),
.B(n_47),
.Y(n_98)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_63),
.B1(n_67),
.B2(n_74),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_26),
.B(n_73),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_71),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_68),
.B1(n_59),
.B2(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_87),
.B1(n_82),
.B2(n_85),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_92),
.B1(n_86),
.B2(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_88),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_121),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_60),
.B(n_72),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_118),
.B(n_63),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_97),
.B1(n_89),
.B2(n_64),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_84),
.B1(n_65),
.B2(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_124),
.B(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_127),
.B1(n_138),
.B2(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_87),
.B1(n_97),
.B2(n_98),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_106),
.B1(n_108),
.B2(n_116),
.Y(n_156)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_98),
.A3(n_86),
.B1(n_92),
.B2(n_99),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_98),
.B(n_83),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_114),
.B(n_76),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_100),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_143),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_143),
.B(n_144),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_104),
.B(n_108),
.C(n_115),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_99),
.B(n_80),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_156),
.B(n_159),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_151),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_119),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_118),
.B1(n_103),
.B2(n_121),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_112),
.B1(n_106),
.B2(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_167),
.B1(n_140),
.B2(n_131),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_115),
.A3(n_114),
.B1(n_112),
.B2(n_110),
.C1(n_105),
.C2(n_58),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_42),
.C(n_40),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_76),
.C(n_46),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_127),
.C(n_130),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_50),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_16),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_65),
.B1(n_50),
.B2(n_39),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_176),
.B1(n_155),
.B2(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_177),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_187),
.Y(n_204)
);

AND2x4_ASAP7_75t_SL g174 ( 
.A(n_151),
.B(n_136),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_160),
.B(n_166),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_146),
.B(n_123),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_123),
.C(n_124),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_122),
.B1(n_65),
.B2(n_24),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_182),
.B1(n_167),
.B2(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_42),
.C(n_77),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_22),
.B(n_19),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_185),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_77),
.C(n_20),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_77),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_77),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_188),
.A2(n_152),
.B1(n_154),
.B2(n_16),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_164),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_165),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_203),
.C(n_205),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_156),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_169),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_178),
.C(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_152),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_22),
.B1(n_16),
.B2(n_2),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_168),
.B1(n_174),
.B2(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_173),
.C(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_184),
.C(n_174),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_172),
.C(n_13),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_220),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_13),
.B(n_12),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_221),
.B(n_2),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_12),
.C(n_1),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_208),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_194),
.B1(n_200),
.B2(n_195),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_226),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_213),
.A2(n_198),
.B(n_202),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_227),
.B(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_204),
.B1(n_189),
.B2(n_3),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_1),
.B(n_2),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_4),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_3),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_11),
.C(n_8),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_3),
.B(n_4),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_214),
.C(n_5),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_239),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_223),
.C(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_241),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_227),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_4),
.C(n_5),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_6),
.C(n_7),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_6),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_235),
.C(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_255),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_230),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_252),
.B(n_7),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_249),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_234),
.B(n_232),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_7),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_9),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_259),
.B(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_9),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_253),
.B(n_251),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_265),
.B(n_253),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_264),
.B1(n_10),
.B2(n_11),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_266),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_10),
.B1(n_11),
.B2(n_266),
.Y(n_271)
);


endmodule