module fake_jpeg_5591_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_15),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_10),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_20),
.B1(n_50),
.B2(n_43),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_65),
.B1(n_72),
.B2(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_34),
.B1(n_28),
.B2(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_62),
.B1(n_53),
.B2(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_38),
.B1(n_29),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_29),
.B1(n_38),
.B2(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_33),
.B1(n_37),
.B2(n_30),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_16),
.B1(n_39),
.B2(n_25),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_85),
.B(n_109),
.C(n_96),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_86),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_37),
.B1(n_39),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_92),
.B1(n_105),
.B2(n_88),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_36),
.B1(n_32),
.B2(n_18),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_89),
.B1(n_93),
.B2(n_88),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_31),
.B(n_11),
.C(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_18),
.B1(n_39),
.B2(n_4),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_44),
.A2(n_31),
.B1(n_11),
.B2(n_4),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_100),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_97),
.B1(n_108),
.B2(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_67),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_51),
.B1(n_43),
.B2(n_20),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_62),
.B(n_21),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_112),
.Y(n_153)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_123),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_121),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_81),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_138),
.B1(n_94),
.B2(n_68),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_91),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_145),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_72),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_142),
.Y(n_172)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_133),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_74),
.B(n_83),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_73),
.Y(n_140)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_78),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_98),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_120),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_149),
.A2(n_169),
.B(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_86),
.B1(n_80),
.B2(n_71),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_160),
.B1(n_165),
.B2(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_179),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_181),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_103),
.B1(n_106),
.B2(n_99),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_143),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_114),
.B1(n_139),
.B2(n_116),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_142),
.B(n_145),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_118),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_142),
.B1(n_118),
.B2(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_112),
.B1(n_127),
.B2(n_131),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_150),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_119),
.C(n_135),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_182),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_143),
.B(n_125),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_192),
.B(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_125),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_125),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_199),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_132),
.B(n_148),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_208),
.B(n_212),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_151),
.A2(n_132),
.B1(n_179),
.B2(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_170),
.B(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_207),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_151),
.B1(n_148),
.B2(n_162),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_210),
.B1(n_180),
.B2(n_155),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_164),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_148),
.A2(n_158),
.B1(n_147),
.B2(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_186),
.B1(n_187),
.B2(n_208),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_147),
.B(n_174),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_226),
.B(n_228),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_232),
.B1(n_236),
.B2(n_231),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_146),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_240),
.C(n_237),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_150),
.B1(n_178),
.B2(n_175),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_175),
.B(n_188),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_192),
.B(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_182),
.B1(n_183),
.B2(n_210),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_232),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_207),
.B1(n_211),
.B2(n_183),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_190),
.B1(n_197),
.B2(n_185),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_184),
.B1(n_202),
.B2(n_199),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_239),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_201),
.A3(n_194),
.B1(n_184),
.B2(n_214),
.C1(n_202),
.C2(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_252),
.B1(n_240),
.B2(n_217),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_259),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_236),
.C(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_219),
.Y(n_254)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_254),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_225),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_230),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_257),
.Y(n_264)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_216),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_SL g259 ( 
.A(n_228),
.B(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_235),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_269),
.Y(n_287)
);

AOI22x1_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_234),
.B1(n_216),
.B2(n_235),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_271),
.B1(n_243),
.B2(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_257),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_243),
.B1(n_249),
.B2(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_215),
.B1(n_227),
.B2(n_249),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_269),
.CI(n_274),
.CON(n_293),
.SN(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_244),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_277),
.B(n_247),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_273),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_252),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_285),
.B(n_291),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_246),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_251),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_262),
.B(n_256),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_294),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_287),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_285),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_260),
.B1(n_267),
.B2(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_300),
.B1(n_280),
.B2(n_271),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_260),
.B1(n_278),
.B2(n_245),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_263),
.B(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_242),
.C(n_276),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_307),
.C(n_309),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_301),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_287),
.C(n_266),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_250),
.C(n_299),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_302),
.B1(n_295),
.B2(n_283),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_276),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_308),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_319),
.CI(n_316),
.CON(n_320),
.SN(n_320)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_321),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_314),
.B(n_313),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_312),
.Y(n_325)
);


endmodule