module fake_aes_4325_n_894 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_894);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_894;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_769;
wire n_818;
wire n_844;
wire n_725;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_703;
wire n_394;
wire n_813;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_685;
wire n_362;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_522;
wire n_883;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_763;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
CKINVDCx16_ASAP7_75t_R g275 ( .A(n_250), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_246), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_62), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_238), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_40), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_189), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_223), .Y(n_285) );
BUFx10_ASAP7_75t_L g286 ( .A(n_202), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_180), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_5), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_104), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_220), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_212), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_11), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_156), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_82), .Y(n_294) );
BUFx10_ASAP7_75t_L g295 ( .A(n_4), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_143), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_69), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_137), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_199), .B(n_217), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_7), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_83), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_157), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_90), .Y(n_305) );
CKINVDCx14_ASAP7_75t_R g306 ( .A(n_164), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_79), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_158), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_89), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_86), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_123), .B(n_95), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_222), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_248), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_51), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_152), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_61), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_197), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_257), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_249), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_55), .Y(n_321) );
INVxp33_ASAP7_75t_SL g322 ( .A(n_150), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_106), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_118), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_195), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_71), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_253), .Y(n_327) );
BUFx5_ASAP7_75t_L g328 ( .A(n_186), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_149), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_213), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_43), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_147), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_65), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_98), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_59), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_107), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_121), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_75), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_53), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_228), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_270), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_172), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_145), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_256), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_174), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_141), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_165), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_138), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_160), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_193), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_201), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_97), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_117), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_35), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_48), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_155), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_251), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_72), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_10), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_261), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_178), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_4), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_148), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_46), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_263), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_255), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_221), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_260), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_264), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_227), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_274), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_20), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_244), .Y(n_374) );
BUFx5_ASAP7_75t_L g375 ( .A(n_182), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_215), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_32), .Y(n_377) );
BUFx10_ASAP7_75t_L g378 ( .A(n_33), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_47), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_56), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_198), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_262), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_146), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_247), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_142), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_266), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_92), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_105), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_27), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_58), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_81), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_205), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_34), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_94), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_168), .Y(n_395) );
BUFx5_ASAP7_75t_L g396 ( .A(n_170), .Y(n_396) );
BUFx10_ASAP7_75t_L g397 ( .A(n_134), .Y(n_397) );
BUFx12f_ASAP7_75t_L g398 ( .A(n_286), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_288), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_328), .Y(n_400) );
BUFx12f_ASAP7_75t_L g401 ( .A(n_378), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_328), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_276), .B(n_0), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_338), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_292), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_328), .Y(n_406) );
AND2x6_ASAP7_75t_L g407 ( .A(n_277), .B(n_19), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_328), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_397), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_283), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_343), .B(n_3), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_302), .B(n_5), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_279), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_280), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_295), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_360), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_398), .B(n_363), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_412), .A2(n_322), .B1(n_306), .B2(n_315), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_410), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_404), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_415), .Y(n_423) );
AND2x6_ASAP7_75t_L g424 ( .A(n_403), .B(n_281), .Y(n_424) );
INVx4_ASAP7_75t_L g425 ( .A(n_407), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_413), .B(n_275), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_413), .B(n_414), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_414), .B(n_305), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_412), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_409), .B(n_327), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_416), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
BUFx10_ASAP7_75t_L g434 ( .A(n_403), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_408), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_431), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_425), .B(n_434), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_425), .B(n_411), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_426), .B(n_411), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_431), .Y(n_440) );
INVx4_ASAP7_75t_L g441 ( .A(n_424), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_428), .B(n_409), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_427), .B(n_429), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_424), .B(n_416), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_419), .B(n_278), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_422), .B(n_282), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_418), .B(n_415), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_430), .B(n_304), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_420), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_423), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_418), .B(n_401), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_424), .B(n_316), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_435), .Y(n_453) );
NAND2xp33_ASAP7_75t_L g454 ( .A(n_424), .B(n_407), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_432), .B(n_405), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_421), .B(n_407), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_421), .B(n_405), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_445), .A2(n_331), .B1(n_350), .B2(n_323), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_443), .B(n_407), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_441), .B(n_284), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_439), .B(n_399), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_441), .B(n_289), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_442), .B(n_399), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_440), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_444), .B(n_300), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_448), .B(n_376), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_452), .A2(n_402), .B1(n_417), .B2(n_329), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_448), .B(n_402), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_454), .A2(n_301), .B(n_417), .Y(n_470) );
INVx5_ASAP7_75t_L g471 ( .A(n_450), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_451), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_438), .A2(n_287), .B1(n_291), .B2(n_290), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_446), .B(n_6), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_455), .B(n_307), .Y(n_475) );
AO21x1_ASAP7_75t_L g476 ( .A1(n_456), .A2(n_296), .B(n_294), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_455), .B(n_309), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_449), .A2(n_298), .B(n_297), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_447), .B(n_354), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_437), .A2(n_382), .B(n_314), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_436), .A2(n_317), .B(n_318), .C(n_313), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_460), .A2(n_457), .B(n_320), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_470), .A2(n_457), .B(n_321), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_471), .B(n_310), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g485 ( .A1(n_467), .A2(n_325), .B(n_312), .Y(n_485) );
OAI21x1_ASAP7_75t_L g486 ( .A1(n_476), .A2(n_324), .B(n_319), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_462), .B(n_332), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_464), .B(n_334), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_472), .B(n_6), .Y(n_489) );
OAI21x1_ASAP7_75t_L g490 ( .A1(n_478), .A2(n_344), .B(n_341), .Y(n_490) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_480), .A2(n_348), .B(n_346), .Y(n_491) );
OAI21x1_ASAP7_75t_L g492 ( .A1(n_459), .A2(n_355), .B(n_352), .Y(n_492) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_469), .A2(n_357), .B(n_356), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_475), .A2(n_362), .B(n_361), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_465), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_471), .Y(n_497) );
AOI211x1_ASAP7_75t_L g498 ( .A1(n_468), .A2(n_366), .B(n_367), .C(n_364), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_481), .B(n_369), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_477), .A2(n_371), .B(n_370), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_466), .A2(n_374), .B(n_372), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_471), .B(n_293), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_461), .A2(n_379), .B(n_377), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_463), .B(n_381), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_473), .A2(n_386), .B(n_388), .C(n_384), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_479), .Y(n_506) );
AOI221x1_ASAP7_75t_L g507 ( .A1(n_458), .A2(n_392), .B1(n_389), .B2(n_410), .C(n_299), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_470), .A2(n_308), .B(n_303), .Y(n_509) );
AOI31xp67_ASAP7_75t_L g510 ( .A1(n_460), .A2(n_330), .A3(n_380), .B(n_333), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_509), .A2(n_311), .B(n_375), .Y(n_512) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_486), .A2(n_336), .B(n_335), .Y(n_513) );
OAI221xp5_ASAP7_75t_SL g514 ( .A1(n_495), .A2(n_347), .B1(n_391), .B2(n_393), .C(n_394), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_506), .B(n_8), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_506), .A2(n_326), .B1(n_339), .B2(n_337), .Y(n_516) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_490), .A2(n_342), .B(n_340), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_497), .Y(n_518) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_492), .A2(n_482), .B(n_491), .Y(n_519) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_507), .A2(n_349), .B(n_345), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_496), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_506), .B(n_9), .Y(n_522) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_483), .A2(n_396), .B(n_375), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_502), .Y(n_524) );
BUFx2_ASAP7_75t_SL g525 ( .A(n_489), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_485), .B(n_351), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_504), .A2(n_375), .B1(n_396), .B2(n_387), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_508), .B(n_9), .Y(n_528) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_493), .A2(n_503), .B(n_500), .Y(n_529) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_510), .A2(n_358), .B(n_353), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_511), .B(n_359), .Y(n_531) );
AOI21x1_ASAP7_75t_L g532 ( .A1(n_493), .A2(n_396), .B(n_387), .Y(n_532) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_494), .A2(n_396), .B(n_387), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_498), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_488), .A2(n_487), .B(n_501), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_504), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_499), .B(n_12), .Y(n_537) );
NAND2xp33_ASAP7_75t_L g538 ( .A(n_505), .B(n_368), .Y(n_538) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_497), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_509), .A2(n_283), .B(n_285), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_495), .B(n_12), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_484), .B(n_283), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_506), .B(n_373), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_508), .B(n_13), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_494), .A2(n_365), .B(n_285), .C(n_383), .Y(n_546) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_509), .A2(n_390), .B(n_385), .Y(n_547) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_509), .A2(n_365), .B(n_421), .Y(n_548) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_509), .A2(n_433), .B(n_22), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_506), .B(n_395), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_508), .B(n_13), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_482), .A2(n_433), .B(n_23), .Y(n_552) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_509), .A2(n_433), .B(n_24), .Y(n_553) );
AO31x2_ASAP7_75t_L g554 ( .A1(n_507), .A2(n_25), .A3(n_26), .B(n_21), .Y(n_554) );
OAI21x1_ASAP7_75t_L g555 ( .A1(n_509), .A2(n_29), .B(n_28), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_508), .B(n_14), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_534), .Y(n_558) );
INVx3_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_556), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_542), .Y(n_561) );
OR2x6_ASAP7_75t_L g562 ( .A(n_528), .B(n_14), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_528), .B(n_15), .Y(n_563) );
INVx5_ASAP7_75t_L g564 ( .A(n_524), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_551), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_545), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_551), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_515), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_539), .Y(n_569) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_532), .A2(n_31), .B(n_30), .Y(n_570) );
NAND2xp33_ASAP7_75t_L g571 ( .A(n_543), .B(n_537), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_541), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_532), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_535), .A2(n_16), .B(n_17), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_522), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_518), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_536), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_540), .B(n_16), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_544), .B(n_17), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_529), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_550), .B(n_18), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_513), .Y(n_585) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_548), .A2(n_18), .B(n_36), .Y(n_586) );
AO21x2_ASAP7_75t_L g587 ( .A1(n_512), .A2(n_37), .B(n_38), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_520), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_523), .B(n_39), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_526), .B(n_41), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_553), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_531), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_527), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_520), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_547), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_547), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_546), .A2(n_42), .B(n_44), .Y(n_599) );
OR2x6_ASAP7_75t_L g600 ( .A(n_519), .B(n_45), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_516), .B(n_49), .Y(n_601) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_552), .A2(n_50), .B(n_52), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_538), .A2(n_54), .B1(n_57), .B2(n_60), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_554), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_530), .B(n_63), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_530), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_514), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_553), .Y(n_611) );
AO21x2_ASAP7_75t_L g612 ( .A1(n_532), .A2(n_64), .B(n_66), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_524), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_534), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_521), .B(n_67), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_535), .A2(n_68), .B(n_70), .Y(n_617) );
INVx11_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_541), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_534), .B(n_73), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_521), .Y(n_621) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_541), .A2(n_74), .B(n_76), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_521), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_521), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_521), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_521), .Y(n_627) );
BUFx3_ASAP7_75t_L g628 ( .A(n_524), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_557), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_569), .B(n_77), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_621), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_618), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_577), .B(n_273), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_568), .B(n_78), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_564), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_609), .A2(n_80), .B1(n_84), .B2(n_85), .C(n_87), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_562), .B(n_88), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_623), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_624), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_625), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_564), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_564), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_563), .B(n_91), .Y(n_645) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_626), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_627), .B(n_93), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_561), .B(n_96), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_575), .B(n_272), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_579), .B(n_99), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_562), .B(n_100), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_615), .Y(n_652) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_588), .Y(n_653) );
AND2x4_ASAP7_75t_L g654 ( .A(n_565), .B(n_101), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_578), .B(n_271), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_560), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_567), .B(n_102), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_562), .B(n_103), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_600), .B(n_108), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_564), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_566), .Y(n_661) );
AO31x2_ASAP7_75t_L g662 ( .A1(n_606), .A2(n_109), .A3(n_110), .B(n_111), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_620), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_580), .B(n_112), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_614), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_620), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_595), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_581), .B(n_116), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_574), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_596), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_583), .B(n_119), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_600), .A2(n_120), .B(n_122), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_574), .Y(n_673) );
INVx3_ASAP7_75t_L g674 ( .A(n_628), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_616), .B(n_124), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_584), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_559), .B(n_269), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_594), .B(n_125), .Y(n_678) );
OAI33xp33_ASAP7_75t_L g679 ( .A1(n_597), .A2(n_126), .A3(n_127), .B1(n_128), .B2(n_129), .B3(n_130), .Y(n_679) );
OAI21x1_ASAP7_75t_L g680 ( .A1(n_582), .A2(n_131), .B(n_132), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_559), .B(n_133), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_613), .B(n_135), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_591), .B(n_136), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_590), .B(n_139), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_573), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_592), .B(n_140), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_604), .Y(n_687) );
INVx3_ASAP7_75t_L g688 ( .A(n_601), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_585), .B(n_144), .Y(n_689) );
INVxp33_ASAP7_75t_L g690 ( .A(n_603), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_588), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_598), .B(n_268), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_607), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_586), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_571), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_573), .B(n_151), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_608), .B(n_267), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_617), .A2(n_153), .B1(n_154), .B2(n_159), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_605), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_582), .B(n_161), .Y(n_700) );
AO21x2_ASAP7_75t_L g701 ( .A1(n_610), .A2(n_162), .B(n_163), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_599), .B(n_166), .Y(n_702) );
OA332x1_ASAP7_75t_L g703 ( .A1(n_617), .A2(n_167), .A3(n_169), .B1(n_171), .B2(n_173), .B3(n_175), .C1(n_176), .C2(n_177), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_612), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_587), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_587), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_589), .B(n_179), .Y(n_708) );
AND2x4_ASAP7_75t_SL g709 ( .A(n_576), .B(n_181), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_642), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_656), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_630), .B(n_593), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_629), .B(n_612), .Y(n_714) );
INVx4_ASAP7_75t_L g715 ( .A(n_636), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_637), .B(n_593), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_661), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_646), .B(n_611), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_632), .B(n_599), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_640), .B(n_572), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_641), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_652), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_676), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_637), .B(n_619), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_665), .B(n_570), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_663), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_688), .B(n_570), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_630), .B(n_666), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_690), .B(n_602), .Y(n_729) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_685), .Y(n_730) );
NAND2x1p5_ASAP7_75t_L g731 ( .A(n_659), .B(n_622), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_685), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_669), .B(n_183), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_674), .B(n_184), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_631), .B(n_185), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_633), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_631), .B(n_187), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_691), .Y(n_738) );
BUFx3_ASAP7_75t_L g739 ( .A(n_660), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_687), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_687), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_634), .B(n_188), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_695), .B(n_190), .Y(n_743) );
BUFx3_ASAP7_75t_L g744 ( .A(n_643), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_647), .B(n_191), .Y(n_745) );
BUFx3_ASAP7_75t_L g746 ( .A(n_644), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_699), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_645), .B(n_192), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_659), .B(n_194), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_693), .B(n_196), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_653), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_651), .B(n_203), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_699), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_658), .B(n_204), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_639), .B(n_206), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_673), .B(n_207), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_694), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_696), .Y(n_758) );
BUFx3_ASAP7_75t_L g759 ( .A(n_635), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_655), .Y(n_760) );
INVx2_ASAP7_75t_SL g761 ( .A(n_682), .Y(n_761) );
BUFx2_ASAP7_75t_L g762 ( .A(n_635), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_704), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_668), .B(n_208), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_706), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_707), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_700), .B(n_209), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_664), .B(n_210), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_671), .B(n_211), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_683), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_705), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_649), .Y(n_772) );
INVxp33_ASAP7_75t_L g773 ( .A(n_744), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_710), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_711), .B(n_654), .Y(n_775) );
AND2x4_ASAP7_75t_L g776 ( .A(n_730), .B(n_709), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_738), .B(n_662), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_721), .B(n_654), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_722), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_751), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_726), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_728), .B(n_712), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_758), .B(n_657), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_729), .B(n_662), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_710), .Y(n_785) );
INVx2_ASAP7_75t_SL g786 ( .A(n_744), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_717), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_746), .B(n_675), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_718), .B(n_686), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_736), .B(n_648), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_730), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_723), .Y(n_792) );
INVx4_ASAP7_75t_L g793 ( .A(n_715), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_746), .B(n_675), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_762), .B(n_681), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_729), .B(n_662), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_753), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_760), .B(n_689), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_719), .B(n_714), .Y(n_799) );
INVxp67_ASAP7_75t_L g800 ( .A(n_727), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_720), .B(n_692), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_732), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_740), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_740), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_741), .Y(n_805) );
NOR2x1_ASAP7_75t_L g806 ( .A(n_715), .B(n_739), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_747), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_772), .B(n_684), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_723), .B(n_708), .Y(n_809) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_759), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_739), .Y(n_811) );
NAND2x1_ASAP7_75t_L g812 ( .A(n_749), .B(n_650), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_716), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_799), .B(n_724), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_786), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_793), .B(n_713), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_779), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_780), .Y(n_818) );
INVx1_ASAP7_75t_SL g819 ( .A(n_811), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_797), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_781), .Y(n_821) );
NAND2x1_ASAP7_75t_L g822 ( .A(n_793), .B(n_749), .Y(n_822) );
INVx1_ASAP7_75t_SL g823 ( .A(n_806), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_773), .A2(n_759), .B1(n_761), .B2(n_731), .Y(n_824) );
OR2x2_ASAP7_75t_L g825 ( .A(n_799), .B(n_724), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_791), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_782), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_810), .B(n_713), .Y(n_828) );
INVxp67_ASAP7_75t_L g829 ( .A(n_802), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_813), .Y(n_830) );
INVx2_ASAP7_75t_SL g831 ( .A(n_788), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_792), .Y(n_832) );
AOI32xp33_ASAP7_75t_L g833 ( .A1(n_794), .A2(n_735), .A3(n_737), .B1(n_767), .B2(n_768), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_787), .B(n_770), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_805), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_803), .Y(n_836) );
BUFx2_ASAP7_75t_SL g837 ( .A(n_819), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_823), .A2(n_776), .B1(n_775), .B2(n_778), .Y(n_838) );
NAND3x2_ASAP7_75t_L g839 ( .A(n_814), .B(n_776), .C(n_795), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_831), .A2(n_784), .B1(n_796), .B2(n_808), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_835), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_817), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_829), .B(n_796), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_816), .A2(n_783), .B1(n_767), .B2(n_798), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g845 ( .A1(n_824), .A2(n_790), .B1(n_800), .B2(n_812), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_826), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_815), .B(n_800), .Y(n_847) );
AND2x4_ASAP7_75t_SL g848 ( .A(n_816), .B(n_827), .Y(n_848) );
OAI211xp5_ASAP7_75t_L g849 ( .A1(n_833), .A2(n_768), .B(n_752), .C(n_754), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_825), .B(n_807), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_820), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_834), .B(n_809), .Y(n_852) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_849), .B(n_818), .C(n_821), .Y(n_853) );
OAI211xp5_ASAP7_75t_L g854 ( .A1(n_839), .A2(n_822), .B(n_828), .C(n_764), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_850), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_847), .A2(n_830), .B1(n_836), .B2(n_832), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_841), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_842), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_843), .B(n_830), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g860 ( .A1(n_845), .A2(n_789), .B1(n_777), .B2(n_836), .Y(n_860) );
OAI321xp33_ASAP7_75t_L g861 ( .A1(n_840), .A2(n_809), .A3(n_777), .B1(n_801), .B2(n_804), .C(n_638), .Y(n_861) );
OAI321xp33_ASAP7_75t_L g862 ( .A1(n_852), .A2(n_769), .A3(n_748), .B1(n_742), .B2(n_785), .C(n_774), .Y(n_862) );
INVxp67_ASAP7_75t_SL g863 ( .A(n_846), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_854), .A2(n_838), .B1(n_844), .B2(n_837), .C(n_851), .Y(n_864) );
NOR2xp67_ASAP7_75t_SL g865 ( .A(n_862), .B(n_672), .Y(n_865) );
OAI21xp33_ASAP7_75t_SL g866 ( .A1(n_863), .A2(n_848), .B(n_702), .Y(n_866) );
AOI222xp33_ASAP7_75t_L g867 ( .A1(n_853), .A2(n_755), .B1(n_750), .B2(n_679), .C1(n_725), .C2(n_745), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_860), .A2(n_678), .B1(n_743), .B2(n_756), .C(n_733), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_855), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_857), .B(n_757), .Y(n_870) );
NAND4xp25_ASAP7_75t_L g871 ( .A(n_864), .B(n_856), .C(n_861), .D(n_859), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_869), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_SL g873 ( .A1(n_865), .A2(n_677), .B(n_858), .C(n_734), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_866), .B(n_743), .Y(n_874) );
OAI211xp5_ASAP7_75t_SL g875 ( .A1(n_867), .A2(n_698), .B(n_667), .C(n_756), .Y(n_875) );
NOR2x1_ASAP7_75t_L g876 ( .A(n_871), .B(n_874), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g877 ( .A(n_873), .B(n_868), .C(n_870), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_872), .B(n_757), .Y(n_878) );
OAI21xp33_ASAP7_75t_L g879 ( .A1(n_876), .A2(n_875), .B(n_733), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_877), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_878), .B(n_771), .Y(n_881) );
NOR3xp33_ASAP7_75t_L g882 ( .A(n_880), .B(n_879), .C(n_881), .Y(n_882) );
AND3x2_ASAP7_75t_L g883 ( .A(n_880), .B(n_703), .C(n_771), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_882), .A2(n_763), .B1(n_701), .B2(n_766), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_883), .Y(n_885) );
AND2x2_ASAP7_75t_SL g886 ( .A(n_885), .B(n_697), .Y(n_886) );
OAI22xp5_ASAP7_75t_SL g887 ( .A1(n_884), .A2(n_680), .B1(n_765), .B2(n_214), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_886), .A2(n_216), .B1(n_218), .B2(n_224), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g889 ( .A1(n_887), .A2(n_225), .B1(n_226), .B2(n_229), .C(n_230), .Y(n_889) );
AOI222xp33_ASAP7_75t_L g890 ( .A1(n_888), .A2(n_231), .B1(n_232), .B2(n_233), .C1(n_234), .C2(n_235), .Y(n_890) );
OAI21xp5_ASAP7_75t_L g891 ( .A1(n_889), .A2(n_236), .B(n_237), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_891), .A2(n_239), .B(n_240), .Y(n_892) );
OR2x6_ASAP7_75t_L g893 ( .A(n_892), .B(n_890), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_893), .A2(n_241), .B1(n_242), .B2(n_243), .Y(n_894) );
endmodule