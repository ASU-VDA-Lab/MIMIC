module fake_netlist_6_977_n_2083 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2083);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2083;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

BUFx8_ASAP7_75t_SL g198 ( 
.A(n_45),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_76),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_64),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_38),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_72),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_13),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_21),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_85),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_54),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_190),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_81),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_167),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_20),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_129),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_82),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_42),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_93),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_15),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_71),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_54),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_150),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_113),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_84),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_66),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_182),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_166),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_7),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_98),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_77),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_67),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_67),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_59),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_30),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_0),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_6),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_128),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_71),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_165),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_138),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_106),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_41),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_80),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_4),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_108),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_88),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_76),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_33),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_62),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_75),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_179),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_30),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_53),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_104),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_12),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_91),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_66),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_74),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_153),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_43),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_134),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_97),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_68),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_27),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_103),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_131),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_162),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_39),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_95),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_116),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_65),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_65),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_52),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_169),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_122),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_189),
.Y(n_313)
);

BUFx4f_ASAP7_75t_SL g314 ( 
.A(n_142),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_40),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_173),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_74),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_87),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_124),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_33),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_39),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_14),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_25),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_92),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_114),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_68),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_105),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_61),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_73),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_154),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_161),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_29),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_191),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_24),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_29),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_25),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_137),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_70),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_37),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_118),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_14),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_117),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_130),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_11),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_86),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_8),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_16),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_141),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_170),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_41),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_1),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_8),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_183),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_52),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_44),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_90),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_140),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_28),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_24),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_16),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_96),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_27),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_72),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_10),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_58),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_111),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_53),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_139),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_23),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_56),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_11),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_22),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_175),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_158),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_168),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_143),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_23),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_18),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_17),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_44),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_136),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_156),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_59),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_127),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_4),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_47),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_180),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_198),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_208),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_259),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_213),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_215),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_220),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_219),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_244),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_357),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_226),
.B(n_0),
.Y(n_408)
);

INVxp33_ASAP7_75t_SL g409 ( 
.A(n_348),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_300),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_221),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_222),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_224),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_267),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_227),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_211),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_228),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_241),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_348),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_268),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_255),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_255),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_1),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_260),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_197),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_242),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_260),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_270),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_262),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_269),
.B(n_2),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_262),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_315),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_269),
.B(n_2),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_245),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_249),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_233),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_257),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_307),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_259),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_251),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_256),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_264),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_340),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_343),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_312),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_271),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_343),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_201),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_273),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_201),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_274),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_314),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_270),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_275),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_302),
.B(n_3),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_315),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_282),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_288),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_301),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_313),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_199),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_342),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_342),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_259),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_233),
.B(n_5),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_317),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_319),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_325),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_237),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_206),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_326),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_329),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_302),
.B(n_5),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_302),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_332),
.Y(n_484)
);

BUFx6f_ASAP7_75t_SL g485 ( 
.A(n_378),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_374),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_315),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_302),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_333),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_237),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_341),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_410),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_393),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_344),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_460),
.B(n_300),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_424),
.B(n_399),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_346),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_347),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_202),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_396),
.B(n_223),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_465),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_403),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_406),
.B(n_408),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_481),
.A2(n_239),
.B(n_223),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_405),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_404),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_473),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_415),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_407),
.A2(n_266),
.B(n_252),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_491),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_475),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_490),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_450),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_492),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_450),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_470),
.B(n_202),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_239),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_398),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

CKINVDCx8_ASAP7_75t_R g540 ( 
.A(n_429),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_413),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_421),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_442),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_413),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_400),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_401),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_452),
.B(n_240),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_425),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_402),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_411),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_406),
.B(n_370),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_471),
.A2(n_263),
.B(n_240),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_452),
.B(n_203),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_412),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_428),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_428),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_431),
.B(n_350),
.Y(n_569)
);

OA21x2_ASAP7_75t_L g570 ( 
.A1(n_432),
.A2(n_266),
.B(n_252),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_449),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_435),
.B(n_370),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_414),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_420),
.B1(n_468),
.B2(n_429),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_572),
.A2(n_467),
.B1(n_426),
.B2(n_409),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_502),
.B(n_416),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_502),
.B(n_489),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_569),
.B(n_300),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_500),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_505),
.B(n_463),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_418),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_419),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_R g585 ( 
.A(n_544),
.B(n_395),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_536),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_536),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_471),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_532),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_539),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_532),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_496),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_499),
.B(n_300),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_499),
.B(n_427),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_503),
.B(n_436),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

BUFx6f_ASAP7_75t_SL g600 ( 
.A(n_537),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_532),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_496),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_532),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_501),
.B(n_263),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_497),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_513),
.B(n_455),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_513),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_563),
.B(n_489),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_500),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_503),
.B(n_438),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_501),
.A2(n_485),
.B1(n_458),
.B2(n_290),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_501),
.A2(n_477),
.B1(n_441),
.B2(n_469),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_505),
.B(n_444),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_509),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_496),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_536),
.B(n_445),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_501),
.A2(n_562),
.B1(n_537),
.B2(n_556),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_496),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_510),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_539),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_537),
.B(n_294),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_563),
.B(n_463),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_510),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_506),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_563),
.B(n_472),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_506),
.B(n_446),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_506),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_546),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_506),
.B(n_451),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_515),
.A2(n_290),
.B1(n_297),
.B2(n_278),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_524),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_524),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_524),
.B(n_294),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_537),
.B(n_303),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_537),
.B(n_303),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_562),
.B(n_537),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

INVx4_ASAP7_75t_SL g646 ( 
.A(n_510),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_454),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_556),
.B(n_300),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_456),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_535),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_540),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_494),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_497),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_561),
.A2(n_462),
.B1(n_464),
.B2(n_459),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_511),
.B(n_466),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_556),
.B(n_300),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_512),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_512),
.B(n_474),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_514),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_538),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_556),
.B(n_392),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_392),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_497),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_510),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_561),
.B(n_468),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_509),
.B(n_457),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_514),
.B(n_478),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_562),
.B(n_232),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_556),
.B(n_392),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_508),
.B(n_472),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_553),
.B(n_392),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_508),
.B(n_479),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_519),
.B(n_480),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_518),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_546),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_510),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_520),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_520),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_510),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_497),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_570),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_523),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_570),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_544),
.B(n_469),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_508),
.B(n_479),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_553),
.B(n_484),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_546),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_498),
.B(n_541),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_498),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_541),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_565),
.B(n_486),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_565),
.B(n_567),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_508),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_498),
.B(n_482),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_508),
.A2(n_485),
.B1(n_278),
.B2(n_390),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_565),
.B(n_482),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_517),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_541),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_541),
.B(n_529),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_555),
.B(n_485),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_497),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_518),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_508),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_493),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_541),
.Y(n_716)
);

NOR2x1p5_ASAP7_75t_L g717 ( 
.A(n_555),
.B(n_486),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_529),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_493),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_566),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_517),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_SL g722 ( 
.A(n_559),
.B(n_485),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_529),
.B(n_366),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_517),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_542),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_672),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_589),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_573),
.B(n_559),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_672),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_642),
.B(n_560),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_721),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_597),
.B(n_560),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_693),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_606),
.A2(n_305),
.B1(n_308),
.B2(n_297),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_642),
.B(n_564),
.Y(n_735)
);

AOI21x1_ASAP7_75t_L g736 ( 
.A1(n_606),
.A2(n_516),
.B(n_534),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_574),
.A2(n_258),
.B1(n_334),
.B2(n_284),
.C(n_316),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_588),
.A2(n_564),
.B1(n_373),
.B2(n_380),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_614),
.A2(n_540),
.B1(n_203),
.B2(n_207),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_598),
.B(n_534),
.Y(n_740)
);

AND3x1_ASAP7_75t_L g741 ( 
.A(n_575),
.B(n_308),
.C(n_305),
.Y(n_741)
);

O2A1O1Ixp5_ASAP7_75t_L g742 ( 
.A1(n_662),
.A2(n_205),
.B(n_209),
.C(n_207),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_576),
.B(n_540),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_589),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_721),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_677),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_642),
.B(n_392),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_588),
.A2(n_381),
.B1(n_386),
.B2(n_371),
.Y(n_748)
);

NOR2x2_ASAP7_75t_L g749 ( 
.A(n_635),
.B(n_204),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_677),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_613),
.B(n_534),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_586),
.B(n_521),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_586),
.B(n_587),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_587),
.B(n_392),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_638),
.A2(n_697),
.B1(n_607),
.B2(n_632),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_583),
.B(n_528),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_584),
.B(n_528),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_589),
.B(n_528),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_714),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_620),
.B(n_693),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_702),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_SL g762 ( 
.A(n_582),
.B(n_521),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_668),
.B(n_544),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_702),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_668),
.B(n_526),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_707),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_662),
.B(n_315),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_638),
.B(n_528),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_703),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_704),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_721),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_701),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_647),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_662),
.B(n_690),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_649),
.B(n_200),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_577),
.A2(n_387),
.B1(n_389),
.B2(n_209),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_690),
.B(n_531),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_701),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_713),
.B(n_526),
.Y(n_780)
);

AO22x1_ASAP7_75t_L g781 ( 
.A1(n_616),
.A2(n_331),
.B1(n_337),
.B2(n_345),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_690),
.B(n_531),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_707),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_656),
.B(n_210),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_708),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_610),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_674),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_690),
.B(n_315),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_607),
.A2(n_390),
.B1(n_364),
.B2(n_345),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_692),
.B(n_531),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_674),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_678),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_678),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_678),
.Y(n_796)
);

OAI221xp5_ASAP7_75t_L g797 ( 
.A1(n_706),
.A2(n_439),
.B1(n_476),
.B2(n_364),
.C(n_337),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_581),
.B(n_542),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_692),
.B(n_531),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_692),
.B(n_533),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_692),
.B(n_533),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_632),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_694),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_621),
.B(n_315),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_577),
.A2(n_516),
.B(n_322),
.C(n_330),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_660),
.B(n_212),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_670),
.B(n_217),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_636),
.A2(n_330),
.B1(n_323),
.B2(n_322),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_611),
.B(n_533),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_611),
.B(n_533),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_626),
.B(n_566),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_704),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_651),
.B(n_323),
.Y(n_814)
);

NOR2x2_ASAP7_75t_L g815 ( 
.A(n_635),
.B(n_218),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_679),
.B(n_225),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_714),
.B(n_671),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_626),
.B(n_566),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_643),
.B(n_644),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_591),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_645),
.B(n_566),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_591),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_694),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_650),
.B(n_629),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_SL g825 ( 
.A(n_582),
.B(n_527),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_581),
.A2(n_361),
.B1(n_214),
.B2(n_216),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_SL g827 ( 
.A1(n_637),
.A2(n_331),
.B1(n_567),
.B2(n_568),
.C(n_549),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_580),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_629),
.B(n_566),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_639),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_714),
.B(n_671),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_708),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_610),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_635),
.A2(n_516),
.B1(n_354),
.B2(n_286),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_629),
.B(n_205),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_601),
.B(n_214),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_L g837 ( 
.A(n_630),
.B(n_315),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_675),
.A2(n_549),
.B(n_568),
.C(n_550),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_592),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_599),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_714),
.B(n_315),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_581),
.A2(n_361),
.B1(n_230),
.B2(n_231),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_601),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_605),
.B(n_725),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_605),
.B(n_216),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_652),
.B(n_230),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_657),
.B(n_231),
.Y(n_847)
);

NAND2x1_ASAP7_75t_L g848 ( 
.A(n_700),
.B(n_493),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_675),
.B(n_229),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_659),
.B(n_234),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_724),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_724),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_661),
.B(n_234),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_635),
.A2(n_250),
.B1(n_276),
.B2(n_362),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_682),
.B(n_250),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_695),
.B(n_530),
.C(n_527),
.Y(n_856)
);

AOI221xp5_ASAP7_75t_L g857 ( 
.A1(n_722),
.A2(n_289),
.B1(n_285),
.B2(n_247),
.C(n_238),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_717),
.A2(n_276),
.B1(n_335),
.B2(n_349),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_612),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_634),
.B(n_235),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_600),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_699),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_684),
.B(n_685),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_579),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_686),
.B(n_286),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_654),
.B(n_236),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_604),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_625),
.A2(n_550),
.B(n_552),
.C(n_558),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_628),
.A2(n_354),
.B1(n_293),
.B2(n_306),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_579),
.Y(n_870)
);

AOI221xp5_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_309),
.B1(n_365),
.B2(n_368),
.C(n_382),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_582),
.B(n_663),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_691),
.B(n_291),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_669),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_680),
.Y(n_875)
);

INVx8_ASAP7_75t_L g876 ( 
.A(n_600),
.Y(n_876)
);

BUFx5_ASAP7_75t_L g877 ( 
.A(n_658),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_631),
.B(n_723),
.Y(n_878)
);

BUFx12f_ASAP7_75t_L g879 ( 
.A(n_663),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_608),
.A2(n_495),
.B(n_493),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_653),
.A2(n_507),
.B(n_495),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_666),
.B(n_291),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_663),
.B(n_530),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_711),
.B(n_246),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_625),
.B(n_293),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_688),
.B(n_306),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_705),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_700),
.B(n_311),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_590),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_700),
.B(n_311),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_720),
.B(n_320),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_600),
.A2(n_320),
.B1(n_353),
.B2(n_358),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_709),
.B(n_327),
.Y(n_893)
);

BUFx12f_ASAP7_75t_L g894 ( 
.A(n_618),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_609),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_680),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_720),
.B(n_248),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_752),
.B(n_618),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_786),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_874),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_887),
.B(n_720),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_733),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_755),
.B(n_709),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_743),
.A2(n_718),
.B1(n_578),
.B2(n_595),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_763),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_744),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_814),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_SL g908 ( 
.A(n_755),
.B(n_522),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_770),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_727),
.B(n_552),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_770),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_774),
.B(n_740),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_SL g913 ( 
.A1(n_860),
.A2(n_578),
.B(n_595),
.C(n_619),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_736),
.A2(n_594),
.B(n_593),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_867),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_790),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_751),
.B(n_709),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_833),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_790),
.B(n_716),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_860),
.B(n_716),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_894),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_726),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_727),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_875),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_726),
.B(n_716),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_728),
.B(n_609),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_798),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_776),
.B(n_784),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_879),
.B(n_872),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_820),
.B(n_554),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_798),
.Y(n_931)
);

AO22x1_ASAP7_75t_L g932 ( 
.A1(n_866),
.A2(n_363),
.B1(n_296),
.B2(n_295),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_762),
.B(n_522),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_729),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_SL g935 ( 
.A(n_857),
.B(n_585),
.C(n_254),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_896),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_760),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_SL g938 ( 
.A1(n_866),
.A2(n_571),
.B1(n_545),
.B2(n_543),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_729),
.A2(n_746),
.B1(n_802),
.B2(n_750),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_780),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_814),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_SL g942 ( 
.A(n_871),
.B(n_545),
.C(n_543),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_728),
.B(n_764),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_896),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_867),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_867),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_746),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_876),
.Y(n_949)
);

AOI22x1_ASAP7_75t_L g950 ( 
.A1(n_830),
.A2(n_619),
.B1(n_603),
.B2(n_594),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_787),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_820),
.B(n_554),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_776),
.B(n_571),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_844),
.B(n_557),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_883),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_814),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_876),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_844),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_784),
.B(n_593),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_732),
.B(n_383),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_807),
.B(n_593),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_789),
.B(n_793),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_805),
.A2(n_849),
.B1(n_739),
.B2(n_791),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_807),
.B(n_594),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_750),
.A2(n_718),
.B1(n_640),
.B2(n_641),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_743),
.B(n_384),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_794),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_761),
.Y(n_968)
);

OR2x2_ASAP7_75t_SL g969 ( 
.A(n_749),
.B(n_327),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_802),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_808),
.B(n_816),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_808),
.A2(n_718),
.B1(n_641),
.B2(n_640),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_816),
.B(n_603),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_795),
.B(n_557),
.Y(n_974)
);

NOR3xp33_ASAP7_75t_SL g975 ( 
.A(n_737),
.B(n_261),
.C(n_253),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_867),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_832),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_813),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_895),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_813),
.B(n_712),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_756),
.B(n_603),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_757),
.B(n_619),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_796),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_738),
.B(n_648),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_741),
.Y(n_986)
);

OR2x6_ASAP7_75t_SL g987 ( 
.A(n_824),
.B(n_265),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_765),
.B(n_206),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_849),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_813),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_825),
.B(n_272),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_884),
.B(n_596),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_753),
.B(n_698),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_767),
.B(n_648),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_753),
.A2(n_673),
.B(n_710),
.C(n_335),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_783),
.B(n_590),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_851),
.Y(n_998)
);

CKINVDCx11_ASAP7_75t_R g999 ( 
.A(n_861),
.Y(n_999)
);

AND3x1_ASAP7_75t_SL g1000 ( 
.A(n_766),
.B(n_353),
.C(n_349),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_852),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_830),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_803),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_897),
.B(n_615),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_804),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_852),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_823),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_862),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_771),
.B(n_277),
.Y(n_1009)
);

INVxp33_ASAP7_75t_L g1010 ( 
.A(n_884),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_897),
.B(n_878),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_862),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_730),
.B(n_596),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_748),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_822),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_828),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_771),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_861),
.B(n_279),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_SL g1019 ( 
.A(n_730),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_839),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_870),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_805),
.A2(n_673),
.B1(n_664),
.B2(n_658),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_813),
.B(n_712),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_840),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_735),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_859),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_819),
.B(n_615),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_735),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_822),
.B(n_358),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_829),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_822),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_837),
.B(n_280),
.Y(n_1032)
);

AND3x1_ASAP7_75t_SL g1033 ( 
.A(n_797),
.B(n_379),
.C(n_362),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_870),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_863),
.B(n_624),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_758),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_778),
.B(n_624),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_769),
.A2(n_379),
.B1(n_712),
.B2(n_627),
.Y(n_1039)
);

INVx4_ASAP7_75t_SL g1040 ( 
.A(n_843),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_856),
.B(n_206),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_782),
.B(n_633),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_775),
.B(n_596),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_843),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_810),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_877),
.B(n_712),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_759),
.B(n_602),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_843),
.B(n_558),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_858),
.B(n_206),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_843),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_815),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_775),
.A2(n_835),
.B1(n_818),
.B2(n_812),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_889),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_811),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_889),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_821),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_885),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_759),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_868),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_773),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_779),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_848),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_785),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_792),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_799),
.B(n_800),
.Y(n_1065)
);

AO21x2_ASAP7_75t_L g1066 ( 
.A1(n_817),
.A2(n_633),
.B(n_681),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_885),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_885),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_836),
.B(n_845),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_864),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_801),
.Y(n_1071)
);

AO21x2_ASAP7_75t_L g1072 ( 
.A1(n_817),
.A2(n_831),
.B(n_768),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_869),
.B(n_281),
.C(n_283),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_877),
.B(n_292),
.Y(n_1074)
);

CKINVDCx14_ASAP7_75t_R g1075 ( 
.A(n_854),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_731),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_745),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_791),
.B(n_734),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_734),
.B(n_655),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_772),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_747),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_846),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_781),
.B(n_567),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_847),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_850),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_853),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_831),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_777),
.B(n_602),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_747),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_877),
.B(n_298),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_855),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_962),
.B(n_768),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_928),
.A2(n_788),
.B(n_742),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_915),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1065),
.A2(n_788),
.B(n_622),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_914),
.A2(n_881),
.B(n_880),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_914),
.A2(n_841),
.B(n_888),
.Y(n_1097)
);

NAND2x1_ASAP7_75t_L g1098 ( 
.A(n_1058),
.B(n_604),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_950),
.A2(n_841),
.B(n_890),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_939),
.A2(n_834),
.B(n_754),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_971),
.B(n_877),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_920),
.A2(n_622),
.B(n_602),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1038),
.A2(n_893),
.B(n_754),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_SL g1104 ( 
.A(n_1058),
.B(n_891),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_962),
.B(n_865),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1011),
.A2(n_891),
.B(n_834),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1064),
.A2(n_622),
.B(n_667),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_963),
.A2(n_809),
.B1(n_886),
.B2(n_882),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_911),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_903),
.A2(n_667),
.B(n_627),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1042),
.A2(n_838),
.B(n_873),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_903),
.A2(n_1052),
.B(n_1081),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1078),
.A2(n_809),
.B(n_806),
.C(n_826),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_917),
.A2(n_667),
.B(n_687),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1046),
.A2(n_681),
.B(n_655),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_912),
.B(n_842),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1010),
.B(n_892),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_966),
.A2(n_806),
.B(n_827),
.C(n_375),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_696),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1002),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_905),
.B(n_937),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1045),
.B(n_1054),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1010),
.B(n_877),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1058),
.B(n_604),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_960),
.A2(n_372),
.B(n_367),
.C(n_360),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_901),
.A2(n_627),
.B(n_604),
.Y(n_1126)
);

NOR2xp67_ASAP7_75t_SL g1127 ( 
.A(n_1067),
.B(n_957),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_944),
.B(n_696),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_911),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_916),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1084),
.B(n_715),
.Y(n_1131)
);

BUFx10_ASAP7_75t_L g1132 ( 
.A(n_900),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1081),
.A2(n_1089),
.B(n_1043),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_915),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1089),
.A2(n_623),
.B1(n_627),
.B2(n_676),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1047),
.A2(n_623),
.B(n_676),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_972),
.A2(n_623),
.B1(n_689),
.B2(n_687),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1046),
.A2(n_925),
.B(n_981),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1087),
.B(n_877),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_926),
.B(n_299),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_935),
.A2(n_388),
.B(n_304),
.C(n_310),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_925),
.A2(n_495),
.B(n_507),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1059),
.A2(n_432),
.A3(n_434),
.B(n_437),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1049),
.A2(n_391),
.B(n_318),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_495),
.B(n_507),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1091),
.B(n_1082),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_434),
.A3(n_437),
.B(n_440),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_993),
.A2(n_904),
.B1(n_1088),
.B2(n_1028),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1085),
.B(n_715),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_959),
.A2(n_507),
.B(n_551),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1047),
.A2(n_964),
.B(n_961),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_981),
.A2(n_547),
.B(n_548),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_973),
.A2(n_676),
.B(n_623),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_965),
.A2(n_440),
.A3(n_447),
.B(n_547),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1023),
.A2(n_547),
.B(n_548),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1023),
.A2(n_547),
.B(n_548),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_898),
.B(n_243),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_977),
.A2(n_548),
.B(n_551),
.Y(n_1158)
);

BUFx2_ASAP7_75t_R g1159 ( 
.A(n_936),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_982),
.A2(n_551),
.B(n_447),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1037),
.A2(n_658),
.B(n_664),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1013),
.A2(n_551),
.A3(n_658),
.B(n_664),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1030),
.A2(n_658),
.B(n_664),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_953),
.B(n_243),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_919),
.A2(n_676),
.B(n_689),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_983),
.A2(n_683),
.B(n_689),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_977),
.A2(n_646),
.B(n_719),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_988),
.B(n_243),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_916),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_SL g1170 ( 
.A(n_915),
.B(n_683),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1002),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_936),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1087),
.B(n_1067),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1025),
.A2(n_689),
.B1(n_687),
.B2(n_683),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1025),
.A2(n_687),
.B1(n_683),
.B2(n_715),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_994),
.A2(n_715),
.B(n_719),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_978),
.A2(n_646),
.B(n_719),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1086),
.B(n_719),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1027),
.A2(n_719),
.B(n_646),
.Y(n_1179)
);

AOI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1014),
.A2(n_321),
.B(n_324),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_909),
.B(n_665),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_978),
.A2(n_646),
.B(n_664),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_908),
.A2(n_378),
.B(n_10),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_975),
.A2(n_355),
.B(n_377),
.C(n_336),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1036),
.A2(n_665),
.B(n_664),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1008),
.A2(n_665),
.B(n_658),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_995),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_L g1188 ( 
.A1(n_913),
.A2(n_665),
.B(n_378),
.C(n_287),
.Y(n_1188)
);

INVx5_ASAP7_75t_L g1189 ( 
.A(n_915),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_946),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_995),
.B(n_665),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1016),
.B(n_665),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_985),
.A2(n_385),
.B(n_338),
.C(n_376),
.Y(n_1193)
);

NOR2x1_ASAP7_75t_SL g1194 ( 
.A(n_946),
.B(n_89),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_913),
.A2(n_1071),
.B(n_934),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_976),
.A2(n_83),
.B(n_195),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1071),
.A2(n_78),
.B(n_101),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1079),
.A2(n_359),
.B(n_356),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_968),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1071),
.A2(n_155),
.B(n_110),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_922),
.A2(n_352),
.B(n_351),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_991),
.A2(n_148),
.B(n_193),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1040),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_991),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1071),
.A2(n_144),
.B(n_192),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1072),
.A2(n_378),
.B(n_187),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_998),
.A2(n_186),
.B(n_184),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_979),
.B(n_181),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1020),
.B(n_287),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1055),
.A2(n_287),
.B(n_243),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_922),
.A2(n_172),
.B(n_171),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_940),
.B(n_955),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_998),
.A2(n_160),
.B(n_135),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1001),
.A2(n_132),
.B(n_126),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1001),
.A2(n_123),
.B(n_119),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1006),
.A2(n_115),
.B(n_112),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_955),
.B(n_287),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_934),
.A2(n_109),
.B(n_12),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_962),
.B(n_9),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1072),
.A2(n_9),
.B(n_17),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1024),
.B(n_18),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1026),
.B(n_19),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_908),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_948),
.A2(n_26),
.B(n_31),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_906),
.B(n_26),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1012),
.A2(n_31),
.A3(n_32),
.B(n_34),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_948),
.A2(n_996),
.B(n_970),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_958),
.B(n_34),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_970),
.A2(n_36),
.B(n_37),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1006),
.A2(n_36),
.B(n_43),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_976),
.A2(n_73),
.B(n_48),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1087),
.B(n_46),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_957),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1069),
.A2(n_1066),
.B(n_997),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1021),
.A2(n_46),
.A3(n_48),
.B(n_49),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1021),
.A2(n_49),
.A3(n_50),
.B(n_51),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_951),
.B(n_50),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1087),
.B(n_55),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_946),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_902),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1067),
.B(n_55),
.Y(n_1241)
);

O2A1O1Ixp5_ASAP7_75t_L g1242 ( 
.A1(n_1017),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1028),
.B(n_57),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_954),
.B(n_1041),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1035),
.A2(n_60),
.B(n_62),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1035),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1053),
.A2(n_60),
.B(n_63),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_976),
.A2(n_63),
.B(n_69),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1040),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1067),
.A2(n_69),
.B1(n_70),
.B2(n_1014),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1031),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1053),
.A2(n_970),
.B(n_1077),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_979),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_979),
.B(n_1031),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1017),
.A2(n_1076),
.B(n_1077),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_990),
.A2(n_1017),
.B(n_947),
.Y(n_1256)
);

AOI211xp5_ASAP7_75t_L g1257 ( 
.A1(n_1180),
.A2(n_942),
.B(n_932),
.C(n_1051),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1140),
.A2(n_938),
.B1(n_980),
.B2(n_1019),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1140),
.B(n_900),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1204),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1246),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1246),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1109),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1129),
.Y(n_1264)
);

NOR2xp67_ASAP7_75t_L g1265 ( 
.A(n_1240),
.B(n_929),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1187),
.B(n_910),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1118),
.A2(n_1070),
.B(n_1063),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1252),
.A2(n_1076),
.B(n_1070),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1148),
.A2(n_1067),
.B1(n_1075),
.B2(n_943),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1255),
.A2(n_1050),
.B(n_1080),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1172),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1118),
.A2(n_1060),
.B(n_1061),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1117),
.A2(n_1075),
.B1(n_931),
.B2(n_927),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1130),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1169),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1240),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1113),
.A2(n_923),
.B(n_1083),
.C(n_990),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_SL g1278 ( 
.A1(n_1113),
.A2(n_1003),
.B(n_984),
.C(n_1007),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1233),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1146),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1255),
.A2(n_1050),
.B(n_1005),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1188),
.A2(n_967),
.B(n_1022),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1108),
.A2(n_986),
.A3(n_1033),
.B(n_1000),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1212),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1173),
.B(n_1029),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1120),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1120),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1125),
.A2(n_969),
.B1(n_918),
.B2(n_899),
.C(n_924),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1183),
.A2(n_1066),
.A3(n_987),
.B(n_1029),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1145),
.A2(n_1050),
.B(n_1057),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1244),
.A2(n_1117),
.B1(n_980),
.B2(n_1217),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1243),
.A2(n_933),
.B1(n_992),
.B2(n_945),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1096),
.A2(n_1150),
.B(n_1097),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1068),
.B(n_1040),
.Y(n_1294)
);

BUFx2_ASAP7_75t_R g1295 ( 
.A(n_1233),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1138),
.A2(n_907),
.B(n_956),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1199),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1099),
.A2(n_941),
.B(n_1029),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1122),
.B(n_910),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1167),
.A2(n_1029),
.B(n_1062),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1177),
.A2(n_1062),
.B(n_947),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1213),
.A2(n_1062),
.B(n_947),
.Y(n_1302)
);

AOI22x1_ASAP7_75t_L g1303 ( 
.A1(n_1106),
.A2(n_1048),
.B1(n_910),
.B2(n_974),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1214),
.A2(n_1062),
.B(n_947),
.Y(n_1304)
);

O2A1O1Ixp5_ASAP7_75t_L g1305 ( 
.A1(n_1188),
.A2(n_1048),
.B(n_974),
.C(n_952),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1171),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1151),
.A2(n_987),
.A3(n_1069),
.B(n_1073),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1171),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1112),
.A2(n_974),
.B(n_1048),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_1253),
.B(n_1044),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1115),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1215),
.A2(n_946),
.B(n_1044),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1121),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1100),
.A2(n_930),
.B(n_952),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1152),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1173),
.B(n_1139),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1116),
.B(n_930),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1172),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1160),
.A2(n_930),
.B(n_952),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1100),
.A2(n_954),
.B(n_1032),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1092),
.A2(n_949),
.B1(n_943),
.B2(n_1015),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1143),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1105),
.B(n_954),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1216),
.A2(n_1044),
.B(n_1031),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1155),
.A2(n_1044),
.B(n_1031),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1143),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1143),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1203),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1143),
.Y(n_1329)
);

BUFx4f_ASAP7_75t_L g1330 ( 
.A(n_1203),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1128),
.B(n_1009),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1178),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1144),
.B(n_945),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1125),
.A2(n_1223),
.B(n_1250),
.C(n_1193),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1131),
.B(n_1105),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1156),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1093),
.A2(n_1133),
.B(n_1101),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1153),
.A2(n_1207),
.B(n_1202),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1105),
.B(n_1034),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1202),
.A2(n_1034),
.B(n_1015),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1092),
.B(n_1219),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1092),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1207),
.A2(n_943),
.B(n_949),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1111),
.A2(n_1032),
.B(n_1090),
.Y(n_1344)
);

BUFx2_ASAP7_75t_SL g1345 ( 
.A(n_1189),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1132),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1103),
.A2(n_949),
.B(n_1074),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1142),
.A2(n_1090),
.B(n_1074),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1119),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1203),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1209),
.B(n_921),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1110),
.A2(n_1009),
.B(n_999),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1132),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1149),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1179),
.A2(n_999),
.B(n_1018),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1227),
.A2(n_1018),
.B(n_992),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1154),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1101),
.A2(n_933),
.B(n_921),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1154),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1154),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1166),
.A2(n_1102),
.B(n_1095),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1230),
.A2(n_1247),
.B(n_1245),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1253),
.B(n_1219),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1157),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_SL g1365 ( 
.A1(n_1141),
.A2(n_1223),
.B(n_1184),
.C(n_1193),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1219),
.B(n_1198),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1176),
.A2(n_1114),
.B(n_1182),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1228),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1154),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1181),
.Y(n_1370)
);

AOI21xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1243),
.A2(n_1164),
.B(n_1168),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1139),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1192),
.Y(n_1373)
);

BUFx8_ASAP7_75t_SL g1374 ( 
.A(n_1159),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1189),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1189),
.B(n_1239),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1094),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_R g1378 ( 
.A(n_1094),
.B(n_1134),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1189),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1126),
.A2(n_1165),
.B(n_1137),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1136),
.A2(n_1107),
.B(n_1135),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1123),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1229),
.A2(n_1184),
.B(n_1141),
.C(n_1237),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1254),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1256),
.A2(n_1186),
.B(n_1123),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1104),
.A2(n_1170),
.B(n_1191),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1211),
.A2(n_1197),
.B(n_1205),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1254),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1221),
.B(n_1222),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1200),
.A2(n_1185),
.B(n_1196),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1225),
.A2(n_1218),
.B(n_1201),
.C(n_1231),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_1190),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1241),
.A2(n_1232),
.B1(n_1238),
.B2(n_1248),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1241),
.A2(n_1238),
.B1(n_1232),
.B2(n_1224),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1242),
.A2(n_1161),
.B(n_1163),
.Y(n_1395)
);

AOI22x1_ASAP7_75t_L g1396 ( 
.A1(n_1208),
.A2(n_1124),
.B1(n_1249),
.B2(n_1251),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1190),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1190),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1175),
.A2(n_1174),
.B(n_1098),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1094),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1124),
.A2(n_1208),
.B(n_1242),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1194),
.B(n_1210),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1210),
.A2(n_1249),
.B(n_1234),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1210),
.A2(n_1127),
.B(n_1234),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1190),
.A2(n_1239),
.B1(n_1251),
.B2(n_1094),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1226),
.B(n_1236),
.Y(n_1406)
);

AOI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1206),
.A2(n_1147),
.B(n_1162),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1147),
.A2(n_1220),
.B(n_1206),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1239),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1134),
.B(n_1220),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1134),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1147),
.A2(n_1162),
.B(n_1235),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1226),
.A2(n_1235),
.B(n_1236),
.Y(n_1413)
);

AO22x2_ASAP7_75t_L g1414 ( 
.A1(n_1226),
.A2(n_1235),
.B1(n_1236),
.B2(n_1147),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1162),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1162),
.A2(n_1235),
.B(n_1236),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1226),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1195),
.A2(n_1252),
.B(n_1255),
.Y(n_1418)
);

NAND2x1_ASAP7_75t_L g1419 ( 
.A(n_1253),
.B(n_979),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1204),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1121),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1195),
.A2(n_1252),
.B(n_1255),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1195),
.A2(n_1252),
.B(n_1255),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1112),
.A2(n_1195),
.B(n_1194),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1285),
.B(n_1392),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1418),
.A2(n_1423),
.B(n_1422),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1258),
.A2(n_1291),
.B1(n_1280),
.B2(n_1317),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1259),
.A2(n_1366),
.B1(n_1273),
.B2(n_1393),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1330),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1333),
.A2(n_1364),
.B1(n_1257),
.B2(n_1366),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1313),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1354),
.B(n_1332),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1418),
.A2(n_1423),
.B(n_1422),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1394),
.A2(n_1331),
.B1(n_1269),
.B2(n_1341),
.Y(n_1434)
);

OR2x6_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_1392),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1330),
.Y(n_1436)
);

NAND2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1346),
.B(n_1328),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1276),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1324),
.A2(n_1312),
.B(n_1304),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1279),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1341),
.B(n_1368),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1279),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1323),
.A2(n_1292),
.B1(n_1342),
.B2(n_1389),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1285),
.B(n_1392),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1371),
.A2(n_1334),
.B1(n_1365),
.B2(n_1288),
.C(n_1421),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1284),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_SL g1447 ( 
.A(n_1346),
.B(n_1328),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1264),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1322),
.A2(n_1329),
.A3(n_1327),
.B(n_1326),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1264),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1383),
.B(n_1391),
.C(n_1351),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1277),
.A2(n_1278),
.B(n_1349),
.C(n_1424),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1323),
.A2(n_1299),
.B1(n_1266),
.B2(n_1265),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1266),
.A2(n_1303),
.B1(n_1356),
.B2(n_1342),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1303),
.A2(n_1356),
.B1(n_1358),
.B2(n_1354),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1271),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1274),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1358),
.A2(n_1382),
.B1(n_1337),
.B2(n_1332),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1274),
.Y(n_1460)
);

CKINVDCx8_ASAP7_75t_R g1461 ( 
.A(n_1345),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1353),
.Y(n_1462)
);

AOI222xp33_ASAP7_75t_L g1463 ( 
.A1(n_1335),
.A2(n_1318),
.B1(n_1382),
.B2(n_1339),
.C1(n_1275),
.C2(n_1373),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1363),
.A2(n_1330),
.B1(n_1285),
.B2(n_1353),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1424),
.A2(n_1361),
.B(n_1309),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1358),
.A2(n_1339),
.B1(n_1363),
.B2(n_1372),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1377),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1275),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1377),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1309),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1328),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1271),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1376),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1262),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1374),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1392),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1309),
.A2(n_1373),
.B1(n_1370),
.B2(n_1372),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1283),
.B(n_1307),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1350),
.B(n_1400),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1296),
.A2(n_1309),
.B1(n_1402),
.B2(n_1410),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1316),
.A2(n_1295),
.B1(n_1321),
.B2(n_1370),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1296),
.B(n_1384),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1283),
.B(n_1307),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1283),
.B(n_1307),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1283),
.B(n_1420),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1262),
.Y(n_1486)
);

NAND2xp33_ASAP7_75t_R g1487 ( 
.A(n_1378),
.B(n_1402),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1350),
.B(n_1400),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1376),
.B(n_1384),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1307),
.B(n_1308),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1316),
.A2(n_1355),
.B1(n_1417),
.B2(n_1352),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1376),
.B(n_1388),
.Y(n_1492)
);

AO31x2_ASAP7_75t_L g1493 ( 
.A1(n_1322),
.A2(n_1326),
.A3(n_1327),
.B(n_1329),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1411),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1388),
.B(n_1355),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1316),
.A2(n_1417),
.B1(n_1352),
.B2(n_1396),
.Y(n_1496)
);

NOR2x1_ASAP7_75t_SL g1497 ( 
.A(n_1345),
.B(n_1409),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1289),
.B(n_1286),
.Y(n_1498)
);

INVx4_ASAP7_75t_L g1499 ( 
.A(n_1409),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1397),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1409),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1305),
.A2(n_1387),
.B(n_1386),
.C(n_1390),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1396),
.A2(n_1417),
.B1(n_1395),
.B2(n_1406),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1397),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1417),
.A2(n_1406),
.B1(n_1395),
.B2(n_1369),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_1405),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1310),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_SL g1508 ( 
.A(n_1398),
.B(n_1375),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1398),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1387),
.A2(n_1379),
.B1(n_1375),
.B2(n_1272),
.Y(n_1510)
);

AOI21xp33_ASAP7_75t_L g1511 ( 
.A1(n_1395),
.A2(n_1314),
.B(n_1272),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1379),
.B(n_1260),
.Y(n_1512)
);

AND2x6_ASAP7_75t_L g1513 ( 
.A(n_1415),
.B(n_1417),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1287),
.B(n_1306),
.Y(n_1514)
);

NOR2x1p5_ASAP7_75t_L g1515 ( 
.A(n_1310),
.B(n_1419),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1419),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1314),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1287),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1413),
.A2(n_1414),
.B1(n_1369),
.B2(n_1360),
.C(n_1357),
.Y(n_1519)
);

OAI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1272),
.A2(n_1267),
.B1(n_1395),
.B2(n_1357),
.C(n_1360),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1261),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1289),
.B(n_1415),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1361),
.A2(n_1381),
.B(n_1344),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1314),
.A2(n_1272),
.B1(n_1267),
.B2(n_1320),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1298),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1359),
.A2(n_1320),
.B1(n_1267),
.B2(n_1282),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1359),
.A2(n_1320),
.B1(n_1267),
.B2(n_1282),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1414),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1289),
.B(n_1298),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1320),
.B(n_1399),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1416),
.B(n_1414),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1344),
.A2(n_1290),
.B1(n_1416),
.B2(n_1390),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1399),
.B(n_1416),
.Y(n_1533)
);

AO21x2_ASAP7_75t_L g1534 ( 
.A1(n_1404),
.A2(n_1338),
.B(n_1407),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1414),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1343),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1401),
.A2(n_1347),
.B1(n_1344),
.B2(n_1348),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1343),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1294),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1282),
.A2(n_1408),
.B1(n_1412),
.B2(n_1344),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1290),
.A2(n_1403),
.B(n_1385),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1362),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1401),
.B(n_1282),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1281),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1412),
.B(n_1403),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1408),
.B(n_1407),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1404),
.B(n_1319),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1408),
.A2(n_1380),
.B1(n_1348),
.B2(n_1347),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1311),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1408),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1270),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1270),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1362),
.B(n_1385),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1300),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1381),
.A2(n_1338),
.B(n_1302),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1362),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1315),
.A2(n_1336),
.B1(n_1340),
.B2(n_1367),
.C(n_1293),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1268),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1268),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1340),
.B(n_1325),
.Y(n_1560)
);

AOI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1367),
.A2(n_1293),
.B1(n_1324),
.B2(n_1312),
.C(n_1304),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1325),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1302),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1301),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1258),
.A2(n_774),
.B1(n_971),
.B2(n_928),
.Y(n_1565)
);

OR2x6_ASAP7_75t_L g1566 ( 
.A(n_1285),
.B(n_1392),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1318),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1284),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1313),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1280),
.A2(n_971),
.B(n_928),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1284),
.B(n_1313),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1341),
.B(n_944),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1263),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1572),
.B(n_1446),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1565),
.A2(n_1427),
.B1(n_1445),
.B2(n_1570),
.C(n_1451),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1427),
.A2(n_1428),
.B1(n_1445),
.B2(n_1463),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1430),
.A2(n_1506),
.B1(n_1452),
.B2(n_1571),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1431),
.B(n_1569),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1563),
.A2(n_1443),
.B1(n_1434),
.B2(n_1441),
.Y(n_1580)
);

BUFx12f_ASAP7_75t_L g1581 ( 
.A(n_1475),
.Y(n_1581)
);

OAI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1454),
.A2(n_1568),
.B1(n_1455),
.B2(n_1438),
.C(n_1472),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1457),
.A2(n_1438),
.B1(n_1481),
.B2(n_1432),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1500),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1432),
.B(n_1518),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1453),
.A2(n_1502),
.B(n_1447),
.C(n_1437),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1521),
.Y(n_1587)
);

AOI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1453),
.A2(n_1456),
.B(n_1459),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1459),
.A2(n_1509),
.B1(n_1466),
.B2(n_1464),
.C(n_1456),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1567),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1448),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1573),
.A2(n_1483),
.B1(n_1484),
.B2(n_1478),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1503),
.A2(n_1465),
.B(n_1508),
.C(n_1496),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1425),
.A2(n_1566),
.B1(n_1435),
.B2(n_1444),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1490),
.A2(n_1468),
.B1(n_1460),
.B2(n_1458),
.Y(n_1597)
);

OAI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1503),
.A2(n_1491),
.B(n_1455),
.C(n_1461),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1495),
.A2(n_1425),
.B1(n_1566),
.B2(n_1435),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1504),
.A2(n_1442),
.B1(n_1440),
.B2(n_1462),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1465),
.A2(n_1477),
.B(n_1523),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1510),
.B(n_1480),
.C(n_1482),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1477),
.A2(n_1528),
.B1(n_1535),
.B2(n_1519),
.C(n_1485),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1444),
.A2(n_1504),
.B1(n_1473),
.B2(n_1429),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1450),
.Y(n_1605)
);

OAI33xp33_ASAP7_75t_L g1606 ( 
.A1(n_1485),
.A2(n_1486),
.A3(n_1474),
.B1(n_1522),
.B2(n_1526),
.B3(n_1527),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1479),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1429),
.A2(n_1436),
.B1(n_1467),
.B2(n_1469),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1512),
.A2(n_1554),
.B1(n_1533),
.B2(n_1494),
.Y(n_1609)
);

CKINVDCx11_ASAP7_75t_R g1610 ( 
.A(n_1471),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1548),
.B(n_1547),
.C(n_1537),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1429),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1519),
.A2(n_1473),
.B(n_1436),
.C(n_1514),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1549),
.A2(n_1497),
.B1(n_1436),
.B2(n_1470),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1479),
.B(n_1488),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1488),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1555),
.A2(n_1533),
.B(n_1548),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1505),
.A2(n_1511),
.B1(n_1520),
.B2(n_1527),
.C(n_1526),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1549),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1498),
.A2(n_1513),
.B1(n_1529),
.B2(n_1507),
.Y(n_1620)
);

AOI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1531),
.A2(n_1541),
.B(n_1525),
.C(n_1555),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1470),
.B(n_1538),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1513),
.A2(n_1507),
.B1(n_1515),
.B2(n_1505),
.Y(n_1623)
);

AOI33xp33_ASAP7_75t_L g1624 ( 
.A1(n_1540),
.A2(n_1524),
.A3(n_1550),
.B1(n_1532),
.B2(n_1546),
.B3(n_1556),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1513),
.A2(n_1476),
.B1(n_1501),
.B2(n_1499),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1513),
.A2(n_1499),
.B1(n_1516),
.B2(n_1536),
.Y(n_1626)
);

BUFx4f_ASAP7_75t_SL g1627 ( 
.A(n_1516),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1517),
.B(n_1449),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1493),
.B(n_1542),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1530),
.A2(n_1562),
.B(n_1557),
.Y(n_1630)
);

INVx3_ASAP7_75t_SL g1631 ( 
.A(n_1536),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1493),
.B(n_1560),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1487),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1520),
.A2(n_1558),
.B1(n_1552),
.B2(n_1551),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1493),
.B(n_1530),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1562),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1544),
.A2(n_1553),
.B1(n_1539),
.B2(n_1534),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1564),
.A2(n_1543),
.B1(n_1557),
.B2(n_1534),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1561),
.B(n_1545),
.C(n_1564),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1439),
.B(n_1426),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1561),
.A2(n_1433),
.B1(n_966),
.B2(n_928),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1565),
.A2(n_971),
.B1(n_928),
.B2(n_966),
.C(n_774),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1521),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1452),
.B(n_1571),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_960),
.B2(n_926),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_960),
.B2(n_926),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1502),
.A2(n_971),
.B(n_928),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1431),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1565),
.A2(n_971),
.B1(n_928),
.B2(n_966),
.C(n_774),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1502),
.A2(n_971),
.B(n_928),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1521),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1495),
.B(n_1309),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1452),
.B(n_1571),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1565),
.A2(n_572),
.B1(n_574),
.B2(n_966),
.C(n_737),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1502),
.A2(n_971),
.B(n_928),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1428),
.A2(n_1258),
.B1(n_774),
.B2(n_966),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1452),
.B(n_1571),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_960),
.B2(n_926),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1448),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1428),
.A2(n_1258),
.B1(n_774),
.B2(n_966),
.Y(n_1669)
);

BUFx5_ASAP7_75t_L g1670 ( 
.A(n_1559),
.Y(n_1670)
);

AOI222xp33_ASAP7_75t_L g1671 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_737),
.B2(n_942),
.C1(n_866),
.C2(n_960),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1502),
.A2(n_971),
.B(n_928),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1565),
.A2(n_572),
.B1(n_574),
.B2(n_966),
.C(n_737),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1429),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1451),
.A2(n_971),
.B(n_928),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1565),
.A2(n_971),
.B1(n_928),
.B2(n_774),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1428),
.A2(n_1258),
.B1(n_774),
.B2(n_966),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1521),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1489),
.B(n_1492),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1565),
.A2(n_966),
.B1(n_971),
.B2(n_928),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1565),
.A2(n_971),
.B1(n_928),
.B2(n_966),
.C(n_774),
.Y(n_1685)
);

CKINVDCx11_ASAP7_75t_R g1686 ( 
.A(n_1567),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1428),
.A2(n_575),
.B1(n_774),
.B2(n_871),
.C(n_857),
.Y(n_1687)
);

AOI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1565),
.A2(n_574),
.B(n_966),
.C(n_572),
.Y(n_1688)
);

A2O1A1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1451),
.A2(n_971),
.B(n_928),
.C(n_774),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1565),
.B(n_1280),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1445),
.A2(n_774),
.B(n_1257),
.C(n_737),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1521),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1565),
.A2(n_572),
.B1(n_574),
.B2(n_966),
.C(n_737),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1565),
.A2(n_572),
.B1(n_574),
.B2(n_966),
.C(n_737),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1565),
.B(n_1280),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1565),
.B(n_1280),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1441),
.B(n_1572),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1635),
.B(n_1628),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1632),
.B(n_1629),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1670),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1657),
.B(n_1617),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1688),
.A2(n_1659),
.B1(n_1675),
.B2(n_1693),
.C(n_1695),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1592),
.B(n_1694),
.Y(n_1705)
);

CKINVDCx16_ASAP7_75t_R g1706 ( 
.A(n_1694),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1630),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1618),
.B(n_1594),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1636),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1611),
.B(n_1602),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1577),
.A2(n_1665),
.B1(n_1645),
.B2(n_1661),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1622),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1593),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1639),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1605),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1577),
.A2(n_1672),
.B1(n_1666),
.B2(n_1665),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1621),
.B(n_1601),
.Y(n_1719)
);

NAND2x1p5_ASAP7_75t_L g1720 ( 
.A(n_1652),
.B(n_1655),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1668),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1603),
.B(n_1620),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1624),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1595),
.B(n_1597),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1588),
.A2(n_1662),
.B(n_1673),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1631),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1641),
.B(n_1599),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1619),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1586),
.B(n_1623),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_SL g1730 ( 
.A(n_1598),
.B(n_1690),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1596),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1648),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1641),
.B(n_1589),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1658),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1664),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1696),
.B(n_1697),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1678),
.A2(n_1625),
.B(n_1575),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1596),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1609),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1698),
.B(n_1626),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1613),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1585),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1579),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1580),
.B(n_1616),
.Y(n_1744)
);

INVxp67_ASAP7_75t_R g1745 ( 
.A(n_1600),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1643),
.A2(n_1651),
.B1(n_1647),
.B2(n_1660),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1679),
.B(n_1647),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1587),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1582),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1646),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1633),
.B(n_1692),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1656),
.Y(n_1752)
);

AOI22x1_ASAP7_75t_L g1753 ( 
.A1(n_1710),
.A2(n_1671),
.B1(n_1584),
.B2(n_1591),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1703),
.A2(n_1667),
.B1(n_1649),
.B2(n_1650),
.C(n_1651),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1713),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1728),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1705),
.B(n_1681),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1721),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1703),
.A2(n_1687),
.B(n_1583),
.C(n_1691),
.Y(n_1759)
);

NAND4xp25_ASAP7_75t_SL g1760 ( 
.A(n_1703),
.B(n_1674),
.C(n_1672),
.D(n_1666),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1713),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1711),
.A2(n_1642),
.B1(n_1685),
.B2(n_1654),
.Y(n_1762)
);

INVx3_ASAP7_75t_SL g1763 ( 
.A(n_1709),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1743),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1710),
.A2(n_1643),
.B1(n_1684),
.B2(n_1683),
.C(n_1645),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1716),
.Y(n_1766)
);

AOI31xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1710),
.A2(n_1674),
.A3(n_1660),
.B(n_1661),
.Y(n_1767)
);

CKINVDCx6p67_ASAP7_75t_R g1768 ( 
.A(n_1728),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_SL g1769 ( 
.A(n_1710),
.B(n_1684),
.C(n_1683),
.Y(n_1769)
);

AOI222xp33_ASAP7_75t_L g1770 ( 
.A1(n_1711),
.A2(n_1680),
.B1(n_1663),
.B2(n_1669),
.C1(n_1676),
.C2(n_1679),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1704),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1711),
.A2(n_1583),
.B1(n_1578),
.B2(n_1608),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1723),
.A2(n_1676),
.B(n_1689),
.C(n_1653),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1728),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1732),
.B(n_1615),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_R g1776 ( 
.A(n_1715),
.B(n_1612),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1715),
.B(n_1578),
.C(n_1574),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1736),
.B(n_1677),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1718),
.A2(n_1606),
.B1(n_1607),
.B2(n_1604),
.C(n_1612),
.Y(n_1779)
);

NAND4xp25_ASAP7_75t_L g1780 ( 
.A(n_1723),
.B(n_1614),
.C(n_1677),
.D(n_1590),
.Y(n_1780)
);

AOI31xp33_ASAP7_75t_L g1781 ( 
.A1(n_1718),
.A2(n_1576),
.A3(n_1682),
.B(n_1590),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1644),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1718),
.A2(n_1746),
.B1(n_1729),
.B2(n_1747),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1742),
.B(n_1644),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1743),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1704),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1721),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1746),
.A2(n_1627),
.B1(n_1682),
.B2(n_1581),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1746),
.A2(n_1610),
.B1(n_1627),
.B2(n_1686),
.C(n_1715),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1732),
.B(n_1734),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1699),
.B(n_1732),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1743),
.Y(n_1792)
);

OAI31xp33_ASAP7_75t_L g1793 ( 
.A1(n_1729),
.A2(n_1708),
.A3(n_1722),
.B(n_1724),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1729),
.A2(n_1722),
.B1(n_1747),
.B2(n_1708),
.Y(n_1794)
);

OAI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1747),
.A2(n_1741),
.B1(n_1749),
.B2(n_1745),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1729),
.A2(n_1722),
.B1(n_1708),
.B2(n_1749),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1720),
.B(n_1719),
.Y(n_1797)
);

BUFx10_ASAP7_75t_L g1798 ( 
.A(n_1726),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1716),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_SL g1800 ( 
.A1(n_1729),
.A2(n_1730),
.B1(n_1708),
.B2(n_1722),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1742),
.B(n_1734),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1728),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1728),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1716),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1734),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1729),
.A2(n_1749),
.B1(n_1733),
.B2(n_1741),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1729),
.A2(n_1730),
.B1(n_1724),
.B2(n_1733),
.Y(n_1807)
);

OAI31xp33_ASAP7_75t_L g1808 ( 
.A1(n_1724),
.A2(n_1741),
.A3(n_1733),
.B(n_1719),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1723),
.A2(n_1720),
.B1(n_1719),
.B2(n_1739),
.C(n_1736),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1758),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1792),
.B(n_1699),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1763),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1791),
.B(n_1764),
.Y(n_1813)
);

AND2x4_ASAP7_75t_SL g1814 ( 
.A(n_1798),
.B(n_1768),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1801),
.B(n_1736),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1771),
.B(n_1719),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_1805),
.Y(n_1817)
);

NOR2x1_ASAP7_75t_L g1818 ( 
.A(n_1809),
.B(n_1750),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1771),
.B(n_1700),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1790),
.B(n_1739),
.Y(n_1820)
);

NAND2x1p5_ASAP7_75t_L g1821 ( 
.A(n_1778),
.B(n_1725),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1776),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1771),
.B(n_1700),
.Y(n_1823)
);

NAND2x1_ASAP7_75t_SL g1824 ( 
.A(n_1786),
.B(n_1702),
.Y(n_1824)
);

AND2x4_ASAP7_75t_SL g1825 ( 
.A(n_1798),
.B(n_1705),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1787),
.B(n_1699),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1700),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1755),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1761),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1759),
.B(n_1725),
.C(n_1724),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1766),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1786),
.B(n_1700),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1702),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1799),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1807),
.B(n_1706),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1701),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.B(n_1702),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1774),
.B(n_1725),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1797),
.B(n_1702),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1775),
.B(n_1707),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1802),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1774),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1757),
.B(n_1707),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1782),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1800),
.B(n_1706),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1757),
.B(n_1707),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1776),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1783),
.B(n_1735),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1798),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1803),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1812),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1810),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1828),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1846),
.B(n_1808),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1846),
.B(n_1748),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1828),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1849),
.B(n_1768),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1810),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1849),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1822),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1825),
.B(n_1803),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1820),
.B(n_1709),
.Y(n_1864)
);

OAI32xp33_ASAP7_75t_L g1865 ( 
.A1(n_1830),
.A2(n_1762),
.A3(n_1777),
.B1(n_1773),
.B2(n_1765),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1819),
.B(n_1704),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1814),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1850),
.B(n_1748),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1814),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1847),
.B(n_1795),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1828),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1850),
.B(n_1748),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1812),
.B(n_1754),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_SL g1874 ( 
.A(n_1836),
.B(n_1712),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1828),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1819),
.B(n_1704),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1830),
.B(n_1748),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1818),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1810),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1847),
.B(n_1793),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1815),
.B(n_1748),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1819),
.B(n_1704),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1836),
.A2(n_1760),
.B1(n_1769),
.B2(n_1762),
.Y(n_1883)
);

NOR3xp33_ASAP7_75t_L g1884 ( 
.A(n_1818),
.B(n_1789),
.C(n_1772),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1829),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1829),
.Y(n_1886)
);

AND2x4_ASAP7_75t_SL g1887 ( 
.A(n_1834),
.B(n_1705),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1829),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1829),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1822),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1810),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1815),
.B(n_1752),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1820),
.B(n_1709),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1823),
.B(n_1704),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1837),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1884),
.B(n_1753),
.C(n_1770),
.Y(n_1896)
);

OAI33xp33_ASAP7_75t_L g1897 ( 
.A1(n_1880),
.A2(n_1870),
.A3(n_1890),
.B1(n_1856),
.B2(n_1877),
.B3(n_1865),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1864),
.B(n_1832),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1853),
.B(n_1873),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1862),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1859),
.B(n_1845),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1859),
.B(n_1845),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1862),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1855),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_R g1906 ( 
.A(n_1853),
.B(n_1706),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1878),
.Y(n_1907)
);

BUFx12f_ASAP7_75t_L g1908 ( 
.A(n_1853),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1883),
.B(n_1861),
.Y(n_1909)
);

AND2x2_ASAP7_75t_SL g1910 ( 
.A(n_1883),
.B(n_1725),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1861),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_R g1912 ( 
.A(n_1863),
.B(n_1756),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1868),
.B(n_1842),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1864),
.B(n_1893),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1855),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1893),
.B(n_1872),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_SL g1917 ( 
.A(n_1865),
.B(n_1796),
.C(n_1794),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1881),
.B(n_1811),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1874),
.B(n_1845),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1892),
.B(n_1842),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_L g1921 ( 
.A(n_1867),
.B(n_1737),
.C(n_1788),
.Y(n_1921)
);

NAND3xp33_ASAP7_75t_L g1922 ( 
.A(n_1857),
.B(n_1796),
.C(n_1794),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1867),
.B(n_1811),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1874),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1869),
.B(n_1811),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1869),
.B(n_1720),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1863),
.B(n_1824),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1858),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1887),
.B(n_1848),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_R g1930 ( 
.A(n_1863),
.B(n_1756),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1858),
.Y(n_1931)
);

NOR2x1p5_ASAP7_75t_L g1932 ( 
.A(n_1863),
.B(n_1780),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1871),
.B(n_1806),
.C(n_1779),
.D(n_1733),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1871),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1875),
.Y(n_1935)
);

NAND2x1_ASAP7_75t_L g1936 ( 
.A(n_1866),
.B(n_1823),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1866),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1875),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1885),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1876),
.B(n_1842),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1911),
.Y(n_1941)
);

OAI32xp33_ASAP7_75t_L g1942 ( 
.A1(n_1909),
.A2(n_1840),
.A3(n_1821),
.B1(n_1720),
.B2(n_1806),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1919),
.B(n_1887),
.Y(n_1943)
);

AOI21xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1896),
.A2(n_1781),
.B(n_1821),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1911),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1906),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1930),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1900),
.Y(n_1948)
);

AOI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1897),
.A2(n_1840),
.B1(n_1816),
.B2(n_1717),
.C(n_1821),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1922),
.B(n_1901),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1904),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1908),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1899),
.B(n_1816),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1897),
.A2(n_1725),
.B1(n_1705),
.B2(n_1727),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1932),
.B(n_1816),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1917),
.B(n_1887),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1917),
.A2(n_1821),
.B(n_1840),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1910),
.A2(n_1840),
.B(n_1737),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1931),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1907),
.B(n_1823),
.Y(n_1960)
);

OAI21xp33_ASAP7_75t_L g1961 ( 
.A1(n_1910),
.A2(n_1933),
.B(n_1907),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1931),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1923),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1902),
.B(n_1827),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1935),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1912),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1937),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1935),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1903),
.B(n_1827),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1925),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1914),
.Y(n_1971)
);

NOR2xp67_ASAP7_75t_SL g1972 ( 
.A(n_1898),
.B(n_1725),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1905),
.Y(n_1973)
);

AOI21xp33_ASAP7_75t_L g1974 ( 
.A1(n_1924),
.A2(n_1725),
.B(n_1851),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1921),
.Y(n_1975)
);

AOI211x1_ASAP7_75t_SL g1976 ( 
.A1(n_1940),
.A2(n_1851),
.B(n_1751),
.C(n_1879),
.Y(n_1976)
);

OAI221xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1924),
.A2(n_1717),
.B1(n_1767),
.B2(n_1727),
.C(n_1839),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1941),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1943),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1977),
.A2(n_1936),
.B1(n_1921),
.B2(n_1929),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_L g1981 ( 
.A1(n_1961),
.A2(n_1717),
.B1(n_1720),
.B2(n_1737),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1948),
.B(n_1916),
.Y(n_1982)
);

INVxp67_ASAP7_75t_L g1983 ( 
.A(n_1941),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1945),
.B(n_1913),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1946),
.B(n_1876),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1956),
.A2(n_1927),
.B1(n_1717),
.B2(n_1926),
.Y(n_1986)
);

NOR2x1_ASAP7_75t_L g1987 ( 
.A(n_1952),
.B(n_1915),
.Y(n_1987)
);

AOI321xp33_ASAP7_75t_L g1988 ( 
.A1(n_1944),
.A2(n_1727),
.A3(n_1714),
.B1(n_1731),
.B2(n_1738),
.C(n_1744),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1959),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1971),
.B(n_1920),
.Y(n_1990)
);

A2O1A1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1956),
.A2(n_1737),
.B(n_1824),
.C(n_1751),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1959),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1970),
.B(n_1918),
.Y(n_1993)
);

NOR2xp67_ASAP7_75t_L g1994 ( 
.A(n_1966),
.B(n_1970),
.Y(n_1994)
);

XOR2x2_ASAP7_75t_L g1995 ( 
.A(n_1947),
.B(n_1730),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1962),
.Y(n_1996)
);

INVxp67_ASAP7_75t_L g1997 ( 
.A(n_1965),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1951),
.B(n_1963),
.Y(n_1998)
);

NAND4xp25_ASAP7_75t_L g1999 ( 
.A(n_1950),
.B(n_1751),
.C(n_1938),
.D(n_1934),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1975),
.B(n_1882),
.Y(n_2000)
);

OR2x6_ASAP7_75t_L g2001 ( 
.A(n_1958),
.B(n_1926),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1943),
.B(n_1882),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1949),
.A2(n_1926),
.B(n_1928),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1942),
.A2(n_1939),
.B(n_1745),
.Y(n_2004)
);

NOR2x1_ASAP7_75t_L g2005 ( 
.A(n_1987),
.B(n_1962),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1994),
.Y(n_2006)
);

A2O1A1Ixp33_ASAP7_75t_L g2007 ( 
.A1(n_1988),
.A2(n_1957),
.B(n_1954),
.C(n_1942),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1981),
.A2(n_1974),
.B(n_1955),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1998),
.B(n_1953),
.Y(n_2009)
);

BUFx2_ASAP7_75t_SL g2010 ( 
.A(n_1995),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1981),
.B(n_1968),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1993),
.B(n_1967),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1978),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1980),
.A2(n_1967),
.B1(n_1960),
.B2(n_1972),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1989),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1985),
.B(n_1973),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1979),
.B(n_1894),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1983),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1982),
.B(n_1964),
.Y(n_2019)
);

OAI322xp33_ASAP7_75t_L g2020 ( 
.A1(n_1983),
.A2(n_1969),
.A3(n_1976),
.B1(n_1817),
.B2(n_1813),
.C1(n_1851),
.C2(n_1972),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1992),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1999),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1996),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1997),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_2005),
.Y(n_2025)
);

OAI321xp33_ASAP7_75t_L g2026 ( 
.A1(n_2014),
.A2(n_2003),
.A3(n_1986),
.B1(n_2001),
.B2(n_1997),
.C(n_1991),
.Y(n_2026)
);

OAI211xp5_ASAP7_75t_SL g2027 ( 
.A1(n_2022),
.A2(n_1991),
.B(n_2004),
.C(n_1990),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2018),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_2024),
.B(n_1984),
.Y(n_2029)
);

NOR3x1_ASAP7_75t_L g2030 ( 
.A(n_2012),
.B(n_2000),
.C(n_1843),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_2024),
.Y(n_2031)
);

XNOR2xp5_ASAP7_75t_SL g2032 ( 
.A(n_2018),
.B(n_1851),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_2007),
.B(n_2002),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2007),
.B(n_1814),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2006),
.B(n_1894),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2016),
.B(n_2001),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2016),
.Y(n_2037)
);

A2O1A1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_2025),
.A2(n_2011),
.B(n_2008),
.C(n_2009),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_2034),
.A2(n_2011),
.B(n_2021),
.C(n_2023),
.Y(n_2039)
);

OAI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2033),
.A2(n_2009),
.B(n_2001),
.Y(n_2040)
);

AOI211xp5_ASAP7_75t_L g2041 ( 
.A1(n_2026),
.A2(n_2020),
.B(n_2015),
.C(n_2013),
.Y(n_2041)
);

AOI221xp5_ASAP7_75t_L g2042 ( 
.A1(n_2027),
.A2(n_2010),
.B1(n_2019),
.B2(n_2017),
.C(n_1844),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_2029),
.A2(n_1844),
.B(n_1891),
.C(n_1854),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2029),
.A2(n_1843),
.B1(n_1889),
.B2(n_1888),
.C(n_1886),
.Y(n_2044)
);

AOI311xp33_ASAP7_75t_L g2045 ( 
.A1(n_2037),
.A2(n_2028),
.A3(n_2036),
.B(n_2035),
.C(n_2030),
.Y(n_2045)
);

NAND3x1_ASAP7_75t_L g2046 ( 
.A(n_2031),
.B(n_1895),
.C(n_1889),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_SL g2047 ( 
.A(n_2032),
.B(n_1814),
.Y(n_2047)
);

A2O1A1Ixp33_ASAP7_75t_L g2048 ( 
.A1(n_2025),
.A2(n_1824),
.B(n_1825),
.C(n_1852),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_2034),
.B(n_1750),
.C(n_1752),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2046),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2038),
.B(n_1885),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2040),
.A2(n_1852),
.B(n_1750),
.C(n_1888),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2042),
.B(n_1886),
.Y(n_2053)
);

OAI311xp33_ASAP7_75t_L g2054 ( 
.A1(n_2039),
.A2(n_1852),
.A3(n_1834),
.B1(n_1841),
.C1(n_1839),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2043),
.Y(n_2055)
);

CKINVDCx6p67_ASAP7_75t_R g2056 ( 
.A(n_2055),
.Y(n_2056)
);

NOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2050),
.B(n_2049),
.Y(n_2057)
);

NAND2x1p5_ASAP7_75t_L g2058 ( 
.A(n_2051),
.B(n_2047),
.Y(n_2058)
);

OAI21xp33_ASAP7_75t_L g2059 ( 
.A1(n_2052),
.A2(n_2041),
.B(n_2048),
.Y(n_2059)
);

NOR2x1_ASAP7_75t_L g2060 ( 
.A(n_2053),
.B(n_2045),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2054),
.A2(n_2044),
.B1(n_1825),
.B2(n_1745),
.Y(n_2061)
);

OA22x2_ASAP7_75t_L g2062 ( 
.A1(n_2050),
.A2(n_1860),
.B1(n_1891),
.B2(n_1854),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_SL g2063 ( 
.A(n_2058),
.B(n_1841),
.C(n_1834),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2059),
.B(n_1841),
.C(n_1839),
.D(n_1740),
.Y(n_2064)
);

NAND2x1p5_ASAP7_75t_L g2065 ( 
.A(n_2057),
.B(n_1726),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2060),
.A2(n_1852),
.B1(n_1825),
.B2(n_1879),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_2056),
.B(n_1852),
.C(n_1752),
.Y(n_2067)
);

AO22x2_ASAP7_75t_L g2068 ( 
.A1(n_2062),
.A2(n_1891),
.B1(n_1854),
.B2(n_1860),
.Y(n_2068)
);

NOR3xp33_ASAP7_75t_SL g2069 ( 
.A(n_2063),
.B(n_2064),
.C(n_2065),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_SL g2070 ( 
.A1(n_2068),
.A2(n_2061),
.B1(n_1726),
.B2(n_1838),
.Y(n_2070)
);

XNOR2x1_ASAP7_75t_L g2071 ( 
.A(n_2066),
.B(n_1740),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_L g2072 ( 
.A(n_2067),
.B(n_1752),
.C(n_1784),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2071),
.A2(n_1879),
.B1(n_1860),
.B2(n_1895),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2073),
.B(n_2069),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_2074),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_2074),
.Y(n_2076)
);

AOI222xp33_ASAP7_75t_L g2077 ( 
.A1(n_2075),
.A2(n_2070),
.B1(n_2072),
.B2(n_1727),
.C1(n_1833),
.C2(n_1827),
.Y(n_2077)
);

NAND3xp33_ASAP7_75t_L g2078 ( 
.A(n_2076),
.B(n_1817),
.C(n_1726),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2078),
.Y(n_2079)
);

OAI222xp33_ASAP7_75t_L g2080 ( 
.A1(n_2077),
.A2(n_1817),
.B1(n_1813),
.B2(n_1826),
.C1(n_1833),
.C2(n_1835),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2079),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_R g2082 ( 
.A1(n_2081),
.A2(n_2080),
.B1(n_1813),
.B2(n_1833),
.C(n_1826),
.Y(n_2082)
);

AOI211xp5_ASAP7_75t_L g2083 ( 
.A1(n_2082),
.A2(n_1726),
.B(n_1831),
.C(n_1835),
.Y(n_2083)
);


endmodule