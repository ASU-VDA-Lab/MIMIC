module fake_jpeg_7787_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_9),
.B(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_24),
.C(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_44),
.B1(n_23),
.B2(n_22),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_46),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_36),
.B1(n_31),
.B2(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_36),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_66),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_71),
.B(n_4),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_33),
.B(n_20),
.C(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_65),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_32),
.B1(n_19),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_38),
.B1(n_47),
.B2(n_21),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_18),
.A3(n_13),
.B1(n_30),
.B2(n_16),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_6),
.Y(n_92)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_73),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_1),
.Y(n_69)
);

NOR2xp67_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_57),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_21),
.B(n_15),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_80),
.B(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_82),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_55),
.B1(n_62),
.B2(n_77),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_38),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_47),
.B1(n_21),
.B2(n_15),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_59),
.B1(n_65),
.B2(n_64),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_72),
.B1(n_69),
.B2(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_72),
.C(n_71),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_80),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_74),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_78),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_80),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_96),
.B1(n_84),
.B2(n_105),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_92),
.C(n_79),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_123),
.B1(n_116),
.B2(n_109),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_97),
.B(n_99),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_120),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_106),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_124),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_93),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_106),
.B1(n_89),
.B2(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_130),
.C(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_115),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_108),
.B(n_119),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_91),
.B1(n_129),
.B2(n_84),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_111),
.C(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_125),
.B(n_6),
.Y(n_138)
);

OAI221xp5_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_134),
.B1(n_75),
.B2(n_5),
.C(n_8),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_11),
.Y(n_141)
);

OAI31xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_139),
.A3(n_11),
.B(n_5),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_136),
.Y(n_143)
);


endmodule