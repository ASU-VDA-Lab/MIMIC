module fake_ariane_2700_n_1427 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1427);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1427;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

INVx1_ASAP7_75t_L g365 ( 
.A(n_71),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_72),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_90),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_248),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_183),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_352),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_255),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_219),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_28),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_194),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_98),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_10),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_151),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_311),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_125),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_171),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_12),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_104),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_284),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_33),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_295),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_187),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_147),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_47),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_24),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_207),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_117),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_6),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_238),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_3),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_184),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_251),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_359),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_231),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_29),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_68),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_73),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_109),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_162),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_203),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_110),
.Y(n_411)
);

BUFx8_ASAP7_75t_SL g412 ( 
.A(n_135),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_213),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_195),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_299),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_304),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_280),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_9),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_30),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_321),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_214),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_56),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_157),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_289),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_96),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_9),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_78),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_19),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_256),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_357),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_285),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_89),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_247),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_60),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_201),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_22),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_286),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_227),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_54),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_12),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_314),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_14),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_4),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_66),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_113),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_230),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_166),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_345),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_164),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_138),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_102),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_22),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_296),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_202),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_52),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_354),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_268),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_149),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_229),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_177),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_216),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_364),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_239),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_143),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_59),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_242),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_215),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_35),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_199),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_101),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_156),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_81),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_356),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_358),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_145),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_282),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_277),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_337),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_265),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_86),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_217),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_121),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_155),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_198),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_322),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_128),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_20),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_85),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_346),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_13),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_241),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_30),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_11),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_33),
.Y(n_499)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_223),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_236),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_180),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_270),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_318),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_120),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_148),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_161),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_348),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_56),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_188),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_193),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_224),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_220),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_234),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_133),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_95),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_54),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_330),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_326),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_1),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_112),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_197),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_80),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_222),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_2),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_141),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_204),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_75),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_92),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_266),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_233),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_309),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_130),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_57),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_185),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_288),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_331),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_131),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_111),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_355),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_106),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_16),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_310),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_24),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_67),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_210),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_281),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_146),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_308),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_362),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_4),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_132),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_341),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_324),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_253),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_225),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_273),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_305),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_267),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_43),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_323),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_41),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_172),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_11),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_118),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_290),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_500),
.B(n_0),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_414),
.B(n_0),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_492),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_473),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_412),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_428),
.Y(n_573)
);

BUFx6f_ASAP7_75t_SL g574 ( 
.A(n_394),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_412),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_379),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_560),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_380),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_405),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_457),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_397),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_403),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_408),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_449),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_461),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_470),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_474),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_497),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_476),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_489),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_504),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_519),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_545),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_374),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_384),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_388),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_394),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

INVxp33_ASAP7_75t_SL g601 ( 
.A(n_392),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_393),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_396),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_418),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_542),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_562),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_419),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_424),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_424),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_500),
.B(n_1),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_430),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_443),
.B(n_2),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_439),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_443),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_444),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_446),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_447),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_482),
.B(n_546),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_460),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_498),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_520),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_517),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_544),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_551),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_564),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_394),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_368),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_450),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_370),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_399),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_450),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_525),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_450),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_371),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_455),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_455),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_372),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_525),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_376),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_366),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_442),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_475),
.Y(n_645)
);

CKINVDCx16_ASAP7_75t_R g646 ( 
.A(n_455),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_367),
.B(n_3),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_510),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_510),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_391),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_365),
.Y(n_652)
);

CKINVDCx16_ASAP7_75t_R g653 ( 
.A(n_391),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_406),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_406),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_369),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_373),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_375),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_R g659 ( 
.A(n_381),
.B(n_382),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_377),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_378),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_386),
.Y(n_662)
);

BUFx2_ASAP7_75t_SL g663 ( 
.A(n_463),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_463),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_383),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_533),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_533),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_608),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_576),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_578),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_579),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_571),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_652),
.A2(n_395),
.B(n_390),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_581),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_580),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_582),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_609),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_614),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_620),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_584),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_653),
.B(n_654),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_583),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_587),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_571),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_623),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_595),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_588),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_600),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_605),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_626),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_606),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_570),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_518),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_R g697 ( 
.A(n_596),
.B(n_404),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_586),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_647),
.B(n_367),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_573),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_590),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_592),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_594),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_635),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_633),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_663),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_630),
.B(n_409),
.Y(n_707)
);

OA21x2_ASAP7_75t_L g708 ( 
.A1(n_656),
.A2(n_422),
.B(n_410),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_641),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_657),
.B(n_432),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_658),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_572),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_660),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_575),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_661),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_625),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_585),
.Y(n_717)
);

XOR2xp5_ASAP7_75t_L g718 ( 
.A(n_591),
.B(n_385),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_593),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_662),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_645),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_612),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_632),
.B(n_423),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_651),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_628),
.Y(n_726)
);

INVxp33_ASAP7_75t_SL g727 ( 
.A(n_659),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_637),
.B(n_427),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_644),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_640),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_577),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_642),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_665),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_655),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_597),
.B(n_387),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_568),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_567),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_610),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_586),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_598),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_602),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_574),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_603),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_569),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_604),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_574),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_607),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_R g749 ( 
.A(n_611),
.B(n_436),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_613),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_615),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_SL g752 ( 
.A(n_664),
.B(n_666),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_733),
.B(n_601),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_705),
.B(n_599),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_730),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_726),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_743),
.B(n_432),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_695),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_682),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_696),
.A2(n_616),
.B1(n_621),
.B2(n_618),
.Y(n_760)
);

AND2x6_ASAP7_75t_L g761 ( 
.A(n_747),
.B(n_434),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_751),
.B(n_634),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_738),
.B(n_646),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_677),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_677),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_705),
.B(n_622),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_730),
.B(n_434),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_677),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_739),
.A2(n_666),
.B1(n_664),
.B2(n_667),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_745),
.B(n_624),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_741),
.Y(n_771)
);

INVxp33_ASAP7_75t_SL g772 ( 
.A(n_670),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_700),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_696),
.A2(n_749),
.B1(n_697),
.B2(n_746),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_737),
.A2(n_667),
.B1(n_631),
.B2(n_629),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_750),
.B(n_398),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_725),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_677),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_678),
.Y(n_779)
);

AND3x2_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_521),
.C(n_629),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

BUFx10_ASAP7_75t_L g782 ( 
.A(n_742),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_745),
.B(n_627),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_734),
.B(n_389),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_731),
.B(n_732),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_707),
.B(n_402),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_729),
.B(n_631),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_744),
.B(n_636),
.Y(n_788)
);

AND2x2_ASAP7_75t_SL g789 ( 
.A(n_716),
.B(n_638),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_671),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_748),
.B(n_639),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_710),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_675),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_678),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_650),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_728),
.B(n_628),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_706),
.B(n_471),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_683),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_727),
.B(n_438),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_689),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_697),
.B(n_454),
.C(n_440),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_698),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_711),
.B(n_506),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_736),
.B(n_400),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_735),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_708),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_464),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_720),
.B(n_472),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_678),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_674),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_678),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_699),
.B(n_541),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_687),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_713),
.B(n_480),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_687),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_723),
.B(n_453),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_691),
.A2(n_566),
.B1(n_527),
.B2(n_532),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_715),
.B(n_505),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_687),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_718),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_687),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_699),
.B(n_692),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_699),
.B(n_401),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_709),
.B(n_538),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_668),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_694),
.B(n_722),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_699),
.B(n_407),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_699),
.B(n_411),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_676),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_679),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_709),
.B(n_539),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_736),
.B(n_413),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_684),
.B(n_415),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_680),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_693),
.B(n_540),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_704),
.B(n_543),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_712),
.B(n_714),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_710),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_708),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_673),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_685),
.B(n_548),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_754),
.B(n_690),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_786),
.B(n_710),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_758),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_774),
.B(n_701),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_806),
.B(n_702),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_767),
.A2(n_749),
.B1(n_710),
.B2(n_708),
.Y(n_848)
);

AO22x1_ASAP7_75t_L g849 ( 
.A1(n_796),
.A2(n_703),
.B1(n_740),
.B2(n_719),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_755),
.B(n_710),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_811),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_763),
.B(n_717),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_781),
.A2(n_559),
.B(n_561),
.C(n_554),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_797),
.B(n_752),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_766),
.B(n_755),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_802),
.A2(n_752),
.B1(n_493),
.B2(n_503),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_798),
.B(n_416),
.Y(n_857)
);

BUFx4f_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_760),
.B(n_698),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_800),
.B(n_417),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_756),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_753),
.B(n_420),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_790),
.A2(n_421),
.B1(n_426),
.B2(n_425),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_831),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_759),
.B(n_672),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_808),
.B(n_762),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_793),
.B(n_429),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_794),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_772),
.B(n_672),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_835),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_799),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_767),
.A2(n_431),
.B1(n_435),
.B2(n_433),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_842),
.B(n_830),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_832),
.B(n_437),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_827),
.B(n_441),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_826),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_823),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_764),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_770),
.B(n_686),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_804),
.B(n_445),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_803),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_767),
.B(n_448),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_783),
.B(n_686),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_826),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_764),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_782),
.B(n_451),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_767),
.B(n_452),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_777),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_809),
.B(n_456),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_815),
.B(n_458),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_782),
.B(n_459),
.Y(n_894)
);

OAI22xp33_ASAP7_75t_L g895 ( 
.A1(n_825),
.A2(n_818),
.B1(n_836),
.B2(n_785),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_SL g896 ( 
.A1(n_769),
.A2(n_465),
.B1(n_466),
.B2(n_462),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_834),
.B(n_467),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_819),
.A2(n_493),
.B1(n_503),
.B2(n_398),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_817),
.A2(n_493),
.B1(n_503),
.B2(n_398),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_787),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_764),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_817),
.B(n_468),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_778),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_778),
.B(n_469),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_787),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_765),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_768),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_795),
.Y(n_908)
);

AND2x6_ASAP7_75t_L g909 ( 
.A(n_807),
.B(n_398),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_795),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_784),
.B(n_477),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_837),
.B(n_779),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_795),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_814),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_839),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_807),
.A2(n_479),
.B(n_478),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_838),
.B(n_481),
.Y(n_917)
);

BUFx6f_ASAP7_75t_SL g918 ( 
.A(n_789),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_788),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_810),
.B(n_483),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_791),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_812),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_775),
.B(n_5),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_814),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_757),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_839),
.A2(n_485),
.B1(n_486),
.B2(n_484),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_813),
.A2(n_503),
.B1(n_493),
.B2(n_488),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_820),
.B(n_487),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_805),
.A2(n_491),
.B1(n_494),
.B2(n_490),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_814),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_833),
.B(n_496),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_816),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_841),
.A2(n_502),
.B(n_507),
.C(n_501),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_816),
.Y(n_934)
);

AND2x6_ASAP7_75t_SL g935 ( 
.A(n_780),
.B(n_821),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_816),
.B(n_822),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_R g937 ( 
.A(n_822),
.B(n_776),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_822),
.B(n_508),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_886),
.B(n_757),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_847),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_847),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_851),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_867),
.B(n_757),
.Y(n_943)
);

CKINVDCx8_ASAP7_75t_R g944 ( 
.A(n_935),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_884),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_854),
.B(n_757),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_859),
.A2(n_824),
.B1(n_828),
.B2(n_829),
.C(n_511),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_843),
.B(n_761),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_860),
.B(n_863),
.Y(n_949)
);

OR2x6_ASAP7_75t_L g950 ( 
.A(n_891),
.B(n_840),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_861),
.B(n_761),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_845),
.B(n_761),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_858),
.B(n_792),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_865),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_SL g955 ( 
.A(n_919),
.B(n_513),
.C(n_512),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_910),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_910),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_900),
.B(n_761),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_871),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_852),
.B(n_776),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_SL g961 ( 
.A(n_875),
.B(n_841),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_862),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_915),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_910),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_850),
.A2(n_792),
.B(n_515),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_921),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_906),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_858),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_915),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_914),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_914),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_870),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_918),
.B(n_776),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_869),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_905),
.B(n_925),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_907),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_792),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_882),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_914),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_849),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_880),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_918),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_923),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_917),
.B(n_516),
.C(n_514),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_873),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_895),
.B(n_522),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_846),
.B(n_523),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_878),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_874),
.B(n_524),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_896),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_855),
.B(n_889),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_881),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_902),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_896),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_856),
.A2(n_776),
.B1(n_528),
.B2(n_529),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_883),
.B(n_565),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_877),
.A2(n_530),
.B1(n_531),
.B2(n_526),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_922),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_880),
.B(n_535),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_901),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_911),
.B(n_536),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_874),
.B(n_537),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_901),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_908),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_894),
.B(n_5),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_897),
.B(n_549),
.C(n_547),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_879),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_887),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_903),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_962),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_SL g1012 ( 
.A(n_1008),
.B(n_844),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_949),
.A2(n_876),
.B1(n_892),
.B2(n_926),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_988),
.A2(n_916),
.B(n_853),
.C(n_857),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_965),
.A2(n_936),
.B(n_908),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_961),
.A2(n_931),
.B(n_904),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_913),
.B(n_888),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_991),
.A2(n_893),
.B1(n_926),
.B2(n_848),
.Y(n_1018)
);

OA22x2_ASAP7_75t_L g1019 ( 
.A1(n_995),
.A2(n_848),
.B1(n_868),
.B2(n_930),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_946),
.A2(n_912),
.B(n_932),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_978),
.B(n_983),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_1008),
.A2(n_924),
.B(n_934),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_962),
.B(n_974),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_968),
.B(n_938),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_979),
.A2(n_928),
.B(n_920),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_974),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_940),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_979),
.A2(n_890),
.B(n_885),
.Y(n_1028)
);

AO31x2_ASAP7_75t_L g1029 ( 
.A1(n_943),
.A2(n_933),
.A3(n_864),
.B(n_909),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1002),
.A2(n_929),
.B(n_899),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_986),
.B(n_909),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_940),
.B(n_909),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_940),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_986),
.B(n_909),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_985),
.B(n_927),
.Y(n_1035)
);

BUFx2_ASAP7_75t_SL g1036 ( 
.A(n_941),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_967),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_948),
.B(n_898),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_987),
.A2(n_552),
.B1(n_553),
.B2(n_550),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_942),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_975),
.B(n_937),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_975),
.B(n_6),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_994),
.B(n_7),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_990),
.A2(n_556),
.B(n_555),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_1001),
.A2(n_61),
.B(n_58),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_966),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_997),
.B(n_7),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_954),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_1001),
.A2(n_999),
.B(n_976),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_963),
.A2(n_558),
.B(n_557),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_945),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_963),
.A2(n_63),
.B(n_62),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_959),
.Y(n_1053)
);

AO21x2_ASAP7_75t_L g1054 ( 
.A1(n_1003),
.A2(n_563),
.B(n_65),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_939),
.B(n_8),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_969),
.A2(n_69),
.B(n_64),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_960),
.A2(n_74),
.B(n_70),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1010),
.A2(n_8),
.B(n_10),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1006),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_1009),
.A2(n_977),
.A3(n_970),
.B(n_947),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_992),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_992),
.A2(n_77),
.B(n_76),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_980),
.B(n_17),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_941),
.B(n_18),
.Y(n_1064)
);

AOI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_998),
.A2(n_950),
.B(n_989),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1007),
.A2(n_1006),
.B(n_984),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_950),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_945),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_SL g1069 ( 
.A1(n_970),
.A2(n_18),
.B(n_19),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1011),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1026),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_1017),
.A2(n_969),
.B(n_953),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1028),
.A2(n_996),
.B(n_957),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1047),
.A2(n_972),
.B(n_955),
.C(n_982),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1018),
.A2(n_958),
.B1(n_951),
.B2(n_993),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1051),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1068),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1014),
.A2(n_1013),
.B(n_1030),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1018),
.A2(n_951),
.B1(n_958),
.B2(n_993),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1037),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1040),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1049),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1023),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1021),
.B(n_944),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_1032),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1025),
.A2(n_957),
.B(n_956),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1048),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1053),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1015),
.A2(n_957),
.B(n_956),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1020),
.A2(n_1022),
.B(n_1045),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1027),
.Y(n_1091)
);

INVx6_ASAP7_75t_L g1092 ( 
.A(n_1033),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_1033),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1057),
.A2(n_964),
.B(n_956),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_1031),
.A2(n_971),
.B(n_964),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1052),
.A2(n_971),
.B(n_964),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1046),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1056),
.A2(n_971),
.B(n_981),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1042),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1016),
.A2(n_1058),
.B(n_1055),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1019),
.B(n_981),
.Y(n_1101)
);

INVx8_ASAP7_75t_L g1102 ( 
.A(n_1032),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_1034),
.A2(n_1004),
.B(n_981),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1062),
.A2(n_1005),
.B(n_1004),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_R g1105 ( 
.A(n_1038),
.B(n_973),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1044),
.A2(n_1005),
.B(n_1004),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1027),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_SL g1108 ( 
.A(n_1036),
.B(n_1005),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_1012),
.A2(n_1000),
.B(n_82),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1067),
.A2(n_83),
.B(n_79),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_1040),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_1058),
.A2(n_87),
.B(n_84),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_1066),
.A2(n_20),
.B(n_21),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1064),
.B(n_21),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1066),
.A2(n_23),
.B(n_25),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1029),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1043),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_1041),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1029),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1069),
.A2(n_91),
.B(n_88),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1035),
.A2(n_94),
.B(n_93),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1024),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_1059),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1050),
.A2(n_99),
.B(n_97),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_1102),
.B(n_1063),
.Y(n_1125)
);

AOI22x1_ASAP7_75t_L g1126 ( 
.A1(n_1078),
.A2(n_1059),
.B1(n_1061),
.B2(n_1039),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1081),
.B(n_23),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1080),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1087),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_SL g1130 ( 
.A(n_1115),
.B(n_1039),
.C(n_1065),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1078),
.A2(n_1060),
.B(n_1029),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_R g1132 ( 
.A(n_1076),
.B(n_100),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1083),
.B(n_1060),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_1076),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1102),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1081),
.B(n_25),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1102),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1070),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1071),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_1115),
.A2(n_1054),
.B1(n_27),
.B2(n_28),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1079),
.A2(n_1060),
.B1(n_1054),
.B2(n_29),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1091),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1088),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_1101),
.B(n_363),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_1077),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1122),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1091),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_1097),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1117),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_1122),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1123),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1092),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1101),
.Y(n_1153)
);

OAI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1075),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1123),
.A2(n_1099),
.B1(n_1118),
.B2(n_1079),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1100),
.A2(n_32),
.B(n_34),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1114),
.B(n_34),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1118),
.B(n_35),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1107),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1090),
.A2(n_105),
.B(n_103),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1100),
.A2(n_36),
.B(n_37),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1111),
.B(n_1085),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1111),
.B(n_36),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1112),
.A2(n_37),
.B(n_38),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1103),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1107),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1122),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1113),
.A2(n_38),
.B(n_39),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1103),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1095),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1112),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1122),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1116),
.A2(n_108),
.B(n_107),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1085),
.B(n_40),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_1095),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1084),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1116),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_SL g1178 ( 
.A1(n_1074),
.A2(n_1082),
.B(n_1119),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_1093),
.B(n_45),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1105),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1107),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1138),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1127),
.B(n_1107),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1126),
.A2(n_1074),
.B1(n_1085),
.B2(n_1092),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1136),
.B(n_1085),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1164),
.A2(n_1086),
.B(n_1089),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1130),
.A2(n_1140),
.B1(n_1153),
.B2(n_1141),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1133),
.B(n_1119),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1157),
.B(n_1092),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1129),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1139),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1167),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1146),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1168),
.A2(n_1130),
.B1(n_1161),
.B2(n_1156),
.C(n_1141),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1172),
.B(n_46),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1168),
.A2(n_1108),
.B1(n_1109),
.B2(n_1082),
.C(n_51),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1155),
.A2(n_1109),
.B1(n_1120),
.B2(n_1106),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1154),
.A2(n_1073),
.B1(n_1110),
.B2(n_1121),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1128),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1162),
.B(n_1104),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1134),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1181),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1144),
.A2(n_1124),
.B1(n_1072),
.B2(n_1105),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1164),
.A2(n_1094),
.A3(n_1096),
.B(n_1098),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1142),
.Y(n_1205)
);

BUFx4f_ASAP7_75t_SL g1206 ( 
.A(n_1166),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1149),
.B(n_48),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1175),
.A2(n_49),
.B(n_50),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1146),
.B(n_49),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1144),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1210)
);

OAI211xp5_ASAP7_75t_L g1211 ( 
.A1(n_1180),
.A2(n_53),
.B(n_55),
.C(n_57),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1144),
.A2(n_53),
.B1(n_55),
.B2(n_114),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1156),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1161),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1160),
.A2(n_126),
.B(n_127),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1131),
.A2(n_129),
.B1(n_134),
.B2(n_136),
.Y(n_1216)
);

AOI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1131),
.A2(n_1171),
.B(n_1133),
.Y(n_1217)
);

AOI221xp5_ASAP7_75t_L g1218 ( 
.A1(n_1176),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.C(n_142),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1132),
.A2(n_144),
.B1(n_150),
.B2(n_152),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1143),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1174),
.A2(n_153),
.B(n_154),
.Y(n_1221)
);

AOI321xp33_ASAP7_75t_L g1222 ( 
.A1(n_1151),
.A2(n_158),
.A3(n_159),
.B1(n_160),
.B2(n_163),
.C(n_165),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1177),
.A2(n_1158),
.B1(n_1163),
.B2(n_1174),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1178),
.A2(n_167),
.B(n_168),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1162),
.A2(n_169),
.B(n_170),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1125),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1175),
.A2(n_176),
.B(n_178),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1158),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_1228)
);

AOI222xp33_ASAP7_75t_L g1229 ( 
.A1(n_1163),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.C1(n_191),
.C2(n_192),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1125),
.A2(n_196),
.B1(n_200),
.B2(n_205),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1150),
.B(n_206),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1150),
.B(n_361),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1147),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1179),
.A2(n_1125),
.B1(n_1148),
.B2(n_1135),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1152),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1173),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1145),
.A2(n_212),
.B1(n_218),
.B2(n_221),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1182),
.B(n_1165),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1191),
.B(n_1152),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1199),
.B(n_1220),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1201),
.B(n_1135),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1190),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1192),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1200),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1200),
.Y(n_1245)
);

AOI211x1_ASAP7_75t_L g1246 ( 
.A1(n_1211),
.A2(n_1159),
.B(n_1137),
.C(n_232),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1235),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1188),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1188),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1186),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1217),
.B(n_1170),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1186),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1224),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1183),
.B(n_1169),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1233),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1204),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1189),
.B(n_1173),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1208),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1208),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1204),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1204),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1225),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1217),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1234),
.B(n_1137),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1210),
.A2(n_226),
.B1(n_228),
.B2(n_235),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1223),
.A2(n_1214),
.B(n_1184),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1193),
.B(n_1185),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1195),
.B(n_1205),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1207),
.B(n_237),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1194),
.A2(n_240),
.B(n_243),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1215),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1187),
.B(n_360),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1209),
.B(n_244),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1202),
.B(n_245),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1193),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1206),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1232),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1231),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1232),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1223),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1184),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1240),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1240),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1280),
.A2(n_1212),
.B1(n_1228),
.B2(n_1213),
.C(n_1196),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1248),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1248),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1266),
.A2(n_1227),
.B(n_1228),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1245),
.B(n_1254),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1238),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1238),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1243),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1266),
.A2(n_1229),
.B1(n_1219),
.B2(n_1218),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1260),
.A2(n_1263),
.B(n_1252),
.Y(n_1293)
);

OAI31xp33_ASAP7_75t_L g1294 ( 
.A1(n_1280),
.A2(n_1221),
.A3(n_1203),
.B(n_1236),
.Y(n_1294)
);

AOI33xp33_ASAP7_75t_L g1295 ( 
.A1(n_1263),
.A2(n_1237),
.A3(n_1216),
.B1(n_1226),
.B2(n_1230),
.B3(n_1198),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1249),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1278),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1254),
.B(n_1197),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1250),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1249),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1250),
.Y(n_1301)
);

OAI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1272),
.A2(n_1222),
.B1(n_1229),
.B2(n_250),
.C(n_252),
.Y(n_1302)
);

NOR4xp25_ASAP7_75t_SL g1303 ( 
.A(n_1277),
.B(n_246),
.C(n_249),
.D(n_254),
.Y(n_1303)
);

INVx5_ASAP7_75t_SL g1304 ( 
.A(n_1266),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1244),
.B(n_1267),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1289),
.B(n_1243),
.Y(n_1306)
);

NAND4xp25_ASAP7_75t_L g1307 ( 
.A(n_1287),
.B(n_1246),
.C(n_1255),
.D(n_1275),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1297),
.B(n_1288),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1293),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1297),
.B(n_1267),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1285),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1286),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1293),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1291),
.B(n_1277),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1304),
.B(n_1278),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1288),
.B(n_1267),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1305),
.B(n_1247),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1292),
.B(n_1279),
.C(n_1281),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1296),
.B(n_1279),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1305),
.B(n_1247),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1300),
.B(n_1281),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1282),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1283),
.Y(n_1323)
);

NAND2xp33_ASAP7_75t_L g1324 ( 
.A(n_1308),
.B(n_1264),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1311),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1308),
.B(n_1268),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1321),
.B(n_1312),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1322),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1319),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1310),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1323),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1306),
.B(n_1289),
.Y(n_1332)
);

NOR5xp2_ASAP7_75t_SL g1333 ( 
.A(n_1307),
.B(n_1304),
.C(n_1302),
.D(n_1265),
.E(n_1241),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1309),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1325),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1328),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_R g1337 ( 
.A(n_1324),
.B(n_1276),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1331),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1327),
.B(n_1318),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1326),
.B(n_1316),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1330),
.B(n_1317),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1284),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1332),
.B(n_1317),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1333),
.A2(n_1304),
.B1(n_1258),
.B2(n_1294),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1329),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1327),
.B(n_1314),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1334),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1334),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1326),
.B(n_1320),
.Y(n_1349)
);

OAI211xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1342),
.A2(n_1295),
.B(n_1299),
.C(n_1301),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1339),
.B(n_1299),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1352)
);

OAI21xp33_ASAP7_75t_L g1353 ( 
.A1(n_1344),
.A2(n_1295),
.B(n_1301),
.Y(n_1353)
);

AOI31xp33_ASAP7_75t_L g1354 ( 
.A1(n_1344),
.A2(n_1315),
.A3(n_1274),
.B(n_1268),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1347),
.A2(n_1269),
.B(n_1270),
.C(n_1259),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1346),
.B(n_1276),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1338),
.Y(n_1357)
);

AOI21xp33_ASAP7_75t_L g1358 ( 
.A1(n_1335),
.A2(n_1293),
.B(n_1259),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1356),
.Y(n_1359)
);

AOI21xp33_ASAP7_75t_L g1360 ( 
.A1(n_1355),
.A2(n_1353),
.B(n_1357),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1350),
.A2(n_1304),
.B1(n_1348),
.B2(n_1298),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1352),
.B(n_1340),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1354),
.A2(n_1348),
.B(n_1345),
.C(n_1273),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1351),
.A2(n_1341),
.B(n_1345),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1358),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1359),
.B(n_1337),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1362),
.Y(n_1367)
);

OAI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1361),
.A2(n_1313),
.B1(n_1309),
.B2(n_1261),
.C(n_1262),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1360),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1364),
.B(n_1349),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1365),
.A2(n_1298),
.B1(n_1273),
.B2(n_1257),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1363),
.A2(n_1337),
.B(n_1340),
.Y(n_1372)
);

AND4x1_ASAP7_75t_L g1373 ( 
.A(n_1367),
.B(n_1274),
.C(n_1343),
.D(n_1320),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1369),
.B(n_1370),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1366),
.A2(n_1303),
.B(n_1313),
.Y(n_1375)
);

NOR4xp25_ASAP7_75t_L g1376 ( 
.A(n_1368),
.B(n_1372),
.C(n_1371),
.D(n_1239),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1369),
.A2(n_1262),
.B(n_1261),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1367),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1369),
.B(n_1290),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1367),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1367),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_SL g1382 ( 
.A(n_1374),
.B(n_1257),
.C(n_1275),
.Y(n_1382)
);

NOR3xp33_ASAP7_75t_L g1383 ( 
.A(n_1379),
.B(n_1256),
.C(n_1252),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1376),
.A2(n_1256),
.B1(n_1253),
.B2(n_1271),
.C(n_1260),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1377),
.A2(n_1256),
.B1(n_1253),
.B2(n_1271),
.C(n_1251),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1377),
.A2(n_1253),
.B1(n_1251),
.B2(n_1242),
.C(n_1290),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1375),
.A2(n_1253),
.B1(n_1244),
.B2(n_259),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1381),
.A2(n_1253),
.B1(n_258),
.B2(n_260),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1378),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1389),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1382),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1388),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1383),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1387),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1386),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1384),
.Y(n_1396)
);

NAND4xp25_ASAP7_75t_SL g1397 ( 
.A(n_1385),
.B(n_1380),
.C(n_1373),
.D(n_262),
.Y(n_1397)
);

NAND4xp75_ASAP7_75t_L g1398 ( 
.A(n_1392),
.B(n_257),
.C(n_261),
.D(n_263),
.Y(n_1398)
);

NOR3xp33_ASAP7_75t_L g1399 ( 
.A(n_1397),
.B(n_1394),
.C(n_1396),
.Y(n_1399)
);

NOR2x1_ASAP7_75t_L g1400 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_SL g1401 ( 
.A(n_1393),
.B(n_264),
.C(n_269),
.Y(n_1401)
);

AND2x2_ASAP7_75t_SL g1402 ( 
.A(n_1395),
.B(n_271),
.Y(n_1402)
);

AOI31xp33_ASAP7_75t_L g1403 ( 
.A1(n_1396),
.A2(n_272),
.A3(n_274),
.B(n_275),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1390),
.Y(n_1404)
);

XOR2x1_ASAP7_75t_L g1405 ( 
.A(n_1404),
.B(n_276),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1398),
.Y(n_1406)
);

NOR4xp25_ASAP7_75t_L g1407 ( 
.A(n_1400),
.B(n_278),
.C(n_279),
.D(n_283),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1402),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1403),
.B(n_293),
.Y(n_1409)
);

NAND5xp2_ASAP7_75t_L g1410 ( 
.A(n_1399),
.B(n_294),
.C(n_297),
.D(n_298),
.E(n_300),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1401),
.B(n_301),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1406),
.B(n_302),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1405),
.Y(n_1413)
);

NOR2x1_ASAP7_75t_L g1414 ( 
.A(n_1410),
.B(n_303),
.Y(n_1414)
);

AOI22x1_ASAP7_75t_L g1415 ( 
.A1(n_1413),
.A2(n_1409),
.B1(n_1407),
.B2(n_1408),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1412),
.B(n_1411),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1414),
.B(n_351),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1416),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1417),
.Y(n_1419)
);

XNOR2xp5_ASAP7_75t_L g1420 ( 
.A(n_1418),
.B(n_1415),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1419),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1420),
.B(n_306),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1421),
.A2(n_307),
.B1(n_312),
.B2(n_313),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1422),
.A2(n_315),
.B1(n_316),
.B2(n_319),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_R g1425 ( 
.A1(n_1424),
.A2(n_1423),
.B1(n_327),
.B2(n_328),
.C(n_329),
.Y(n_1425)
);

OAI221xp5_ASAP7_75t_R g1426 ( 
.A1(n_1425),
.A2(n_325),
.B1(n_332),
.B2(n_334),
.C(n_335),
.Y(n_1426)
);

AOI211xp5_ASAP7_75t_L g1427 ( 
.A1(n_1426),
.A2(n_338),
.B(n_339),
.C(n_340),
.Y(n_1427)
);


endmodule