module fake_jpeg_9557_n_175 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_34),
.Y(n_48)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_20),
.B1(n_29),
.B2(n_18),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_24),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_60),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_63),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_30),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_30),
.B(n_33),
.C(n_35),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_73),
.B1(n_25),
.B2(n_26),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_45),
.B(n_51),
.C(n_40),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_75),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_82),
.B(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_35),
.C(n_49),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_58),
.C(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_43),
.B1(n_54),
.B2(n_32),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_90),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_54),
.B1(n_38),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_38),
.B1(n_26),
.B2(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_1),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_67),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_14),
.B(n_37),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_38),
.B1(n_14),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_64),
.B1(n_59),
.B2(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_79),
.C(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_76),
.B1(n_85),
.B2(n_80),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_86),
.B1(n_78),
.B2(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_37),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_119),
.C(n_120),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_118),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_82),
.B(n_2),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_82),
.C(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_99),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_1),
.B(n_3),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_101),
.C(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_109),
.C(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_138),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_124),
.B1(n_112),
.B2(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_108),
.C(n_100),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_108),
.C(n_94),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_114),
.B1(n_118),
.B2(n_115),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_136),
.A2(n_119),
.B1(n_123),
.B2(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_127),
.B1(n_130),
.B2(n_116),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_6),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_64),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_107),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_131),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_1),
.B(n_4),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_135),
.C(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_155),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_13),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_12),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_9),
.C(n_11),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_156),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_156),
.B(n_146),
.Y(n_159)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_8),
.B1(n_139),
.B2(n_148),
.C(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_154),
.C(n_162),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_140),
.C(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_142),
.B1(n_147),
.B2(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_157),
.C(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_167),
.B(n_8),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_8),
.Y(n_175)
);


endmodule