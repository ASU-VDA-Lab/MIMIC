module fake_jpeg_3462_n_650 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_441;
wire n_161;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_0),
.B(n_3),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_6),
.B(n_17),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_59),
.B(n_75),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

INVx2_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_64),
.B(n_23),
.Y(n_154)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_17),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_67),
.Y(n_152)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_70),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_72),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_73),
.Y(n_184)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_76),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_77),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_78),
.B(n_79),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_18),
.B(n_17),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_97),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_19),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_24),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_101),
.B(n_127),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_103),
.Y(n_185)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_111),
.Y(n_189)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_20),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_138),
.B(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_140),
.B(n_15),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_145),
.B(n_150),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_154),
.B(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_59),
.B(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_171),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_168),
.B(n_172),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_170),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_93),
.B(n_22),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_74),
.B(n_22),
.Y(n_172)
);

OR2x4_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_27),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_173),
.A2(n_30),
.B(n_48),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_54),
.B1(n_57),
.B2(n_28),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g255 ( 
.A1(n_174),
.A2(n_119),
.B1(n_117),
.B2(n_116),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_60),
.B(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_221),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_61),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_198),
.Y(n_231)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_191),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_69),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_70),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_211),
.Y(n_257)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_200),
.Y(n_293)
);

INVx6_ASAP7_75t_SL g203 ( 
.A(n_129),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g290 ( 
.A(n_203),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_102),
.A2(n_54),
.B1(n_57),
.B2(n_21),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_205),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_90),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_20),
.B1(n_53),
.B2(n_52),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_42),
.B1(n_28),
.B2(n_35),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_130),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_98),
.B(n_21),
.C(n_53),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_215),
.B(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_73),
.B(n_56),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_115),
.B(n_56),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_194),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_226),
.B(n_229),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_201),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_233),
.B(n_235),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_144),
.B(n_36),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_237),
.Y(n_361)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_156),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_240),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_241),
.Y(n_355)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_135),
.Y(n_242)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_154),
.A2(n_36),
.B1(n_42),
.B2(n_47),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_243),
.A2(n_255),
.B1(n_262),
.B2(n_301),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_244),
.A2(n_250),
.B1(n_254),
.B2(n_281),
.Y(n_332)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_148),
.Y(n_245)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_153),
.Y(n_249)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_249),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_146),
.A2(n_109),
.B1(n_108),
.B2(n_91),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_147),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_252),
.Y(n_347)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_77),
.B1(n_99),
.B2(n_95),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

CKINVDCx6p67_ASAP7_75t_R g324 ( 
.A(n_260),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_147),
.A2(n_52),
.B1(n_47),
.B2(n_45),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_263),
.B(n_305),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_264),
.B(n_270),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_144),
.B(n_45),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_279),
.Y(n_312)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_136),
.Y(n_267)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_269),
.B(n_282),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_178),
.B(n_30),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_149),
.B(n_218),
.Y(n_321)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_273),
.B(n_278),
.Y(n_344)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_139),
.Y(n_274)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_133),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_276),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_146),
.A2(n_94),
.B1(n_48),
.B2(n_16),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_277),
.A2(n_283),
.B1(n_284),
.B2(n_294),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_137),
.B(n_16),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_152),
.B(n_15),
.Y(n_279)
);

AOI22x1_ASAP7_75t_SL g281 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_208),
.B(n_1),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_155),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_195),
.Y(n_285)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_166),
.B(n_177),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_286),
.B(n_298),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_167),
.B(n_7),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_152),
.Y(n_291)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_189),
.Y(n_292)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_176),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_174),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_295),
.A2(n_302),
.B1(n_303),
.B2(n_238),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_143),
.B(n_10),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_132),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_223),
.A2(n_13),
.B1(n_192),
.B2(n_163),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_184),
.A2(n_13),
.B1(n_186),
.B2(n_196),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_157),
.A2(n_13),
.B1(n_142),
.B2(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_212),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_189),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_193),
.B(n_224),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_186),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_232),
.B(n_219),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_311),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_252),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_206),
.B1(n_218),
.B2(n_216),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_313),
.A2(n_360),
.B1(n_290),
.B2(n_284),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_320),
.B(n_336),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_321),
.B(n_255),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_162),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_327),
.B(n_356),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_265),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_225),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_357),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_277),
.B(n_149),
.CI(n_181),
.CON(n_342),
.SN(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_238),
.B(n_281),
.C(n_257),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_231),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_345),
.B(n_351),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_240),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_202),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_227),
.B(n_131),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_269),
.B(n_132),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_230),
.B(n_197),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_292),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_254),
.A2(n_216),
.B1(n_206),
.B2(n_196),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_180),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_290),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_303),
.B(n_301),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_368),
.A2(n_378),
.B(n_398),
.Y(n_434)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_308),
.Y(n_371)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_371),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_372),
.A2(n_387),
.B1(n_399),
.B2(n_331),
.Y(n_442)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_350),
.A2(n_354),
.B1(n_321),
.B2(n_310),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_411),
.B1(n_318),
.B2(n_358),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_347),
.A2(n_287),
.B(n_255),
.Y(n_378)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_346),
.Y(n_380)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_381),
.B(n_406),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_290),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_382),
.B(n_391),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_384),
.A2(n_385),
.B(n_400),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_329),
.A2(n_243),
.B(n_241),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_332),
.A2(n_283),
.B1(n_294),
.B2(n_248),
.Y(n_387)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_389),
.Y(n_417)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_275),
.B1(n_239),
.B2(n_306),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_331),
.B1(n_361),
.B2(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g394 ( 
.A(n_329),
.B(n_234),
.C(n_280),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_394),
.B(n_409),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_395),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_274),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_401),
.Y(n_421)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_397),
.A2(n_402),
.B1(n_403),
.B2(n_405),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_287),
.B(n_300),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_245),
.B1(n_267),
.B2(n_214),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_357),
.B(n_300),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_312),
.B(n_261),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_404),
.A2(n_343),
.B1(n_324),
.B2(n_330),
.Y(n_444)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_315),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_309),
.B(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_407),
.A2(n_412),
.B1(n_355),
.B2(n_353),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_410),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_293),
.C(n_228),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_311),
.A2(n_225),
.B1(n_169),
.B2(n_197),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_340),
.B(n_169),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_413),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_414),
.A2(n_419),
.B1(n_420),
.B2(n_423),
.Y(n_464)
);

AOI32xp33_ASAP7_75t_L g415 ( 
.A1(n_377),
.A2(n_342),
.A3(n_366),
.B1(n_339),
.B2(n_344),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_342),
.B1(n_334),
.B2(n_361),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_416),
.A2(n_426),
.B1(n_430),
.B2(n_432),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_367),
.B1(n_378),
.B2(n_383),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_404),
.A2(n_317),
.B1(n_319),
.B2(n_242),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_328),
.Y(n_425)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_425),
.A2(n_437),
.B(n_443),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_319),
.B1(n_349),
.B2(n_338),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_381),
.A2(n_328),
.B(n_325),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_429),
.B(n_425),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_392),
.A2(n_349),
.B1(n_338),
.B2(n_325),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_368),
.A2(n_365),
.B1(n_362),
.B2(n_326),
.Y(n_432)
);

AO21x2_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_324),
.B(n_362),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_398),
.A2(n_324),
.B(n_330),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_438),
.A2(n_446),
.B(n_413),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_442),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_388),
.B(n_370),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_444),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_383),
.A2(n_365),
.B(n_326),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_355),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_448),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_483),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_394),
.C(n_409),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_486),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_421),
.B(n_369),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_455),
.B(n_459),
.Y(n_513)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_427),
.Y(n_456)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_458),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_451),
.B(n_405),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_428),
.Y(n_461)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_466),
.A2(n_476),
.B(n_434),
.Y(n_493)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_467),
.Y(n_507)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_307),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_470),
.B(n_475),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_414),
.A2(n_413),
.B1(n_386),
.B2(n_371),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_471),
.A2(n_473),
.B1(n_487),
.B2(n_430),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_447),
.B(n_451),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_477),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_420),
.A2(n_411),
.B1(n_386),
.B2(n_373),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_447),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_375),
.B(n_389),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_443),
.B(n_390),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_478),
.B(n_488),
.Y(n_518)
);

INVx13_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_479),
.Y(n_489)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_480),
.Y(n_519)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_446),
.B(n_403),
.CI(n_391),
.CON(n_481),
.SN(n_481)
);

FAx1_ASAP7_75t_SL g521 ( 
.A(n_481),
.B(n_417),
.CI(n_422),
.CON(n_521),
.SN(n_521)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

AND2x2_ASAP7_75t_SL g484 ( 
.A(n_418),
.B(n_397),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_484),
.Y(n_492)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_435),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_440),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_380),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_429),
.A2(n_374),
.B1(n_395),
.B2(n_337),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_307),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_493),
.A2(n_501),
.B(n_509),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_517),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_464),
.A2(n_465),
.B1(n_471),
.B2(n_453),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_495),
.A2(n_498),
.B1(n_502),
.B2(n_505),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_464),
.A2(n_416),
.B1(n_425),
.B2(n_437),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_497),
.A2(n_483),
.B1(n_482),
.B2(n_481),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_429),
.B1(n_423),
.B2(n_437),
.Y(n_498)
);

FAx1_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_418),
.CI(n_437),
.CON(n_501),
.SN(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_468),
.A2(n_437),
.B1(n_432),
.B2(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_445),
.Y(n_504)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_466),
.A2(n_437),
.B1(n_445),
.B2(n_419),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_441),
.Y(n_508)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_508),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_474),
.A2(n_444),
.B(n_440),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_510),
.A2(n_480),
.B1(n_463),
.B2(n_439),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_486),
.B(n_441),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_512),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_469),
.B(n_454),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_515),
.B(n_253),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_410),
.Y(n_516)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_474),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_433),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_467),
.B(n_436),
.Y(n_522)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_522),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_462),
.C(n_484),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_538),
.C(n_519),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_495),
.A2(n_487),
.B1(n_484),
.B2(n_462),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_526),
.A2(n_542),
.B1(n_546),
.B2(n_506),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g564 ( 
.A(n_528),
.B(n_539),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_474),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_544),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_530),
.A2(n_531),
.B1(n_540),
.B2(n_501),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_497),
.A2(n_482),
.B1(n_476),
.B2(n_481),
.Y(n_531)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_537),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_484),
.C(n_457),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_499),
.B(n_456),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_498),
.A2(n_461),
.B1(n_460),
.B2(n_485),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_499),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_541),
.B(n_550),
.Y(n_572)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_491),
.Y(n_543)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_543),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_511),
.B(n_431),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_545),
.A2(n_505),
.B(n_501),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_490),
.A2(n_439),
.B1(n_431),
.B2(n_433),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_547),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_489),
.B(n_436),
.Y(n_548)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_548),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_511),
.B(n_479),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_549),
.B(n_553),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_490),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_520),
.A2(n_479),
.B1(n_379),
.B2(n_337),
.Y(n_551)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_551),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_149),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_552),
.B(n_494),
.Y(n_565)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_556),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_527),
.A2(n_517),
.B(n_493),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_557),
.A2(n_571),
.B(n_521),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_559),
.A2(n_532),
.B1(n_526),
.B2(n_545),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_548),
.B(n_489),
.Y(n_562)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_562),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_502),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_568),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_552),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_547),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_566),
.B(n_534),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_544),
.B(n_519),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_524),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_569),
.A2(n_573),
.B1(n_576),
.B2(n_533),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_575),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_527),
.A2(n_492),
.B(n_518),
.C(n_521),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

XOR2x1_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_492),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_572),
.B(n_513),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_578),
.B(n_579),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_570),
.B(n_528),
.C(n_525),
.Y(n_579)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_580),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_538),
.C(n_535),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_582),
.B(n_588),
.Y(n_610)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_583),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_586),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_561),
.A2(n_540),
.B1(n_530),
.B2(n_531),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_555),
.B(n_536),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_589),
.B(n_592),
.C(n_594),
.Y(n_600)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_555),
.Y(n_590)
);

BUFx24_ASAP7_75t_SL g605 ( 
.A(n_590),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_561),
.A2(n_518),
.B1(n_523),
.B2(n_503),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_573),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_539),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_593),
.A2(n_571),
.B(n_569),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_559),
.B(n_546),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_564),
.B(n_506),
.C(n_503),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_565),
.C(n_560),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_563),
.C(n_568),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_597),
.B(n_598),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_563),
.C(n_576),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_585),
.B(n_557),
.C(n_564),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_599),
.B(n_604),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_601),
.A2(n_606),
.B(n_587),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_603),
.B(n_507),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g606 ( 
.A1(n_577),
.A2(n_562),
.B(n_556),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_582),
.B(n_575),
.C(n_560),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_607),
.B(n_609),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_581),
.A2(n_554),
.B1(n_558),
.B2(n_500),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_611),
.A2(n_583),
.B1(n_593),
.B2(n_595),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_615),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_614),
.A2(n_622),
.B(n_276),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_597),
.B(n_587),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_596),
.A2(n_554),
.B1(n_500),
.B2(n_496),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_617),
.B(n_618),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_601),
.A2(n_600),
.B1(n_610),
.B2(n_602),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_586),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_620),
.B(n_621),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_598),
.B(n_496),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_601),
.A2(n_507),
.B(n_258),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_623),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_599),
.A2(n_272),
.B1(n_236),
.B2(n_296),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_624),
.B(n_256),
.Y(n_625)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_625),
.Y(n_634)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_626),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_614),
.A2(n_605),
.B1(n_268),
.B2(n_259),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_627),
.B(n_629),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_260),
.C(n_160),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_621),
.B(n_160),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g636 ( 
.A(n_631),
.B(n_620),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_630),
.B(n_615),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_636),
.Y(n_641)
);

OAI221xp5_ASAP7_75t_L g639 ( 
.A1(n_628),
.A2(n_619),
.B1(n_613),
.B2(n_622),
.C(n_260),
.Y(n_639)
);

AOI31xp33_ASAP7_75t_L g642 ( 
.A1(n_639),
.A2(n_629),
.A3(n_626),
.B(n_627),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_638),
.A2(n_632),
.B(n_633),
.Y(n_640)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_640),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_642),
.B(n_643),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_637),
.B(n_160),
.C(n_161),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_644),
.A2(n_641),
.B(n_645),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_646),
.B(n_634),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_207),
.B1(n_161),
.B2(n_180),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_161),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_133),
.B(n_180),
.Y(n_650)
);


endmodule