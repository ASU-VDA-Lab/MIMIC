module fake_jpeg_10590_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_1),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_7),
.A2(n_1),
.B(n_2),
.Y(n_12)
);

NAND2x1_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_16),
.Y(n_20)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_8),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_15)
);

CKINVDCx11_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_5),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_6),
.B(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_21),
.B(n_17),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_20),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_13),
.C(n_20),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_22),
.B(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_27)
);


endmodule