module fake_jpeg_22886_n_229 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_37),
.B(n_15),
.C(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_28),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_53),
.B1(n_56),
.B2(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_27),
.B1(n_18),
.B2(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_70),
.B1(n_71),
.B2(n_51),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_37),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_67),
.B(n_76),
.C(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_40),
.A2(n_33),
.B1(n_31),
.B2(n_38),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_33),
.B1(n_15),
.B2(n_34),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_0),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_68),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_51),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_87),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_54),
.B1(n_43),
.B2(n_65),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_49),
.B1(n_41),
.B2(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_74),
.B1(n_56),
.B2(n_46),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_101),
.B1(n_113),
.B2(n_117),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_105),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_59),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_57),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.C(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_41),
.B1(n_48),
.B2(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_65),
.B1(n_54),
.B2(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_91),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_22),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_43),
.B1(n_55),
.B2(n_38),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_31),
.C(n_52),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_92),
.C(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_128),
.B1(n_137),
.B2(n_25),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_79),
.B(n_84),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_138),
.B(n_116),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_125),
.C(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_84),
.B1(n_85),
.B2(n_95),
.Y(n_128)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_85),
.B1(n_47),
.B2(n_52),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_61),
.B(n_35),
.C(n_23),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_78),
.B1(n_81),
.B2(n_28),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_133),
.B1(n_104),
.B2(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_78),
.B1(n_47),
.B2(n_61),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_140),
.B(n_152),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_138),
.B1(n_120),
.B2(n_35),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_145),
.B1(n_148),
.B2(n_157),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_16),
.B1(n_24),
.B2(n_17),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_24),
.B1(n_21),
.B2(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_24),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_125),
.C(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_135),
.B1(n_119),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_25),
.B1(n_23),
.B2(n_20),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_172),
.C(n_173),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_141),
.B(n_157),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_153),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_165),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_20),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_122),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_25),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_23),
.C(n_20),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_23),
.C(n_20),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_1),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_181),
.C(n_174),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_177),
.B(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_172),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_144),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_147),
.B1(n_141),
.B2(n_156),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_168),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_141),
.B1(n_151),
.B2(n_145),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_162),
.B1(n_173),
.B2(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_168),
.B1(n_160),
.B2(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_175),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_167),
.C(n_2),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_197),
.C(n_184),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_7),
.B(n_12),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_185),
.B1(n_184),
.B2(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_189),
.B1(n_3),
.B2(n_5),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.C(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_1),
.C(n_2),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_196),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_212),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_195),
.B(n_188),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_193),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_206),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_197),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_213),
.B(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_217),
.B(n_202),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_204),
.Y(n_217)
);

OAI321xp33_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_222),
.A3(n_9),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_189),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_SL g225 ( 
.A1(n_223),
.A2(n_224),
.A3(n_11),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_220),
.C(n_221),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_10),
.B(n_11),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_11),
.B(n_13),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_3),
.B(n_225),
.C(n_209),
.Y(n_229)
);


endmodule