module real_aes_1119_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_0), .B(n_123), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_1), .A2(n_117), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_2), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_3), .B(n_123), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_4), .B(n_134), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_5), .B(n_134), .Y(n_209) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_7), .B(n_134), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_8), .Y(n_734) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_9), .B(n_132), .Y(n_185) );
AND2x2_ASAP7_75t_L g442 ( .A(n_10), .B(n_179), .Y(n_442) );
AND2x2_ASAP7_75t_L g450 ( .A(n_11), .B(n_146), .Y(n_450) );
INVx2_ASAP7_75t_L g114 ( .A(n_12), .Y(n_114) );
AOI221x1_ASAP7_75t_L g116 ( .A1(n_13), .A2(n_25), .B1(n_117), .B2(n_123), .C(n_130), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_14), .B(n_134), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g412 ( .A(n_15), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_16), .B(n_123), .Y(n_181) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_179), .B(n_180), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_18), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_19), .B(n_112), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_20), .B(n_134), .Y(n_193) );
AO21x1_ASAP7_75t_L g204 ( .A1(n_21), .A2(n_123), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_22), .B(n_123), .Y(n_481) );
INVx1_ASAP7_75t_L g416 ( .A(n_23), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_24), .A2(n_87), .B1(n_123), .B2(n_511), .Y(n_510) );
NAND2x1_ASAP7_75t_L g142 ( .A(n_26), .B(n_134), .Y(n_142) );
NAND2x1_ASAP7_75t_L g172 ( .A(n_27), .B(n_132), .Y(n_172) );
OR2x2_ASAP7_75t_L g115 ( .A(n_28), .B(n_84), .Y(n_115) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_28), .A2(n_84), .B(n_114), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_29), .B(n_132), .Y(n_167) );
AOI221xp5_ASAP7_75t_L g100 ( .A1(n_30), .A2(n_101), .B1(n_720), .B2(n_723), .C(n_724), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_30), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_31), .B(n_134), .Y(n_184) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_32), .A2(n_146), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_33), .B(n_132), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_34), .A2(n_117), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_35), .B(n_134), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_36), .A2(n_117), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g118 ( .A(n_37), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g129 ( .A(n_37), .B(n_122), .Y(n_129) );
INVx1_ASAP7_75t_L g519 ( .A(n_37), .Y(n_519) );
OR2x6_ASAP7_75t_L g414 ( .A(n_38), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_39), .B(n_123), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_40), .B(n_123), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_41), .B(n_134), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_42), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_43), .B(n_132), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_44), .B(n_123), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_45), .A2(n_117), .B(n_446), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_46), .A2(n_117), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_47), .B(n_132), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_48), .B(n_132), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_49), .B(n_123), .Y(n_455) );
INVx1_ASAP7_75t_L g121 ( .A(n_50), .Y(n_121) );
INVx1_ASAP7_75t_L g126 ( .A(n_50), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_51), .B(n_134), .Y(n_448) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_52), .A2(n_99), .B1(n_727), .B2(n_738), .C1(n_746), .C2(n_750), .Y(n_98) );
OAI22xp33_ASAP7_75t_SL g740 ( .A1(n_52), .A2(n_418), .B1(n_419), .B2(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_52), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_53), .Y(n_725) );
AND2x2_ASAP7_75t_L g472 ( .A(n_54), .B(n_112), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_55), .B(n_132), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_56), .B(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_57), .B(n_132), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_58), .A2(n_117), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_59), .B(n_123), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_60), .B(n_123), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_61), .A2(n_117), .B(n_463), .Y(n_462) );
AO21x1_ASAP7_75t_L g206 ( .A1(n_62), .A2(n_117), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g487 ( .A(n_63), .B(n_113), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_64), .B(n_123), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_65), .B(n_132), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_66), .B(n_123), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_67), .B(n_132), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_68), .A2(n_92), .B1(n_117), .B2(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g157 ( .A(n_69), .B(n_113), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_70), .B(n_134), .Y(n_484) );
INVx1_ASAP7_75t_L g119 ( .A(n_71), .Y(n_119) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
AND2x2_ASAP7_75t_L g176 ( .A(n_72), .B(n_146), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_73), .B(n_132), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_74), .A2(n_117), .B(n_476), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_75), .A2(n_117), .B(n_429), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_76), .A2(n_117), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g467 ( .A(n_77), .B(n_113), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_78), .B(n_112), .Y(n_508) );
INVx1_ASAP7_75t_L g417 ( .A(n_79), .Y(n_417) );
AND2x2_ASAP7_75t_L g161 ( .A(n_80), .B(n_146), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_81), .B(n_123), .Y(n_195) );
AND2x2_ASAP7_75t_L g432 ( .A(n_82), .B(n_179), .Y(n_432) );
AND2x2_ASAP7_75t_L g205 ( .A(n_83), .B(n_186), .Y(n_205) );
AND2x2_ASAP7_75t_L g149 ( .A(n_85), .B(n_146), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_86), .B(n_132), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_88), .B(n_134), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_89), .B(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_90), .A2(n_117), .B(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_91), .A2(n_117), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_93), .B(n_134), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_94), .B(n_134), .Y(n_166) );
BUFx2_ASAP7_75t_L g486 ( .A(n_95), .Y(n_486) );
BUFx2_ASAP7_75t_L g735 ( .A(n_96), .Y(n_735) );
BUFx2_ASAP7_75t_SL g754 ( .A(n_96), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_97), .A2(n_117), .B(n_183), .Y(n_182) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_409), .B1(n_418), .B2(n_718), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_103), .A2(n_411), .B1(n_419), .B2(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_321), .Y(n_103) );
AND4x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_233), .C(n_260), .D(n_295), .Y(n_104) );
AOI221xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_158), .B1(n_198), .B2(n_213), .C(n_217), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_137), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_108), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g274 ( .A(n_109), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g329 ( .A(n_109), .B(n_284), .Y(n_329) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g232 ( .A(n_110), .B(n_150), .Y(n_232) );
AND2x4_ASAP7_75t_L g268 ( .A(n_110), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_110), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g199 ( .A(n_111), .Y(n_199) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_111), .Y(n_371) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_136), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_112), .A2(n_163), .B(n_164), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_112), .Y(n_175) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_112), .A2(n_116), .B(n_136), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_112), .A2(n_427), .B(n_428), .Y(n_426) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_112), .A2(n_510), .B(n_516), .Y(n_509) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x4_ASAP7_75t_L g186 ( .A(n_114), .B(n_115), .Y(n_186) );
AND2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
BUFx3_ASAP7_75t_L g515 ( .A(n_118), .Y(n_515) );
AND2x6_ASAP7_75t_L g132 ( .A(n_119), .B(n_125), .Y(n_132) );
INVx2_ASAP7_75t_L g521 ( .A(n_119), .Y(n_521) );
AND2x4_ASAP7_75t_L g517 ( .A(n_120), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g134 ( .A(n_121), .B(n_127), .Y(n_134) );
INVx2_ASAP7_75t_L g513 ( .A(n_121), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_122), .Y(n_514) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_135), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_132), .B(n_486), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_135), .A2(n_142), .B(n_143), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_135), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_135), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_135), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_135), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_135), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_135), .A2(n_430), .B(n_431), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_135), .A2(n_439), .B(n_440), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_135), .A2(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_135), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_135), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_135), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_135), .A2(n_484), .B(n_485), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_SL g226 ( .A1(n_137), .A2(n_199), .B(n_227), .C(n_231), .Y(n_226) );
AND2x2_ASAP7_75t_L g247 ( .A(n_137), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_137), .B(n_199), .Y(n_387) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_150), .Y(n_137) );
INVx2_ASAP7_75t_L g267 ( .A(n_138), .Y(n_267) );
BUFx3_ASAP7_75t_L g283 ( .A(n_138), .Y(n_283) );
INVxp67_ASAP7_75t_L g287 ( .A(n_138), .Y(n_287) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_149), .Y(n_138) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_139), .A2(n_145), .B(n_149), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_145), .A2(n_151), .B(n_157), .Y(n_150) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_145), .A2(n_151), .B(n_157), .Y(n_212) );
AO21x1_ASAP7_75t_SL g460 ( .A1(n_145), .A2(n_461), .B(n_467), .Y(n_460) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_145), .A2(n_461), .B(n_467), .Y(n_494) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_147), .A2(n_444), .B(n_450), .Y(n_443) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx4f_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx2_ASAP7_75t_L g266 ( .A(n_150), .Y(n_266) );
AND2x2_ASAP7_75t_L g272 ( .A(n_150), .B(n_245), .Y(n_272) );
AND2x2_ASAP7_75t_L g298 ( .A(n_150), .B(n_267), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_152), .B(n_156), .Y(n_151) );
AOI211xp5_ASAP7_75t_L g295 ( .A1(n_158), .A2(n_296), .B(n_299), .C(n_309), .Y(n_295) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_177), .Y(n_158) );
OAI321xp33_ASAP7_75t_L g270 ( .A1(n_159), .A2(n_218), .A3(n_271), .B1(n_273), .B2(n_274), .C(n_276), .Y(n_270) );
AND2x2_ASAP7_75t_L g391 ( .A(n_159), .B(n_366), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_159), .Y(n_394) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_168), .Y(n_159) );
INVx5_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_160), .B(n_230), .Y(n_229) );
NOR2x1_ASAP7_75t_SL g261 ( .A(n_160), .B(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g306 ( .A(n_160), .Y(n_306) );
AND2x2_ASAP7_75t_L g408 ( .A(n_160), .B(n_178), .Y(n_408) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g215 ( .A(n_168), .B(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_168), .Y(n_225) );
INVx4_ASAP7_75t_L g230 ( .A(n_168), .Y(n_230) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_175), .B(n_176), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AOI21x1_ASAP7_75t_L g435 ( .A1(n_175), .A2(n_436), .B(n_442), .Y(n_435) );
INVx1_ASAP7_75t_L g273 ( .A(n_177), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_R g376 ( .A1(n_177), .A2(n_215), .B(n_247), .C(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g396 ( .A(n_177), .B(n_221), .Y(n_396) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_187), .Y(n_177) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
INVx2_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
OR2x2_ASAP7_75t_L g239 ( .A(n_178), .B(n_230), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_178), .B(n_262), .Y(n_308) );
BUFx3_ASAP7_75t_L g315 ( .A(n_178), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_179), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_186), .Y(n_180) );
INVx1_ASAP7_75t_SL g189 ( .A(n_186), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_186), .B(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_186), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_186), .A2(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g278 ( .A(n_187), .Y(n_278) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_187), .Y(n_291) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
INVx1_ASAP7_75t_L g333 ( .A(n_188), .Y(n_333) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_196), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_189), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_189), .A2(n_190), .B(n_196), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_195), .Y(n_190) );
AND2x2_ASAP7_75t_L g234 ( .A(n_198), .B(n_235), .Y(n_234) );
OAI31xp33_ASAP7_75t_L g385 ( .A1(n_198), .A2(n_386), .A3(n_388), .B(n_391), .Y(n_385) );
INVx1_ASAP7_75t_SL g403 ( .A(n_198), .Y(n_403) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AOI21xp33_ASAP7_75t_L g217 ( .A1(n_199), .A2(n_218), .B(n_226), .Y(n_217) );
NAND2x1_ASAP7_75t_L g297 ( .A(n_199), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g326 ( .A(n_199), .Y(n_326) );
INVx2_ASAP7_75t_L g275 ( .A(n_200), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_200), .B(n_258), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_200), .B(n_257), .Y(n_367) );
NOR2xp33_ASAP7_75t_SL g375 ( .A(n_200), .B(n_326), .Y(n_375) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_201), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g255 ( .A(n_201), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g284 ( .A(n_201), .B(n_266), .Y(n_284) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g248 ( .A(n_202), .Y(n_248) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
OAI21x1_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_206), .B(n_210), .Y(n_203) );
INVx1_ASAP7_75t_L g211 ( .A(n_205), .Y(n_211) );
INVx2_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_212), .Y(n_316) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
AND2x2_ASAP7_75t_L g331 ( .A(n_214), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g242 ( .A(n_215), .B(n_236), .Y(n_242) );
INVx2_ASAP7_75t_SL g290 ( .A(n_215), .Y(n_290) );
INVx4_ASAP7_75t_L g221 ( .A(n_216), .Y(n_221) );
AND2x2_ASAP7_75t_L g319 ( .A(n_216), .B(n_262), .Y(n_319) );
AND2x2_ASAP7_75t_SL g337 ( .A(n_216), .B(n_332), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_216), .B(n_230), .Y(n_354) );
INVx1_ASAP7_75t_L g360 ( .A(n_218), .Y(n_360) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_222), .Y(n_218) );
INVx1_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
OR2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
OR2x2_ASAP7_75t_L g344 ( .A(n_220), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g374 ( .A(n_220), .B(n_262), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_221), .B(n_224), .Y(n_250) );
AND2x2_ASAP7_75t_L g342 ( .A(n_221), .B(n_332), .Y(n_342) );
AND2x4_ASAP7_75t_L g404 ( .A(n_221), .B(n_283), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
INVx2_ASAP7_75t_L g228 ( .A(n_223), .Y(n_228) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2xp67_ASAP7_75t_SL g227 ( .A(n_228), .B(n_229), .Y(n_227) );
OAI322xp33_ASAP7_75t_SL g240 ( .A1(n_228), .A2(n_241), .A3(n_243), .B1(n_246), .B2(n_249), .C1(n_251), .C2(n_253), .Y(n_240) );
INVx1_ASAP7_75t_L g398 ( .A(n_228), .Y(n_398) );
OR2x2_ASAP7_75t_L g251 ( .A(n_229), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g277 ( .A(n_230), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_230), .B(n_278), .Y(n_293) );
INVx2_ASAP7_75t_L g320 ( .A(n_230), .Y(n_320) );
AND2x4_ASAP7_75t_L g332 ( .A(n_230), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_SL g335 ( .A(n_232), .B(n_248), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_238), .B(n_240), .Y(n_233) );
AND2x2_ASAP7_75t_L g301 ( .A(n_235), .B(n_268), .Y(n_301) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_236), .B(n_390), .Y(n_389) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_237), .B(n_256), .Y(n_341) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g249 ( .A(n_239), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_242), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g377 ( .A(n_244), .B(n_341), .Y(n_377) );
NOR4xp25_ASAP7_75t_L g381 ( .A(n_244), .B(n_258), .C(n_298), .D(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g258 ( .A(n_245), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_269), .Y(n_294) );
AND2x4_ASAP7_75t_L g358 ( .A(n_245), .B(n_269), .Y(n_358) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_248), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
OR2x2_ASAP7_75t_L g347 ( .A(n_255), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g401 ( .A(n_255), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_256), .B(n_268), .Y(n_302) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AOI211xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_263), .B(n_270), .C(n_285), .Y(n_260) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_266), .B(n_269), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_267), .B(n_272), .Y(n_271) );
BUFx2_ASAP7_75t_L g349 ( .A(n_267), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g364 ( .A(n_268), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B(n_280), .Y(n_276) );
AND2x4_ASAP7_75t_L g313 ( .A(n_277), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g407 ( .A(n_277), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_SL g311 ( .A(n_283), .Y(n_311) );
AND2x2_ASAP7_75t_L g370 ( .A(n_284), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g384 ( .A(n_284), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_288), .B(n_292), .C(n_294), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_286), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g362 ( .A(n_287), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g383 ( .A(n_287), .B(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g372 ( .A(n_290), .B(n_314), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_293), .A2(n_300), .B1(n_302), .B2(n_303), .Y(n_299) );
INVx1_ASAP7_75t_SL g390 ( .A(n_294), .Y(n_390) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_305), .B(n_314), .Y(n_356) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_308), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_316), .B2(n_317), .Y(n_309) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_SL g323 ( .A1(n_314), .A2(n_324), .B(n_327), .Y(n_323) );
AND2x2_ASAP7_75t_L g352 ( .A(n_314), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND3x2_ASAP7_75t_L g318 ( .A(n_315), .B(n_319), .C(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g380 ( .A(n_315), .B(n_337), .Y(n_380) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_366), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_322), .B(n_378), .Y(n_321) );
NAND4xp25_ASAP7_75t_L g322 ( .A(n_323), .B(n_338), .C(n_359), .D(n_376), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_334), .B2(n_336), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_330), .A2(n_344), .B1(n_364), .B2(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_334), .A2(n_357), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_343), .B2(n_346), .C(n_350), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_356), .B2(n_357), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_353), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_353), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_365), .B2(n_367), .C(n_368), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_364), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_373), .B2(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_374), .A2(n_394), .B(n_395), .C(n_397), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_385), .C(n_392), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_399), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_392) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
CKINVDCx11_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
OR2x6_ASAP7_75t_SL g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x6_ASAP7_75t_SL g719 ( .A(n_412), .B(n_414), .Y(n_719) );
OR2x2_ASAP7_75t_L g726 ( .A(n_412), .B(n_414), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_412), .B(n_413), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx4_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_626), .Y(n_419) );
NOR3xp33_ASAP7_75t_SL g420 ( .A(n_421), .B(n_549), .C(n_584), .Y(n_420) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_451), .B(n_501), .C(n_539), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_433), .Y(n_423) );
AND2x2_ASAP7_75t_L g532 ( .A(n_424), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_424), .B(n_538), .Y(n_572) );
AND2x2_ASAP7_75t_L g597 ( .A(n_424), .B(n_552), .Y(n_597) );
INVx4_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g504 ( .A(n_425), .Y(n_504) );
OR2x2_ASAP7_75t_L g535 ( .A(n_425), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g543 ( .A(n_425), .B(n_443), .Y(n_543) );
AND2x2_ASAP7_75t_L g551 ( .A(n_425), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g578 ( .A(n_425), .B(n_579), .Y(n_578) );
NOR2x1_ASAP7_75t_L g589 ( .A(n_425), .B(n_581), .Y(n_589) );
AND2x4_ASAP7_75t_L g606 ( .A(n_425), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g644 ( .A(n_425), .Y(n_644) );
AND2x4_ASAP7_75t_SL g649 ( .A(n_425), .B(n_434), .Y(n_649) );
OR2x6_ASAP7_75t_L g425 ( .A(n_426), .B(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_433), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_433), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_443), .Y(n_433) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_434), .Y(n_544) );
INVx2_ASAP7_75t_L g580 ( .A(n_434), .Y(n_580) );
INVx1_ASAP7_75t_L g607 ( .A(n_434), .Y(n_607) );
AND2x2_ASAP7_75t_L g706 ( .A(n_434), .B(n_616), .Y(n_706) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_435), .Y(n_538) );
AND2x2_ASAP7_75t_L g552 ( .A(n_435), .B(n_443), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
INVx2_ASAP7_75t_L g581 ( .A(n_443), .Y(n_581) );
INVx2_ASAP7_75t_L g616 ( .A(n_443), .Y(n_616) );
OR2x2_ASAP7_75t_L g701 ( .A(n_443), .B(n_533), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_449), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_468), .B(n_488), .C(n_495), .Y(n_451) );
INVx2_ASAP7_75t_SL g590 ( .A(n_452), .Y(n_590) );
AND2x2_ASAP7_75t_L g596 ( .A(n_452), .B(n_469), .Y(n_596) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g492 ( .A(n_453), .Y(n_492) );
INVx1_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
INVx2_ASAP7_75t_L g523 ( .A(n_453), .Y(n_523) );
AND2x2_ASAP7_75t_L g547 ( .A(n_453), .B(n_471), .Y(n_547) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_453), .Y(n_576) );
OR2x2_ASAP7_75t_L g656 ( .A(n_453), .B(n_479), .Y(n_656) );
AND2x2_ASAP7_75t_L g522 ( .A(n_460), .B(n_523), .Y(n_522) );
NOR2x1_ASAP7_75t_SL g554 ( .A(n_460), .B(n_479), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g568 ( .A(n_469), .B(n_491), .Y(n_568) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
OR2x2_ASAP7_75t_L g500 ( .A(n_470), .B(n_479), .Y(n_500) );
BUFx2_ASAP7_75t_L g524 ( .A(n_470), .Y(n_524) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_470), .B(n_576), .Y(n_575) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
AND2x2_ASAP7_75t_L g553 ( .A(n_471), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g563 ( .A(n_471), .Y(n_563) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_471), .B(n_479), .Y(n_601) );
OR2x2_ASAP7_75t_L g676 ( .A(n_471), .B(n_493), .Y(n_676) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_SL g489 ( .A(n_479), .Y(n_489) );
AND2x2_ASAP7_75t_L g548 ( .A(n_479), .B(n_493), .Y(n_548) );
AND2x2_ASAP7_75t_L g619 ( .A(n_479), .B(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g640 ( .A(n_479), .Y(n_640) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_487), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g562 ( .A(n_491), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
BUFx2_ASAP7_75t_L g557 ( .A(n_492), .Y(n_557) );
AND2x2_ASAP7_75t_L g529 ( .A(n_493), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g620 ( .A(n_493), .Y(n_620) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
OR2x2_ASAP7_75t_L g566 ( .A(n_497), .B(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_SL g608 ( .A(n_497), .B(n_609), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g645 ( .A1(n_497), .A2(n_524), .A3(n_646), .B1(n_648), .B2(n_651), .C1(n_653), .C2(n_655), .Y(n_645) );
AND2x2_ASAP7_75t_L g710 ( .A(n_497), .B(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_498), .B(n_524), .Y(n_534) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_499), .A2(n_586), .A3(n_590), .B1(n_591), .B2(n_594), .C1(n_596), .C2(n_597), .Y(n_585) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g637 ( .A(n_500), .B(n_590), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_500), .A2(n_697), .B1(n_699), .B2(n_702), .Y(n_696) );
OR2x2_ASAP7_75t_L g714 ( .A(n_500), .B(n_663), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_524), .B(n_525), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
AOI221xp5_ASAP7_75t_SL g564 ( .A1(n_503), .A2(n_540), .B1(n_565), .B2(n_568), .C(n_569), .Y(n_564) );
AND2x2_ASAP7_75t_L g591 ( .A(n_503), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_504), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g633 ( .A(n_504), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g662 ( .A(n_505), .Y(n_662) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_522), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_506), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g604 ( .A(n_506), .Y(n_604) );
OR2x2_ASAP7_75t_L g611 ( .A(n_506), .B(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g654 ( .A(n_507), .B(n_616), .Y(n_654) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
AND2x4_ASAP7_75t_L g533 ( .A(n_508), .B(n_509), .Y(n_533) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
NOR2x1p5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_522), .B(n_583), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_522), .B(n_563), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_522), .Y(n_663) );
INVx1_ASAP7_75t_L g530 ( .A(n_523), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_531), .B1(n_534), .B2(n_535), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_SL g641 ( .A(n_529), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_530), .B(n_554), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_532), .B(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_SL g570 ( .A(n_532), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_532), .B(n_691), .Y(n_690) );
BUFx3_ASAP7_75t_L g558 ( .A(n_533), .Y(n_558) );
INVx2_ASAP7_75t_L g588 ( .A(n_533), .Y(n_588) );
AND2x2_ASAP7_75t_L g631 ( .A(n_533), .B(n_615), .Y(n_631) );
INVx1_ASAP7_75t_L g545 ( .A(n_535), .Y(n_545) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI21xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_545), .B(n_546), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g624 ( .A(n_543), .Y(n_624) );
INVx2_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g609 ( .A(n_548), .B(n_563), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_548), .A2(n_646), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_564), .Y(n_549) );
AOI32xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .A3(n_555), .B1(n_559), .B2(n_562), .Y(n_550) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_551), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_551), .A2(n_640), .B1(n_658), .B2(n_660), .C(n_666), .Y(n_657) );
AND2x2_ASAP7_75t_L g677 ( .A(n_551), .B(n_558), .Y(n_677) );
BUFx2_ASAP7_75t_L g561 ( .A(n_552), .Y(n_561) );
INVx1_ASAP7_75t_L g686 ( .A(n_552), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_552), .Y(n_691) );
INVx1_ASAP7_75t_SL g684 ( .A(n_553), .Y(n_684) );
INVx2_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
AND2x2_ASAP7_75t_L g679 ( .A(n_555), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g651 ( .A(n_557), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g623 ( .A(n_558), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_558), .B(n_649), .Y(n_671) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g583 ( .A(n_563), .Y(n_583) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g573 ( .A(n_567), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g582 ( .A(n_567), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g687 ( .A(n_568), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B1(n_577), .B2(n_582), .Y(n_569) );
INVx2_ASAP7_75t_SL g661 ( .A(n_571), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_571), .B(n_700), .Y(n_702) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_573), .A2(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g646 ( .A(n_578), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g593 ( .A(n_579), .Y(n_593) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g635 ( .A(n_581), .Y(n_635) );
INVx1_ASAP7_75t_L g680 ( .A(n_582), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_598), .C(n_621), .Y(n_584) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
AND2x2_ASAP7_75t_L g665 ( .A(n_587), .B(n_606), .Y(n_665) );
OR2x2_ASAP7_75t_L g704 ( .A(n_587), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_588), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g600 ( .A(n_590), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g667 ( .A(n_593), .B(n_604), .Y(n_667) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_596), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B1(n_606), .B2(n_608), .C(n_610), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_599), .A2(n_622), .B(n_625), .Y(n_621) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g652 ( .A(n_601), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_601), .B(n_695), .Y(n_694) );
INVxp33_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g613 ( .A(n_609), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B1(n_614), .B2(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g716 ( .A(n_612), .Y(n_716) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g695 ( .A(n_620), .Y(n_695) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_672), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_645), .C(n_657), .D(n_669), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_632), .B(n_636), .C(n_638), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g668 ( .A(n_631), .Y(n_668) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_633), .A2(n_639), .B(n_642), .Y(n_638) );
INVx2_ASAP7_75t_L g717 ( .A(n_634), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_635), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g650 ( .A(n_635), .Y(n_650) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OR2x2_ASAP7_75t_L g712 ( .A(n_640), .B(n_676), .Y(n_712) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_647), .Y(n_683) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g653 ( .A(n_649), .B(n_654), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_649), .A2(n_679), .B(n_681), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_649), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g707 ( .A(n_649), .Y(n_707) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .C(n_688), .D(n_709), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_685), .B2(n_687), .Y(n_681) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI211xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_692), .B(n_696), .C(n_703), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_707), .B(n_708), .Y(n_703) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_713), .B(n_715), .Y(n_709) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx3_ASAP7_75t_SL g722 ( .A(n_718), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_719), .Y(n_718) );
CKINVDCx6p67_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_736), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_732), .B(n_735), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_SL g749 ( .A(n_733), .B(n_735), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_733), .A2(n_752), .B(n_755), .Y(n_751) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx3_ASAP7_75t_L g742 ( .A(n_737), .Y(n_742) );
BUFx2_ASAP7_75t_L g745 ( .A(n_737), .Y(n_745) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_742), .B(n_743), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx2_ASAP7_75t_L g755 ( .A(n_745), .Y(n_755) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx11_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx8_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
endmodule