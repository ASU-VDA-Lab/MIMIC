module fake_ariane_2282_n_26 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_26);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_26;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_17;
wire n_18;
wire n_11;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

AND3x2_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_7),
.C(n_0),
.Y(n_10)
);

NAND3xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_2),
.C(n_6),
.Y(n_11)
);

NAND2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_4),
.Y(n_12)
);

OAI22xp33_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_3),
.B1(n_6),
.B2(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

O2A1O1Ixp5_ASAP7_75t_SL g15 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.C(n_8),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_9),
.B(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_12),
.Y(n_17)
);

BUFx2_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_13),
.B(n_11),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_16),
.C(n_20),
.Y(n_24)
);

AO22x2_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_22),
.B1(n_18),
.B2(n_8),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_22),
.B(n_21),
.Y(n_26)
);


endmodule