module fake_jpeg_28819_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_12),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_6),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_7),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_17),
.B1(n_33),
.B2(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_57),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_5),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_38),
.B1(n_45),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_67),
.B1(n_16),
.B2(n_22),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_49),
.C(n_38),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_81),
.Y(n_88)
);

OAI211xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_20),
.B(n_30),
.C(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_8),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_9),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_94),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_36),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_25),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_15),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_91),
.C(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_26),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_84),
.B(n_89),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_104),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_88),
.B(n_97),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_85),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_86),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_109),
.Y(n_110)
);


endmodule