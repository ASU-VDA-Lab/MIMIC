module fake_jpeg_12181_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_19),
.B(n_1),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_17),
.B(n_4),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_15),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_36),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_32),
.B1(n_39),
.B2(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_15),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

FAx1_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_27),
.CI(n_23),
.CON(n_50),
.SN(n_50)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_53),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_14),
.B(n_24),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_21),
.B1(n_18),
.B2(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_29),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_29),
.A2(n_17),
.B1(n_23),
.B2(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_3),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_4),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_36),
.B1(n_30),
.B2(n_11),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_55),
.B1(n_52),
.B2(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_7),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_12),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_59),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_44),
.B(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_67),
.B1(n_66),
.B2(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_100),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_62),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_83),
.B1(n_72),
.B2(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_92),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_80),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_99),
.C(n_87),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_104),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_101),
.C(n_95),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.C(n_109),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_97),
.C(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_120),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_105),
.B1(n_81),
.B2(n_108),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_106),
.Y(n_121)
);

NAND4xp25_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.C(n_123),
.D(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_105),
.A3(n_64),
.B1(n_71),
.B2(n_70),
.C1(n_85),
.C2(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_76),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_51),
.A3(n_46),
.B1(n_73),
.B2(n_68),
.C1(n_125),
.C2(n_54),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_54),
.C(n_48),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B(n_46),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_30),
.Y(n_132)
);


endmodule