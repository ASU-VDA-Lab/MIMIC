module fake_jpeg_10341_n_132 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_SL g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx4f_ASAP7_75t_SL g12 ( 
.A(n_1),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_29),
.B1(n_10),
.B2(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp67_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_4),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_15),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_4),
.CON(n_29),
.SN(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_10),
.B1(n_18),
.B2(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_41),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_10),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_28),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_15),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_58),
.B1(n_51),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_49),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_25),
.C(n_17),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_30),
.B(n_35),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_26),
.B1(n_57),
.B2(n_16),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_5),
.B(n_6),
.Y(n_73)
);

NOR4xp25_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_79),
.B1(n_72),
.B2(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_82),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_62),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_23),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_85),
.C(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_81),
.C(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_99),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_88),
.B1(n_69),
.B2(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_100),
.B(n_86),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_62),
.C(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_115),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_62),
.C(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_96),
.B1(n_95),
.B2(n_69),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_101),
.B(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_107),
.B(n_105),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_119),
.B(n_20),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_120),
.Y(n_124)
);

AOI31xp67_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_104),
.A3(n_61),
.B(n_17),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_112),
.C(n_39),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_128),
.Y(n_130)
);

NOR2xp67_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_9),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_25),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_127),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_130),
.Y(n_132)
);


endmodule