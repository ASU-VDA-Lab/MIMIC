module fake_jpeg_24630_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_0),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_8),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_48),
.B1(n_33),
.B2(n_18),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_25),
.B1(n_31),
.B2(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_34),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_57),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_18),
.B1(n_17),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_22),
.B1(n_17),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_90),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_73),
.B1(n_84),
.B2(n_92),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_88),
.B1(n_62),
.B2(n_75),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_82),
.B(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_27),
.B1(n_33),
.B2(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_14),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_37),
.B1(n_35),
.B2(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_19),
.B1(n_20),
.B2(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_37),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_66),
.B1(n_60),
.B2(n_61),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_87),
.B1(n_82),
.B2(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_108),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_45),
.B1(n_44),
.B2(n_63),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_117),
.B1(n_89),
.B2(n_92),
.Y(n_148)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_109),
.B1(n_112),
.B2(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_44),
.B1(n_64),
.B2(n_53),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_116),
.Y(n_125)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_91),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_76),
.A2(n_85),
.B1(n_94),
.B2(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_80),
.Y(n_149)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_134),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_120),
.C(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_124),
.C(n_133),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_81),
.C(n_70),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_70),
.B(n_72),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_142),
.B(n_145),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_72),
.C(n_92),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_82),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_98),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_147),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_73),
.B1(n_71),
.B2(n_80),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_117),
.B1(n_104),
.B2(n_19),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_110),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_92),
.C(n_42),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_97),
.C(n_95),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_53),
.B(n_92),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_92),
.B1(n_35),
.B2(n_82),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_149),
.B(n_35),
.Y(n_180)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_117),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_112),
.CI(n_97),
.CON(n_151),
.SN(n_151)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_172),
.B1(n_127),
.B2(n_119),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_169),
.C(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_115),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_107),
.B1(n_98),
.B2(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_99),
.C(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_101),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_80),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_58),
.B(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_134),
.B1(n_132),
.B2(n_122),
.C(n_127),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_133),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_182),
.C(n_185),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_142),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_180),
.B(n_177),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_124),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_129),
.C(n_144),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_196),
.C(n_199),
.Y(n_216)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_136),
.B1(n_139),
.B2(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_192),
.B1(n_198),
.B2(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_136),
.B1(n_146),
.B2(n_137),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_178),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_153),
.C(n_160),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_148),
.B1(n_141),
.B2(n_128),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_128),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_151),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_166),
.B1(n_163),
.B2(n_170),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_171),
.C(n_164),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_168),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_213),
.C(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_188),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_59),
.B1(n_65),
.B2(n_24),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_175),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_220),
.B(n_221),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_224),
.B1(n_187),
.B2(n_58),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_167),
.B1(n_151),
.B2(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_20),
.B1(n_65),
.B2(n_58),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_222),
.B1(n_226),
.B2(n_58),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_162),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_176),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_225),
.C(n_184),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_156),
.B1(n_174),
.B2(n_161),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_138),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_35),
.CI(n_58),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_185),
.C(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_194),
.C(n_200),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_203),
.B1(n_205),
.B2(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_192),
.C(n_190),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_235),
.C(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_193),
.C(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_237),
.B1(n_221),
.B2(n_219),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_214),
.C(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_65),
.B1(n_59),
.B2(n_51),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_208),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_224),
.B1(n_226),
.B2(n_211),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_59),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_9),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_255),
.C(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_8),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_232),
.C(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_3),
.C(n_4),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_234),
.B1(n_238),
.B2(n_10),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_265),
.B1(n_7),
.B2(n_11),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_16),
.B(n_8),
.Y(n_260)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_263),
.A3(n_13),
.B1(n_15),
.B2(n_5),
.C(n_6),
.Y(n_274)
);

NAND4xp25_ASAP7_75t_SL g262 ( 
.A(n_256),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_4),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_246),
.B(n_250),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_254),
.B(n_6),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_15),
.B1(n_7),
.B2(n_10),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_3),
.C(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_251),
.C(n_5),
.Y(n_269)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_270),
.C(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_7),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_262),
.B(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_13),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_5),
.C(n_258),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_278),
.B(n_282),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_271),
.CI(n_272),
.CON(n_288),
.SN(n_288)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_283),
.B(n_280),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_269),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_285),
.B(n_281),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_288),
.C(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_291),
.Y(n_292)
);


endmodule