module fake_jpeg_28380_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12f_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_51),
.Y(n_88)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_27),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx2_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_33),
.B1(n_16),
.B2(n_23),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_20),
.B1(n_28),
.B2(n_33),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_87),
.Y(n_115)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_29),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_62),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_88),
.B(n_1),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_66),
.B1(n_45),
.B2(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_110),
.B1(n_114),
.B2(n_30),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_77),
.B1(n_70),
.B2(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_116),
.B1(n_33),
.B2(n_16),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_17),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_113),
.C(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_32),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_117),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_66),
.B1(n_61),
.B2(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_84),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_51),
.C(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_20),
.B1(n_16),
.B2(n_33),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_126),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_79),
.B1(n_71),
.B2(n_88),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_125),
.B(n_129),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_114),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

XNOR2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_31),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_134),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_107),
.Y(n_149)
);

CKINVDCx6p67_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_32),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_71),
.B1(n_27),
.B2(n_31),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_16),
.B1(n_18),
.B2(n_30),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_18),
.B1(n_30),
.B2(n_32),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_31),
.C(n_25),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_123),
.C(n_134),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_97),
.A3(n_112),
.B1(n_96),
.B2(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_112),
.B(n_117),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_145),
.B(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_163),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_164),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_95),
.B(n_111),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_166),
.B(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_126),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_105),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_172),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_175),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_92),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_142),
.B1(n_129),
.B2(n_118),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_181),
.B1(n_158),
.B2(n_170),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_182),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_134),
.B1(n_99),
.B2(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_193),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_151),
.B(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_141),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_158),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_168),
.B(n_163),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_140),
.B(n_101),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_144),
.B1(n_143),
.B2(n_94),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_202),
.B1(n_157),
.B2(n_156),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_110),
.B1(n_106),
.B2(n_103),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_165),
.C(n_171),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_204),
.C(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_167),
.C(n_175),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_146),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_211),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_177),
.B1(n_181),
.B2(n_184),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_223),
.B(n_224),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_187),
.C(n_176),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_157),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_103),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_31),
.C(n_21),
.Y(n_246)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_2),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_176),
.B1(n_182),
.B2(n_178),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_218),
.B1(n_21),
.B2(n_31),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_185),
.B(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_238),
.B1(n_241),
.B2(n_245),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_197),
.B1(n_193),
.B2(n_200),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_187),
.B(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_183),
.B1(n_179),
.B2(n_116),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_179),
.B(n_11),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_15),
.B(n_3),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_18),
.B1(n_2),
.B2(n_0),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_204),
.C(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_213),
.C(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_256),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_205),
.Y(n_253)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_225),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_21),
.C(n_25),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_25),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_230),
.B1(n_245),
.B2(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_236),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_10),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_238),
.B1(n_240),
.B2(n_242),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_253),
.B1(n_237),
.B2(n_2),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_250),
.C(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_271),
.A2(n_243),
.B1(n_235),
.B2(n_254),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_285),
.B1(n_267),
.B2(n_266),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_9),
.B(n_4),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_284),
.B(n_7),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_10),
.C(n_5),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_273),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_263),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_7),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_280),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_298),
.B(n_295),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_278),
.B(n_275),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_302),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_287),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_301),
.B(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_299),
.B1(n_283),
.B2(n_12),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_8),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_2),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_8),
.B(n_13),
.Y(n_308)
);


endmodule