module real_aes_1639_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_964, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_965, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_964;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_965;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_865;
wire n_666;
wire n_551;
wire n_884;
wire n_537;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_744;
wire n_384;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_552;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_727;
wire n_397;
wire n_749;
wire n_385;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_0), .A2(n_340), .B1(n_418), .B2(n_688), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_1), .A2(n_260), .B1(n_457), .B2(n_737), .Y(n_736) );
AOI222xp33_ASAP7_75t_L g915 ( .A1(n_2), .A2(n_916), .B1(n_934), .B2(n_938), .C1(n_940), .C2(n_960), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_2), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_3), .A2(n_302), .B1(n_412), .B2(n_685), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_4), .A2(n_61), .B1(n_509), .B2(n_510), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_5), .A2(n_343), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_6), .A2(n_171), .B1(n_457), .B2(n_460), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_7), .A2(n_261), .B1(n_390), .B2(n_695), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_8), .A2(n_40), .B1(n_440), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_9), .A2(n_320), .B1(n_464), .B2(n_645), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_10), .A2(n_28), .B1(n_409), .B2(n_624), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_11), .A2(n_296), .B1(n_362), .B2(n_379), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_12), .A2(n_92), .B1(n_729), .B2(n_730), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_13), .A2(n_77), .B1(n_385), .B2(n_386), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_14), .A2(n_188), .B1(n_362), .B2(n_379), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_15), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_16), .A2(n_347), .B1(n_679), .B2(n_710), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_17), .A2(n_151), .B1(n_435), .B2(n_438), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g808 ( .A1(n_18), .A2(n_248), .B1(n_392), .B2(n_697), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_19), .A2(n_203), .B1(n_450), .B2(n_454), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_20), .A2(n_50), .B1(n_665), .B2(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_21), .A2(n_183), .B1(n_498), .B2(n_499), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_22), .A2(n_125), .B1(n_688), .B2(n_712), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_23), .A2(n_338), .B1(n_492), .B2(n_493), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_24), .A2(n_127), .B1(n_528), .B2(n_529), .Y(n_527) );
AO22x2_ASAP7_75t_L g476 ( .A1(n_25), .A2(n_477), .B1(n_500), .B2(n_501), .Y(n_476) );
INVx1_ASAP7_75t_L g500 ( .A(n_25), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_26), .A2(n_185), .B1(n_645), .B2(n_780), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_27), .A2(n_227), .B1(n_450), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_29), .A2(n_172), .B1(n_566), .B2(n_568), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_30), .A2(n_238), .B1(n_390), .B2(n_392), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_31), .B(n_489), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_32), .A2(n_176), .B1(n_443), .B2(n_446), .Y(n_442) );
AO222x2_ASAP7_75t_L g922 ( .A1(n_33), .A2(n_133), .B1(n_233), .B2(n_679), .C1(n_682), .C2(n_710), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_34), .A2(n_126), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_35), .A2(n_314), .B1(n_685), .B2(n_686), .Y(n_925) );
INVx1_ASAP7_75t_L g654 ( .A(n_36), .Y(n_654) );
INVx1_ASAP7_75t_SL g377 ( .A(n_37), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_37), .B(n_47), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_38), .A2(n_225), .B1(n_670), .B2(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_39), .A2(n_54), .B1(n_528), .B2(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_41), .A2(n_307), .B1(n_513), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_42), .A2(n_192), .B1(n_418), .B2(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_43), .A2(n_87), .B1(n_412), .B2(n_685), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_44), .B(n_558), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_45), .A2(n_219), .B1(n_617), .B2(n_695), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_46), .B(n_682), .Y(n_847) );
AO22x2_ASAP7_75t_L g372 ( .A1(n_47), .A2(n_326), .B1(n_366), .B2(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_48), .A2(n_199), .B1(n_563), .B2(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_49), .B(n_682), .Y(n_681) );
XOR2xp5_ASAP7_75t_L g764 ( .A(n_51), .B(n_765), .Y(n_764) );
XOR2xp5_ASAP7_75t_L g813 ( .A(n_51), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_52), .A2(n_91), .B1(n_450), .B2(n_452), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_53), .B(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_55), .A2(n_121), .B1(n_577), .B2(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g378 ( .A(n_56), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_57), .A2(n_90), .B1(n_435), .B2(n_438), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_58), .A2(n_103), .B1(n_379), .B2(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_59), .A2(n_204), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g828 ( .A1(n_60), .A2(n_310), .B1(n_485), .B2(n_755), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_62), .A2(n_184), .B1(n_568), .B2(n_877), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_63), .A2(n_136), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_64), .A2(n_335), .B1(n_524), .B2(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_65), .A2(n_274), .B1(n_499), .B2(n_672), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_66), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_67), .A2(n_231), .B1(n_385), .B2(n_386), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_68), .A2(n_168), .B1(n_685), .B2(n_686), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_69), .A2(n_169), .B1(n_443), .B2(n_524), .Y(n_607) );
AO22x2_ASAP7_75t_L g369 ( .A1(n_70), .A2(n_180), .B1(n_366), .B2(n_370), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_71), .A2(n_344), .B1(n_401), .B2(n_405), .Y(n_400) );
AO22x1_ASAP7_75t_L g516 ( .A1(n_72), .A2(n_270), .B1(n_517), .B2(n_520), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_73), .A2(n_322), .B1(n_394), .B2(n_666), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_74), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g953 ( .A1(n_75), .A2(n_135), .B1(n_386), .B2(n_619), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_76), .A2(n_152), .B1(n_576), .B2(n_577), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_78), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_79), .A2(n_148), .B1(n_785), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_80), .A2(n_220), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_81), .A2(n_312), .B1(n_679), .B2(n_680), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_82), .A2(n_213), .B1(n_487), .B2(n_556), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g928 ( .A1(n_83), .A2(n_119), .B1(n_386), .B2(n_929), .Y(n_928) );
AOI222xp33_ASAP7_75t_L g861 ( .A1(n_84), .A2(n_96), .B1(n_187), .B2(n_418), .C1(n_419), .C2(n_682), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_85), .A2(n_268), .B1(n_362), .B2(n_379), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_86), .A2(n_191), .B1(n_362), .B2(n_695), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_88), .A2(n_348), .B1(n_418), .B2(n_419), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_89), .A2(n_333), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_93), .A2(n_228), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_94), .A2(n_166), .B1(n_436), .B2(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_95), .A2(n_140), .B1(n_604), .B2(n_619), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_97), .A2(n_118), .B1(n_385), .B2(n_386), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_98), .A2(n_254), .B1(n_510), .B2(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_99), .A2(n_202), .B1(n_379), .B2(n_697), .Y(n_855) );
OA22x2_ASAP7_75t_L g856 ( .A1(n_100), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_100), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_101), .A2(n_107), .B1(n_695), .B2(n_697), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_102), .A2(n_277), .B1(n_362), .B2(n_695), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_104), .A2(n_131), .B1(n_493), .B2(n_528), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_105), .A2(n_211), .B1(n_577), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_106), .A2(n_328), .B1(n_385), .B2(n_386), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_108), .A2(n_290), .B1(n_496), .B2(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_109), .A2(n_223), .B1(n_362), .B2(n_379), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_110), .A2(n_190), .B1(n_409), .B2(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_111), .A2(n_247), .B1(n_429), .B2(n_514), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_112), .A2(n_246), .B1(n_833), .B2(n_834), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_113), .A2(n_145), .B1(n_430), .B2(n_881), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_114), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_115), .A2(n_329), .B1(n_362), .B2(n_397), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_116), .A2(n_206), .B1(n_679), .B2(n_680), .Y(n_678) );
AO22x2_ASAP7_75t_L g365 ( .A1(n_117), .A2(n_273), .B1(n_366), .B2(n_367), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_120), .A2(n_224), .B1(n_464), .B2(n_526), .Y(n_525) );
XOR2x2_ASAP7_75t_L g358 ( .A(n_122), .B(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_123), .A2(n_311), .B1(n_570), .B2(n_573), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_124), .A2(n_141), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_128), .A2(n_161), .B1(n_390), .B2(n_392), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_129), .A2(n_300), .B1(n_379), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_130), .A2(n_201), .B1(n_484), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_132), .A2(n_332), .B1(n_536), .B2(n_537), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_134), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_137), .A2(n_146), .B1(n_695), .B2(n_697), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_138), .A2(n_263), .B1(n_528), .B2(n_642), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_139), .A2(n_163), .B1(n_409), .B2(n_412), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_142), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_143), .A2(n_170), .B1(n_412), .B2(n_685), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_144), .A2(n_285), .B1(n_392), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_147), .A2(n_317), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_149), .A2(n_165), .B1(n_218), .B2(n_466), .C1(n_467), .C2(n_468), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_150), .A2(n_303), .B1(n_468), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_153), .A2(n_318), .B1(n_385), .B2(n_386), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_154), .A2(n_257), .B1(n_679), .B2(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_155), .B(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_156), .A2(n_198), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_157), .A2(n_295), .B1(n_679), .B2(n_680), .Y(n_804) );
AO22x2_ASAP7_75t_L g700 ( .A1(n_158), .A2(n_701), .B1(n_714), .B2(n_715), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_158), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_159), .B(n_533), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_160), .A2(n_234), .B1(n_394), .B2(n_397), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_162), .A2(n_181), .B1(n_566), .B2(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_164), .B(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_167), .A2(n_284), .B1(n_679), .B2(n_680), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_173), .A2(n_264), .B1(n_419), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_174), .A2(n_301), .B1(n_401), .B2(n_487), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_175), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_177), .A2(n_214), .B1(n_556), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_178), .A2(n_194), .B1(n_480), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_179), .A2(n_226), .B1(n_688), .B2(n_712), .Y(n_805) );
INVx1_ASAP7_75t_L g903 ( .A(n_180), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_182), .A2(n_280), .B1(n_430), .B2(n_596), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_186), .A2(n_281), .B1(n_390), .B2(n_392), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_189), .A2(n_349), .B1(n_362), .B2(n_379), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_193), .A2(n_242), .B1(n_379), .B2(n_528), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_195), .A2(n_241), .B1(n_412), .B2(n_685), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_196), .A2(n_298), .B1(n_642), .B2(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_197), .B(n_682), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_200), .A2(n_269), .B1(n_553), .B2(n_555), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_205), .A2(n_209), .B1(n_551), .B2(n_591), .Y(n_590) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_207), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_208), .B(n_558), .Y(n_557) );
XNOR2x1_ASAP7_75t_L g725 ( .A(n_210), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g913 ( .A(n_212), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_215), .A2(n_286), .B1(n_429), .B2(n_481), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_216), .A2(n_342), .B1(n_390), .B2(n_392), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_217), .A2(n_279), .B1(n_537), .B2(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g914 ( .A(n_221), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_222), .A2(n_426), .B1(n_469), .B2(n_470), .Y(n_425) );
INVx1_ASAP7_75t_L g470 ( .A(n_222), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_229), .A2(n_331), .B1(n_624), .B2(n_662), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_230), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_232), .B(n_422), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_235), .A2(n_276), .B1(n_741), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g585 ( .A(n_236), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_237), .A2(n_294), .B1(n_555), .B2(n_593), .Y(n_745) );
XNOR2x1_ASAP7_75t_L g844 ( .A(n_239), .B(n_845), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_240), .A2(n_291), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_243), .A2(n_272), .B1(n_385), .B2(n_386), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_244), .A2(n_278), .B1(n_640), .B2(n_784), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_245), .A2(n_292), .B1(n_480), .B2(n_744), .Y(n_772) );
XOR2x2_ASAP7_75t_L g544 ( .A(n_249), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_250), .A2(n_346), .B1(n_487), .B2(n_556), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_251), .A2(n_309), .B1(n_409), .B2(n_513), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_252), .A2(n_339), .B1(n_576), .B2(n_779), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_253), .A2(n_258), .B1(n_602), .B2(n_604), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g748 ( .A(n_255), .B(n_749), .Y(n_748) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_255), .B(n_749), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g924 ( .A1(n_256), .A2(n_271), .B1(n_688), .B2(n_712), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_259), .A2(n_262), .B1(n_362), .B2(n_379), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_265), .A2(n_297), .B1(n_392), .B2(n_617), .Y(n_692) );
OA22x2_ASAP7_75t_L g610 ( .A1(n_266), .A2(n_611), .B1(n_612), .B2(n_627), .Y(n_610) );
INVx1_ASAP7_75t_L g627 ( .A(n_266), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_267), .B(n_533), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_273), .B(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_275), .A2(n_324), .B1(n_498), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_282), .A2(n_306), .B1(n_392), .B2(n_572), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_283), .A2(n_315), .B1(n_468), .B2(n_554), .Y(n_826) );
INVx3_ASAP7_75t_L g366 ( .A(n_287), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_288), .A2(n_305), .B1(n_732), .B2(n_733), .Y(n_731) );
XOR2x1_ASAP7_75t_L g631 ( .A(n_289), .B(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_293), .A2(n_316), .B1(n_570), .B2(n_606), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_299), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_304), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_308), .B(n_489), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_313), .Y(n_789) );
OAI22xp5_ASAP7_75t_SL g940 ( .A1(n_319), .A2(n_941), .B1(n_958), .B2(n_959), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_319), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_321), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_323), .A2(n_330), .B1(n_685), .B2(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g698 ( .A(n_325), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_327), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g898 ( .A(n_334), .Y(n_898) );
NAND2xp5_ASAP7_75t_SL g912 ( .A(n_334), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g899 ( .A(n_336), .Y(n_899) );
AND2x2_ASAP7_75t_R g962 ( .A(n_336), .B(n_898), .Y(n_962) );
INVx1_ASAP7_75t_L g515 ( .A(n_337), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_337), .A2(n_507), .B1(n_539), .B2(n_964), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_337), .A2(n_522), .B1(n_531), .B2(n_965), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_337), .B(n_516), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_341), .B(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_345), .B(n_422), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_894), .B(n_905), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_580), .Y(n_351) );
AOI21xp33_ASAP7_75t_SL g894 ( .A1(n_352), .A2(n_580), .B(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_544), .B1(n_578), .B2(n_579), .Y(n_352) );
INVx1_ASAP7_75t_L g579 ( .A(n_353), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_472), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
AO22x2_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B1(n_425), .B2(n_471), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
XNOR2x1_ASAP7_75t_L g503 ( .A(n_358), .B(n_504), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_399), .C(n_416), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_384), .C(n_389), .D(n_393), .Y(n_360) );
AND2x6_ASAP7_75t_L g362 ( .A(n_363), .B(n_371), .Y(n_362) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g396 ( .A(n_363), .B(n_380), .Y(n_396) );
AND2x2_ASAP7_75t_L g424 ( .A(n_363), .B(n_415), .Y(n_424) );
AND2x2_ASAP7_75t_L g445 ( .A(n_363), .B(n_371), .Y(n_445) );
AND2x4_ASAP7_75t_L g459 ( .A(n_363), .B(n_391), .Y(n_459) );
AND2x2_ASAP7_75t_L g617 ( .A(n_363), .B(n_391), .Y(n_617) );
AND2x4_ASAP7_75t_L g682 ( .A(n_363), .B(n_415), .Y(n_682) );
AND2x2_ASAP7_75t_L g697 ( .A(n_363), .B(n_380), .Y(n_697) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g383 ( .A(n_365), .Y(n_383) );
AND2x2_ASAP7_75t_L g388 ( .A(n_365), .B(n_369), .Y(n_388) );
AND2x4_ASAP7_75t_L g398 ( .A(n_365), .B(n_368), .Y(n_398) );
INVx2_ASAP7_75t_L g367 ( .A(n_366), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_366), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_366), .Y(n_373) );
OAI22x1_ASAP7_75t_L g375 ( .A1(n_366), .A2(n_376), .B1(n_377), .B2(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_366), .Y(n_376) );
INVxp67_ASAP7_75t_L g420 ( .A(n_368), .Y(n_420) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g382 ( .A(n_369), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g385 ( .A(n_371), .B(n_382), .Y(n_385) );
AND2x2_ASAP7_75t_L g418 ( .A(n_371), .B(n_398), .Y(n_418) );
AND2x4_ASAP7_75t_L g437 ( .A(n_371), .B(n_398), .Y(n_437) );
AND2x2_ASAP7_75t_L g451 ( .A(n_371), .B(n_382), .Y(n_451) );
AND2x2_ASAP7_75t_L g712 ( .A(n_371), .B(n_398), .Y(n_712) );
AND2x2_ASAP7_75t_SL g929 ( .A(n_371), .B(n_382), .Y(n_929) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx2_ASAP7_75t_L g381 ( .A(n_372), .Y(n_381) );
BUFx2_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
AND2x2_ASAP7_75t_L g415 ( .A(n_372), .B(n_375), .Y(n_415) );
AND2x4_ASAP7_75t_L g380 ( .A(n_374), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g391 ( .A(n_375), .B(n_381), .Y(n_391) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
AND2x6_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
AND2x4_ASAP7_75t_L g392 ( .A(n_380), .B(n_388), .Y(n_392) );
AND2x4_ASAP7_75t_L g397 ( .A(n_380), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g448 ( .A(n_380), .B(n_382), .Y(n_448) );
AND2x4_ASAP7_75t_L g464 ( .A(n_380), .B(n_388), .Y(n_464) );
AND2x2_ASAP7_75t_L g695 ( .A(n_380), .B(n_398), .Y(n_695) );
AND2x2_ASAP7_75t_L g411 ( .A(n_382), .B(n_391), .Y(n_411) );
AND2x4_ASAP7_75t_L g685 ( .A(n_382), .B(n_391), .Y(n_685) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AND2x4_ASAP7_75t_L g454 ( .A(n_387), .B(n_388), .Y(n_454) );
AND2x2_ASAP7_75t_L g403 ( .A(n_388), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_388), .B(n_404), .Y(n_680) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_388), .B(n_404), .Y(n_710) );
AND2x2_ASAP7_75t_L g407 ( .A(n_391), .B(n_398), .Y(n_407) );
AND2x4_ASAP7_75t_L g679 ( .A(n_391), .B(n_398), .Y(n_679) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_SL g462 ( .A(n_395), .Y(n_462) );
INVx2_ASAP7_75t_L g492 ( .A(n_395), .Y(n_492) );
INVx3_ASAP7_75t_SL g528 ( .A(n_395), .Y(n_528) );
INVx4_ASAP7_75t_L g572 ( .A(n_395), .Y(n_572) );
INVx2_ASAP7_75t_SL g672 ( .A(n_395), .Y(n_672) );
INVx8_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g460 ( .A(n_397), .Y(n_460) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_397), .Y(n_493) );
INVx2_ASAP7_75t_L g530 ( .A(n_397), .Y(n_530) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_397), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g556 ( .A(n_402), .Y(n_556) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx12f_ASAP7_75t_L g468 ( .A(n_403), .Y(n_468) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g769 ( .A(n_406), .Y(n_769) );
INVx2_ASAP7_75t_L g884 ( .A(n_406), .Y(n_884) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx5_ASAP7_75t_L g467 ( .A(n_407), .Y(n_467) );
BUFx3_ASAP7_75t_L g487 ( .A(n_407), .Y(n_487) );
BUFx3_ASAP7_75t_L g554 ( .A(n_407), .Y(n_554) );
INVx2_ASAP7_75t_SL g597 ( .A(n_409), .Y(n_597) );
INVx4_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g549 ( .A(n_410), .Y(n_549) );
INVx2_ASAP7_75t_L g662 ( .A(n_410), .Y(n_662) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_411), .Y(n_429) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
AND2x4_ASAP7_75t_L g433 ( .A(n_413), .B(n_415), .Y(n_433) );
AND2x2_ASAP7_75t_L g686 ( .A(n_413), .B(n_415), .Y(n_686) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g419 ( .A(n_415), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g440 ( .A(n_415), .B(n_420), .Y(n_440) );
AND2x2_ASAP7_75t_L g688 ( .A(n_415), .B(n_420), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_421), .Y(n_416) );
INVx4_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
INVx3_ASAP7_75t_L g489 ( .A(n_423), .Y(n_489) );
BUFx2_ASAP7_75t_L g534 ( .A(n_423), .Y(n_534) );
INVx3_ASAP7_75t_SL g560 ( .A(n_423), .Y(n_560) );
INVx4_ASAP7_75t_SL g752 ( .A(n_423), .Y(n_752) );
INVx6_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g471 ( .A(n_425), .Y(n_471) );
INVx1_ASAP7_75t_L g469 ( .A(n_426), .Y(n_469) );
NAND4xp75_ASAP7_75t_L g426 ( .A(n_427), .B(n_441), .C(n_455), .D(n_465), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_434), .Y(n_427) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
BUFx3_ASAP7_75t_L g514 ( .A(n_433), .Y(n_514) );
BUFx6f_ASAP7_75t_SL g624 ( .A(n_433), .Y(n_624) );
BUFx4f_ASAP7_75t_L g744 ( .A(n_433), .Y(n_744) );
BUFx4f_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g536 ( .A(n_436), .Y(n_536) );
BUFx2_ASAP7_75t_L g551 ( .A(n_436), .Y(n_551) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
BUFx2_ASAP7_75t_L g755 ( .A(n_437), .Y(n_755) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
INVx2_ASAP7_75t_L g537 ( .A(n_439), .Y(n_537) );
INVx2_ASAP7_75t_L g591 ( .A(n_439), .Y(n_591) );
INVx1_ASAP7_75t_L g659 ( .A(n_439), .Y(n_659) );
INVx2_ASAP7_75t_SL g741 ( .A(n_439), .Y(n_741) );
INVx6_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .Y(n_441) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g665 ( .A(n_444), .Y(n_665) );
INVx2_ASAP7_75t_SL g732 ( .A(n_444), .Y(n_732) );
INVx3_ASAP7_75t_L g761 ( .A(n_444), .Y(n_761) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
BUFx2_ASAP7_75t_L g785 ( .A(n_445), .Y(n_785) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g524 ( .A(n_447), .Y(n_524) );
INVx2_ASAP7_75t_SL g640 ( .A(n_447), .Y(n_640) );
INVx2_ASAP7_75t_L g666 ( .A(n_447), .Y(n_666) );
INVx2_ASAP7_75t_SL g733 ( .A(n_447), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_447), .A2(n_782), .B1(n_783), .B2(n_786), .Y(n_781) );
INVx2_ASAP7_75t_L g836 ( .A(n_447), .Y(n_836) );
INVx8_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g519 ( .A(n_451), .Y(n_519) );
BUFx3_ASAP7_75t_L g619 ( .A(n_451), .Y(n_619) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g568 ( .A(n_453), .Y(n_568) );
INVx3_ASAP7_75t_L g670 ( .A(n_453), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_453), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
INVx2_ASAP7_75t_L g834 ( .A(n_453), .Y(n_834) );
INVx5_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g520 ( .A(n_454), .Y(n_520) );
BUFx2_ASAP7_75t_L g604 ( .A(n_454), .Y(n_604) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_461), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
INVx1_ASAP7_75t_SL g576 ( .A(n_458), .Y(n_576) );
INVx2_ASAP7_75t_L g600 ( .A(n_458), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_458), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_775) );
INVx6_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx3_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
BUFx3_ASAP7_75t_L g645 ( .A(n_459), .Y(n_645) );
BUFx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g499 ( .A(n_464), .Y(n_499) );
BUFx2_ASAP7_75t_SL g577 ( .A(n_464), .Y(n_577) );
INVx2_ASAP7_75t_L g738 ( .A(n_464), .Y(n_738) );
BUFx3_ASAP7_75t_L g780 ( .A(n_464), .Y(n_780) );
BUFx3_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
INVx2_ASAP7_75t_L g886 ( .A(n_468), .Y(n_886) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_502), .B(n_542), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_475), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g501 ( .A(n_477), .Y(n_501) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .C(n_486), .D(n_488), .Y(n_478) );
BUFx6f_ASAP7_75t_SL g881 ( .A(n_480), .Y(n_881) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g889 ( .A(n_484), .Y(n_889) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_487), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .C(n_495), .D(n_497), .Y(n_490) );
INVx1_ASAP7_75t_L g794 ( .A(n_492), .Y(n_794) );
INVx2_ASAP7_75t_L g574 ( .A(n_493), .Y(n_574) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
INVx2_ASAP7_75t_L g564 ( .A(n_496), .Y(n_564) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g543 ( .A(n_503), .Y(n_543) );
NAND4xp75_ASAP7_75t_L g504 ( .A(n_505), .B(n_538), .C(n_540), .D(n_541), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_521), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .C(n_516), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g539 ( .A(n_512), .Y(n_539) );
BUFx6f_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g603 ( .A(n_518), .Y(n_603) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_518), .Y(n_735) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g567 ( .A(n_519), .Y(n_567) );
INVx1_ASAP7_75t_L g833 ( .A(n_519), .Y(n_833) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_522), .B(n_531), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .C(n_527), .Y(n_522) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g642 ( .A(n_530), .Y(n_642) );
INVx1_ASAP7_75t_L g730 ( .A(n_530), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .Y(n_531) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g578 ( .A(n_544), .Y(n_578) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_546), .B(n_561), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_552), .D(n_557), .Y(n_546) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g594 ( .A(n_554), .Y(n_594) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI21xp33_ASAP7_75t_SL g824 ( .A1(n_559), .A2(n_825), .B(n_826), .Y(n_824) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_560), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .C(n_569), .D(n_575), .Y(n_561) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_572), .Y(n_729) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_574), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
XNOR2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_721), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_647), .B1(n_717), .B2(n_718), .Y(n_581) );
INVx1_ASAP7_75t_L g717 ( .A(n_582), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_630), .B1(n_631), .B2(n_646), .Y(n_582) );
INVx1_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_608), .B1(n_628), .B2(n_629), .Y(n_583) );
INVx2_ASAP7_75t_L g628 ( .A(n_584), .Y(n_628) );
XNOR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_598), .Y(n_586) );
NAND4xp25_ASAP7_75t_SL g587 ( .A(n_588), .B(n_590), .C(n_592), .D(n_595), .Y(n_587) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .C(n_605), .D(n_607), .Y(n_598) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_603), .Y(n_790) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g629 ( .A(n_610), .Y(n_629) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g612 ( .A(n_613), .B(n_621), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .C(n_620), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
BUFx2_ASAP7_75t_L g877 ( .A(n_619), .Y(n_877) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .C(n_625), .D(n_626), .Y(n_621) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_638), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .C(n_636), .D(n_637), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .C(n_643), .D(n_644), .Y(n_638) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OA22x2_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_699), .B2(n_716), .Y(n_649) );
OA22x2_ASAP7_75t_L g720 ( .A1(n_650), .A2(n_651), .B1(n_699), .B2(n_716), .Y(n_720) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OA22x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_673), .B2(n_674), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
XNOR2x2_ASAP7_75t_SL g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .C(n_660), .D(n_661), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .C(n_669), .D(n_671), .Y(n_663) );
INVx3_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
XOR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_698), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_689), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_683), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_678), .B(n_681), .Y(n_677) );
INVx2_ASAP7_75t_SL g945 ( .A(n_682), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVxp67_ASAP7_75t_L g716 ( .A(n_699), .Y(n_716) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g715 ( .A(n_701), .Y(n_715) );
NOR2xp67_ASAP7_75t_L g701 ( .A(n_702), .B(n_707), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .C(n_705), .D(n_706), .Y(n_702) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_708), .B(n_709), .C(n_711), .D(n_713), .Y(n_707) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
XNOR2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_817), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_763), .B1(n_815), .B2(n_816), .Y(n_722) );
INVx2_ASAP7_75t_L g815 ( .A(n_723), .Y(n_815) );
OA22x2_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_746), .B2(n_747), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_739), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_731), .C(n_734), .D(n_736), .Y(n_727) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .C(n_743), .D(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_748), .A2(n_799), .B1(n_800), .B2(n_812), .Y(n_798) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_757), .Y(n_749) );
NAND4xp25_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .C(n_754), .D(n_756), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .C(n_760), .D(n_762), .Y(n_757) );
INVx3_ASAP7_75t_SL g816 ( .A(n_763), .Y(n_816) );
OA22x2_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_796), .B1(n_797), .B2(n_813), .Y(n_763) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_774), .C(n_787), .Y(n_765) );
AND3x1_ASAP7_75t_L g814 ( .A(n_766), .B(n_774), .C(n_787), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_771), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_770), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_781), .Y(n_774) );
INVxp67_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
BUFx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_807), .Y(n_801) );
NAND4xp25_ASAP7_75t_SL g802 ( .A(n_803), .B(n_804), .C(n_805), .D(n_806), .Y(n_802) );
NAND4xp25_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .C(n_810), .D(n_811), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_841), .B1(n_892), .B2(n_893), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_819), .Y(n_892) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
XNOR2x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_840), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_830), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_837), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVxp33_ASAP7_75t_L g893 ( .A(n_841), .Y(n_893) );
AO22x2_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_871), .B2(n_891), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AO22x2_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_856), .B1(n_869), .B2(n_870), .Y(n_843) );
INVx1_ASAP7_75t_L g869 ( .A(n_844), .Y(n_869) );
OR2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_851), .Y(n_845) );
NAND4xp25_ASAP7_75t_SL g846 ( .A(n_847), .B(n_848), .C(n_849), .D(n_850), .Y(n_846) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .C(n_854), .D(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g870 ( .A(n_856), .Y(n_870) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2x1_ASAP7_75t_L g859 ( .A(n_860), .B(n_864), .Y(n_859) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .C(n_863), .Y(n_860) );
NAND4xp25_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .C(n_867), .D(n_868), .Y(n_864) );
INVx1_ASAP7_75t_L g891 ( .A(n_871), .Y(n_891) );
XOR2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_890), .Y(n_871) );
NOR2x1_ASAP7_75t_L g872 ( .A(n_873), .B(n_879), .Y(n_872) );
NAND4xp25_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .C(n_876), .D(n_878), .Y(n_873) );
NAND4xp25_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .C(n_883), .D(n_887), .Y(n_879) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_897), .B(n_901), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
INVx1_ASAP7_75t_L g910 ( .A(n_899), .Y(n_910) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_914), .B(n_915), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
AND2x2_ASAP7_75t_SL g908 ( .A(n_909), .B(n_911), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
OR2x2_ASAP7_75t_L g939 ( .A(n_910), .B(n_911), .Y(n_939) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
XNOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
AND2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_926), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_931), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_930), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_935), .Y(n_934) );
CKINVDCx20_ASAP7_75t_R g935 ( .A(n_936), .Y(n_935) );
CKINVDCx6p67_ASAP7_75t_R g936 ( .A(n_937), .Y(n_936) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_939), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_941), .Y(n_959) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
NAND2x1_ASAP7_75t_L g942 ( .A(n_943), .B(n_951), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_944), .B(n_948), .Y(n_943) );
OAI21xp5_ASAP7_75t_SL g944 ( .A1(n_945), .A2(n_946), .B(n_947), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_949), .B(n_950), .Y(n_948) );
NOR2x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_955), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
INVx1_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
endmodule