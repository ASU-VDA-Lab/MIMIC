module real_jpeg_7390_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_1),
.B(n_185),
.C(n_188),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_1),
.A2(n_34),
.B1(n_172),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_1),
.B(n_124),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_46),
.B1(n_227),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_54),
.B1(n_57),
.B2(n_62),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_43),
.B1(n_62),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_3),
.Y(n_146)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_5),
.A2(n_76),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_76),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_47),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_11),
.A2(n_48),
.B1(n_97),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_12),
.A2(n_103),
.B1(n_126),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_126),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_176),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_175),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_18),
.B(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_74),
.C(n_106),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_19),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_45),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_20),
.B(n_45),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.A3(n_29),
.B1(n_33),
.B2(n_38),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_22),
.A2(n_131),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_23),
.Y(n_129)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_26),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_33),
.A2(n_34),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_34),
.B(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_34),
.B(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_40),
.A2(n_102),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B(n_63),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_46),
.B(n_68),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_46),
.A2(n_202),
.B(n_204),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_46),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_46),
.A2(n_65),
.B1(n_212),
.B2(n_227),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_47),
.Y(n_145)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_52),
.Y(n_153)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_52),
.Y(n_239)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_60),
.Y(n_229)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_66),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_74),
.B(n_106),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_83),
.B1(n_95),
.B2(n_96),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_75),
.A2(n_83),
.B1(n_95),
.B2(n_192),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_83),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_83),
.A2(n_95),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_86),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_124),
.B2(n_125),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_110),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_162),
.B2(n_163),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_155),
.B2(n_161),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_150),
.B(n_154),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_173),
.B2(n_174),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B(n_168),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_243),
.B(n_247),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_208),
.B(n_242),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_195),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_179),
.B(n_195),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_223),
.B(n_241),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_222),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_233),
.B(n_240),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);


endmodule