module fake_netlist_1_5884_n_22 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_0), .B(n_1), .Y(n_11) );
NAND3xp33_ASAP7_75t_L g12 ( .A(n_2), .B(n_4), .C(n_0), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_8), .B(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_1), .Y(n_15) );
AO31x2_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_2), .A3(n_3), .B(n_7), .Y(n_16) );
NOR2x1_ASAP7_75t_L g17 ( .A(n_15), .B(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AOI221xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_13), .B1(n_16), .B2(n_3), .C(n_10), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_19), .B(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NAND2x1p5_ASAP7_75t_L g22 ( .A(n_21), .B(n_9), .Y(n_22) );
endmodule