module real_aes_12232_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_0), .A2(n_461), .B1(n_464), .B2(n_473), .C(n_476), .Y(n_460) );
AOI21xp33_ASAP7_75t_L g531 ( .A1(n_0), .A2(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g897 ( .A(n_1), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_1), .A2(n_70), .B1(n_924), .B2(n_925), .C(n_926), .Y(n_923) );
INVx1_ASAP7_75t_L g835 ( .A(n_2), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_2), .A2(n_30), .B1(n_740), .B2(n_865), .C(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_3), .A2(n_245), .B1(n_299), .B2(n_526), .Y(n_904) );
INVx1_ASAP7_75t_L g936 ( .A(n_3), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_4), .A2(n_72), .B1(n_643), .B2(n_644), .Y(n_651) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_4), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_5), .A2(n_299), .B(n_972), .Y(n_1084) );
INVx1_ASAP7_75t_L g1102 ( .A(n_5), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_6), .A2(n_60), .B1(n_1110), .B2(n_1132), .Y(n_1131) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_7), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_8), .Y(n_261) );
AND2x2_ASAP7_75t_L g351 ( .A(n_8), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g406 ( .A(n_8), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_8), .B(n_184), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g955 ( .A1(n_9), .A2(n_146), .B1(n_287), .B2(n_607), .C(n_902), .Y(n_955) );
INVx1_ASAP7_75t_L g991 ( .A(n_9), .Y(n_991) );
INVx1_ASAP7_75t_L g388 ( .A(n_10), .Y(n_388) );
INVxp67_ASAP7_75t_L g729 ( .A(n_11), .Y(n_729) );
OAI222xp33_ASAP7_75t_L g744 ( .A1(n_11), .A2(n_45), .B1(n_234), .B2(n_313), .C1(n_586), .C2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g397 ( .A(n_12), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_13), .A2(n_22), .B1(n_482), .B2(n_485), .C(n_486), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_13), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_14), .A2(n_78), .B1(n_784), .B2(n_786), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_14), .A2(n_31), .B1(n_350), .B2(n_411), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_15), .A2(n_210), .B1(n_821), .B2(n_839), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_15), .A2(n_64), .B1(n_519), .B2(n_598), .C(n_874), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g901 ( .A1(n_16), .A2(n_37), .B1(n_519), .B2(n_749), .C(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g938 ( .A(n_16), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_17), .A2(n_64), .B1(n_841), .B2(n_843), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_17), .A2(n_210), .B1(n_756), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_18), .A2(n_69), .B1(n_1132), .B2(n_1146), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_19), .Y(n_1342) );
AOI221xp5_ASAP7_75t_L g1399 ( .A1(n_20), .A2(n_206), .B1(n_874), .B2(n_971), .C(n_972), .Y(n_1399) );
INVx1_ASAP7_75t_L g1420 ( .A(n_20), .Y(n_1420) );
OAI221xp5_ASAP7_75t_L g1064 ( .A1(n_21), .A2(n_512), .B1(n_1065), .B2(n_1070), .C(n_1075), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_21), .A2(n_166), .B1(n_813), .B2(n_1098), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_22), .Y(n_541) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_23), .A2(n_141), .B1(n_402), .B2(n_812), .C(n_813), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_23), .A2(n_205), .B1(n_451), .B2(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g282 ( .A(n_24), .Y(n_282) );
OR2x2_ASAP7_75t_L g441 ( .A(n_24), .B(n_330), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_25), .A2(n_174), .B1(n_577), .B2(n_578), .C(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g590 ( .A(n_25), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_26), .A2(n_118), .B1(n_1122), .B2(n_1128), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_27), .A2(n_59), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g806 ( .A(n_27), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_28), .A2(n_218), .B1(n_865), .B2(n_1029), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1039 ( .A1(n_28), .A2(n_218), .B1(n_925), .B2(n_926), .C(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g730 ( .A(n_29), .Y(n_730) );
INVx1_ASAP7_75t_L g834 ( .A(n_30), .Y(n_834) );
OAI222xp33_ASAP7_75t_L g822 ( .A1(n_31), .A2(n_141), .B1(n_148), .B2(n_657), .C1(n_823), .C2(n_825), .Y(n_822) );
BUFx2_ASAP7_75t_L g284 ( .A(n_32), .Y(n_284) );
BUFx2_ASAP7_75t_L g318 ( .A(n_32), .Y(n_318) );
INVx1_ASAP7_75t_L g332 ( .A(n_32), .Y(n_332) );
OR2x2_ASAP7_75t_L g484 ( .A(n_32), .B(n_413), .Y(n_484) );
INVx1_ASAP7_75t_L g1169 ( .A(n_33), .Y(n_1169) );
INVx1_ASAP7_75t_L g1006 ( .A(n_34), .Y(n_1006) );
INVx1_ASAP7_75t_L g556 ( .A(n_35), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_36), .A2(n_153), .B1(n_414), .B2(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g522 ( .A(n_36), .Y(n_522) );
INVx1_ASAP7_75t_L g931 ( .A(n_37), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_38), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_39), .A2(n_65), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1422 ( .A1(n_39), .A2(n_65), .B1(n_486), .B2(n_924), .C(n_925), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_40), .A2(n_131), .B1(n_663), .B2(n_673), .Y(n_1083) );
INVx1_ASAP7_75t_L g1103 ( .A(n_40), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_41), .A2(n_171), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_41), .A2(n_223), .B1(n_311), .B2(n_682), .C(n_685), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_42), .A2(n_82), .B1(n_432), .B2(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_42), .A2(n_82), .B1(n_503), .B2(n_507), .Y(n_502) );
INVx1_ASAP7_75t_L g713 ( .A(n_43), .Y(n_713) );
INVx1_ASAP7_75t_L g1206 ( .A(n_44), .Y(n_1206) );
INVxp67_ASAP7_75t_L g727 ( .A(n_45), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_46), .A2(n_186), .B1(n_784), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1045 ( .A(n_46), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_47), .A2(n_54), .B1(n_849), .B2(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g878 ( .A(n_47), .Y(n_878) );
INVx1_ASAP7_75t_L g566 ( .A(n_48), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_49), .Y(n_333) );
INVx1_ASAP7_75t_L g794 ( .A(n_50), .Y(n_794) );
OAI221xp5_ASAP7_75t_L g815 ( .A1(n_50), .A2(n_79), .B1(n_816), .B2(n_818), .C(n_819), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_51), .A2(n_94), .B1(n_1122), .B2(n_1128), .Y(n_1149) );
INVx1_ASAP7_75t_L g467 ( .A(n_52), .Y(n_467) );
AOI21xp33_ASAP7_75t_L g518 ( .A1(n_52), .A2(n_519), .B(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_53), .A2(n_87), .B1(n_647), .B2(n_648), .Y(n_650) );
INVxp33_ASAP7_75t_SL g694 ( .A(n_53), .Y(n_694) );
INVx1_ASAP7_75t_L g872 ( .A(n_54), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_55), .A2(n_166), .B1(n_507), .B2(n_510), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_55), .A2(n_240), .B1(n_1092), .B2(n_1096), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_56), .A2(n_66), .B1(n_519), .B2(n_750), .C(n_874), .Y(n_1019) );
INVxp67_ASAP7_75t_SL g1048 ( .A(n_56), .Y(n_1048) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_57), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_58), .A2(n_182), .B1(n_311), .B2(n_312), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_58), .A2(n_244), .B1(n_347), .B2(n_357), .Y(n_346) );
INVx1_ASAP7_75t_L g804 ( .A(n_59), .Y(n_804) );
INVx1_ASAP7_75t_L g1338 ( .A(n_61), .Y(n_1338) );
AOI221xp5_ASAP7_75t_L g1372 ( .A1(n_61), .A2(n_119), .B1(n_1373), .B2(n_1374), .C(n_1375), .Y(n_1372) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_62), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_63), .A2(n_104), .B1(n_1122), .B2(n_1128), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_66), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_67), .A2(n_236), .B1(n_526), .B2(n_876), .Y(n_1409) );
INVx1_ASAP7_75t_L g1425 ( .A(n_67), .Y(n_1425) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_68), .A2(n_123), .B1(n_390), .B2(n_562), .C(n_563), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_68), .A2(n_83), .B1(n_601), .B2(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g898 ( .A(n_70), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_71), .Y(n_470) );
INVxp33_ASAP7_75t_L g692 ( .A(n_72), .Y(n_692) );
INVx1_ASAP7_75t_L g565 ( .A(n_73), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_73), .A2(n_123), .B1(n_595), .B2(n_596), .C(n_598), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_74), .A2(n_137), .B1(n_761), .B2(n_763), .C(n_764), .Y(n_760) );
OAI221xp5_ASAP7_75t_L g766 ( .A1(n_74), .A2(n_154), .B1(n_767), .B2(n_768), .C(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g1349 ( .A(n_75), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_75), .A2(n_248), .B1(n_292), .B2(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g281 ( .A(n_76), .Y(n_281) );
INVx1_ASAP7_75t_L g330 ( .A(n_76), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_77), .A2(n_227), .B1(n_609), .B2(n_784), .Y(n_956) );
INVx1_ASAP7_75t_L g999 ( .A(n_77), .Y(n_999) );
INVx1_ASAP7_75t_L g814 ( .A(n_78), .Y(n_814) );
INVx1_ASAP7_75t_L g793 ( .A(n_79), .Y(n_793) );
INVx1_ASAP7_75t_L g1015 ( .A(n_80), .Y(n_1015) );
INVx1_ASAP7_75t_L g581 ( .A(n_81), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_81), .A2(n_174), .B1(n_586), .B2(n_588), .C(n_589), .Y(n_585) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_83), .Y(n_564) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_84), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_84), .A2(n_198), .B1(n_665), .B2(n_667), .Y(n_664) );
NAND2xp33_ASAP7_75t_SL g895 ( .A(n_85), .B(n_786), .Y(n_895) );
INVx1_ASAP7_75t_L g919 ( .A(n_85), .Y(n_919) );
INVx1_ASAP7_75t_L g1071 ( .A(n_86), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_86), .A2(n_149), .B1(n_813), .B2(n_1090), .Y(n_1089) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_87), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_88), .A2(n_142), .B1(n_497), .B2(n_500), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_88), .A2(n_192), .B1(n_288), .B2(n_526), .Y(n_530) );
INVx1_ASAP7_75t_L g573 ( .A(n_89), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_89), .A2(n_133), .B1(n_534), .B2(n_606), .C(n_607), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_90), .A2(n_106), .B1(n_1122), .B2(n_1128), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_91), .A2(n_192), .B1(n_490), .B2(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g528 ( .A(n_91), .Y(n_528) );
XNOR2xp5_ASAP7_75t_L g703 ( .A(n_92), .B(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_92), .A2(n_189), .B1(n_1122), .B2(n_1128), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1150 ( .A1(n_93), .A2(n_121), .B1(n_1132), .B2(n_1146), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_94), .A2(n_1061), .B1(n_1105), .B2(n_1106), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_94), .Y(n_1105) );
INVxp67_ASAP7_75t_L g711 ( .A(n_95), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_95), .A2(n_156), .B1(n_519), .B2(n_749), .C(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_96), .Y(n_889) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_97), .A2(n_548), .B(n_583), .Y(n_547) );
INVx1_ASAP7_75t_L g617 ( .A(n_97), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_98), .A2(n_155), .B1(n_684), .B2(n_763), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g802 ( .A1(n_98), .A2(n_414), .B(n_474), .Y(n_802) );
INVx1_ASAP7_75t_L g1137 ( .A(n_99), .Y(n_1137) );
INVx1_ASAP7_75t_L g582 ( .A(n_100), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_101), .A2(n_216), .B1(n_1026), .B2(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1038 ( .A(n_101), .Y(n_1038) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_102), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_103), .A2(n_193), .B1(n_299), .B2(n_874), .C(n_972), .Y(n_1024) );
INVx1_ASAP7_75t_L g1037 ( .A(n_103), .Y(n_1037) );
INVx1_ASAP7_75t_L g253 ( .A(n_105), .Y(n_253) );
AO22x1_ASAP7_75t_SL g1134 ( .A1(n_107), .A2(n_195), .B1(n_1122), .B2(n_1128), .Y(n_1134) );
INVx1_ASAP7_75t_L g912 ( .A(n_108), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g1412 ( .A(n_109), .Y(n_1412) );
INVx1_ASAP7_75t_L g1204 ( .A(n_110), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_111), .A2(n_175), .B1(n_845), .B2(n_847), .Y(n_844) );
INVx1_ASAP7_75t_L g879 ( .A(n_111), .Y(n_879) );
AO221x2_ASAP7_75t_L g1163 ( .A1(n_112), .A2(n_235), .B1(n_1110), .B2(n_1164), .C(n_1165), .Y(n_1163) );
OAI221xp5_ASAP7_75t_SL g569 ( .A1(n_113), .A2(n_214), .B1(n_570), .B2(n_571), .C(n_572), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_113), .A2(n_214), .B1(n_287), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_114), .A2(n_177), .B1(n_756), .B2(n_966), .Y(n_1400) );
INVx1_ASAP7_75t_L g1417 ( .A(n_114), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_115), .Y(n_1367) );
CKINVDCx5p33_ASAP7_75t_R g1359 ( .A(n_116), .Y(n_1359) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_117), .A2(n_199), .B1(n_292), .B2(n_789), .Y(n_894) );
INVx1_ASAP7_75t_L g922 ( .A(n_117), .Y(n_922) );
XOR2xp5_ASAP7_75t_L g457 ( .A(n_118), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g1343 ( .A(n_119), .Y(n_1343) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_120), .Y(n_1362) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_122), .A2(n_157), .B1(n_239), .B2(n_500), .C1(n_707), .C2(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g738 ( .A(n_122), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_124), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_125), .Y(n_854) );
INVx1_ASAP7_75t_L g882 ( .A(n_126), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_127), .B(n_773), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_128), .A2(n_246), .B1(n_607), .B2(n_971), .C(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g979 ( .A(n_128), .Y(n_979) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_129), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g1079 ( .A(n_130), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_131), .A2(n_229), .B1(n_493), .B2(n_497), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_132), .A2(n_225), .B1(n_286), .B2(n_291), .Y(n_285) );
INVx1_ASAP7_75t_L g370 ( .A(n_132), .Y(n_370) );
INVx1_ASAP7_75t_L g575 ( .A(n_133), .Y(n_575) );
INVx1_ASAP7_75t_L g961 ( .A(n_134), .Y(n_961) );
OAI221xp5_ASAP7_75t_L g983 ( .A1(n_134), .A2(n_211), .B1(n_485), .B2(n_984), .C(n_986), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g1411 ( .A(n_135), .Y(n_1411) );
INVx1_ASAP7_75t_L g853 ( .A(n_136), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_136), .A2(n_207), .B1(n_288), .B2(n_314), .Y(n_867) );
OAI332xp33_ASAP7_75t_L g709 ( .A1(n_137), .A2(n_473), .A3(n_710), .B1(n_715), .B2(n_721), .B3(n_728), .C1(n_733), .C2(n_734), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_138), .A2(n_230), .B1(n_1132), .B2(n_1146), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_139), .A2(n_1393), .B1(n_1432), .B2(n_1433), .Y(n_1392) );
CKINVDCx5p33_ASAP7_75t_R g1432 ( .A(n_139), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_140), .Y(n_1406) );
INVx1_ASAP7_75t_L g536 ( .A(n_142), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_143), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_144), .Y(n_658) );
INVx1_ASAP7_75t_L g1018 ( .A(n_145), .Y(n_1018) );
INVx1_ASAP7_75t_L g995 ( .A(n_146), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_147), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_148), .A2(n_205), .B1(n_562), .B2(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1067 ( .A(n_149), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_150), .A2(n_159), .B1(n_292), .B2(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g797 ( .A(n_150), .Y(n_797) );
XOR2x2_ASAP7_75t_L g618 ( .A(n_151), .B(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_152), .A2(n_244), .B1(n_298), .B2(n_304), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_152), .A2(n_182), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g517 ( .A(n_153), .Y(n_517) );
INVx1_ASAP7_75t_L g759 ( .A(n_154), .Y(n_759) );
INVx1_ASAP7_75t_L g801 ( .A(n_155), .Y(n_801) );
INVx1_ASAP7_75t_L g716 ( .A(n_156), .Y(n_716) );
INVx1_ASAP7_75t_L g754 ( .A(n_157), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g1074 ( .A1(n_158), .A2(n_287), .B(n_520), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_158), .A2(n_228), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
INVx1_ASAP7_75t_L g798 ( .A(n_159), .Y(n_798) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_160), .Y(n_255) );
AND3x2_ASAP7_75t_L g1114 ( .A(n_160), .B(n_253), .C(n_1115), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_160), .B(n_253), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_161), .A2(n_220), .B1(n_1110), .B2(n_1132), .Y(n_1174) );
CKINVDCx5p33_ASAP7_75t_R g1340 ( .A(n_162), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1407 ( .A1(n_163), .A2(n_208), .B1(n_750), .B2(n_1384), .C(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1428 ( .A(n_163), .Y(n_1428) );
INVx2_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
INVx1_ASAP7_75t_L g1030 ( .A(n_165), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_167), .Y(n_634) );
INVx1_ASAP7_75t_L g552 ( .A(n_168), .Y(n_552) );
INVxp33_ASAP7_75t_SL g636 ( .A(n_169), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_169), .A2(n_209), .B1(n_670), .B2(n_672), .C(n_674), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_170), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_171), .A2(n_190), .B1(n_609), .B2(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g1115 ( .A(n_172), .Y(n_1115) );
INVx1_ASAP7_75t_L g1139 ( .A(n_173), .Y(n_1139) );
INVx1_ASAP7_75t_L g863 ( .A(n_175), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_176), .A2(n_238), .B1(n_414), .B2(n_472), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_176), .A2(n_238), .B1(n_510), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g1421 ( .A(n_177), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_178), .A2(n_221), .B1(n_298), .B2(n_304), .Y(n_297) );
INVx1_ASAP7_75t_L g382 ( .A(n_178), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_179), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g1398 ( .A(n_180), .Y(n_1398) );
INVx1_ASAP7_75t_L g1352 ( .A(n_181), .Y(n_1352) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_181), .A2(n_241), .B1(n_520), .B2(n_1373), .C(n_1384), .Y(n_1383) );
CKINVDCx20_ASAP7_75t_R g1166 ( .A(n_183), .Y(n_1166) );
INVx1_ASAP7_75t_L g268 ( .A(n_184), .Y(n_268) );
INVx2_ASAP7_75t_L g352 ( .A(n_184), .Y(n_352) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_185), .B(n_656), .Y(n_1062) );
INVx1_ASAP7_75t_L g1051 ( .A(n_186), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_187), .A2(n_1010), .B1(n_1058), .B2(n_1059), .Y(n_1009) );
INVx1_ASAP7_75t_L g1059 ( .A(n_187), .Y(n_1059) );
INVx1_ASAP7_75t_L g856 ( .A(n_188), .Y(n_856) );
AOI21xp33_ASAP7_75t_L g868 ( .A1(n_188), .A2(n_534), .B(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_190), .A2(n_223), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_191), .A2(n_194), .B1(n_1109), .B2(n_1202), .C(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1035 ( .A(n_193), .Y(n_1035) );
AOI222xp33_ASAP7_75t_L g1331 ( .A1(n_194), .A2(n_1332), .B1(n_1390), .B2(n_1392), .C1(n_1434), .C2(n_1436), .Y(n_1331) );
XNOR2x1_ASAP7_75t_L g1333 ( .A(n_194), .B(n_1334), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g958 ( .A(n_196), .Y(n_958) );
INVx1_ASAP7_75t_L g417 ( .A(n_197), .Y(n_417) );
INVxp67_ASAP7_75t_SL g626 ( .A(n_198), .Y(n_626) );
INVx1_ASAP7_75t_L g917 ( .A(n_199), .Y(n_917) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_200), .B(n_274), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_201), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_202), .Y(n_959) );
INVx1_ASAP7_75t_L g631 ( .A(n_203), .Y(n_631) );
INVx1_ASAP7_75t_L g393 ( .A(n_204), .Y(n_393) );
INVx1_ASAP7_75t_L g1418 ( .A(n_206), .Y(n_1418) );
INVx1_ASAP7_75t_L g857 ( .A(n_207), .Y(n_857) );
INVx1_ASAP7_75t_L g1426 ( .A(n_208), .Y(n_1426) );
INVxp33_ASAP7_75t_SL g628 ( .A(n_209), .Y(n_628) );
INVx1_ASAP7_75t_L g962 ( .A(n_211), .Y(n_962) );
INVx1_ASAP7_75t_L g741 ( .A(n_212), .Y(n_741) );
INVx1_ASAP7_75t_L g975 ( .A(n_213), .Y(n_975) );
INVx1_ASAP7_75t_L g1023 ( .A(n_215), .Y(n_1023) );
INVx1_ASAP7_75t_L g1034 ( .A(n_216), .Y(n_1034) );
INVx1_ASAP7_75t_L g718 ( .A(n_217), .Y(n_718) );
INVx1_ASAP7_75t_L g1113 ( .A(n_219), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_219), .B(n_1125), .Y(n_1130) );
INVx1_ASAP7_75t_L g378 ( .A(n_221), .Y(n_378) );
INVx2_ASAP7_75t_L g265 ( .A(n_222), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g969 ( .A(n_224), .Y(n_969) );
INVx1_ASAP7_75t_L g364 ( .A(n_225), .Y(n_364) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_226), .A2(n_299), .B(n_534), .Y(n_896) );
INVx1_ASAP7_75t_L g921 ( .A(n_226), .Y(n_921) );
INVx1_ASAP7_75t_L g989 ( .A(n_227), .Y(n_989) );
INVx1_ASAP7_75t_L g1069 ( .A(n_228), .Y(n_1069) );
INVx1_ASAP7_75t_L g1081 ( .A(n_229), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1344 ( .A1(n_231), .A2(n_232), .B1(n_708), .B2(n_1040), .C(n_1345), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_231), .A2(n_232), .B1(n_667), .B2(n_1371), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_233), .Y(n_1360) );
INVxp67_ASAP7_75t_L g722 ( .A(n_234), .Y(n_722) );
INVx1_ASAP7_75t_L g1429 ( .A(n_236), .Y(n_1429) );
INVx1_ASAP7_75t_L g1413 ( .A(n_237), .Y(n_1413) );
INVx1_ASAP7_75t_L g742 ( .A(n_239), .Y(n_742) );
OAI211xp5_ASAP7_75t_SL g1076 ( .A1(n_240), .A2(n_503), .B(n_1077), .C(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g1354 ( .A(n_241), .Y(n_1354) );
BUFx3_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
INVx1_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
BUFx3_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
INVx1_ASAP7_75t_L g933 ( .A(n_245), .Y(n_933) );
INVx1_ASAP7_75t_L g981 ( .A(n_246), .Y(n_981) );
INVx1_ASAP7_75t_L g1014 ( .A(n_247), .Y(n_1014) );
INVx1_ASAP7_75t_L g1356 ( .A(n_248), .Y(n_1356) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_269), .B(n_1107), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
AND2x4_ASAP7_75t_L g1391 ( .A(n_251), .B(n_257), .Y(n_1391) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_SL g1435 ( .A(n_252), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_252), .B(n_254), .Y(n_1440) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_254), .B(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_268), .Y(n_385) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g474 ( .A(n_261), .B(n_475), .Y(n_474) );
OR2x6_ASAP7_75t_L g262 ( .A(n_263), .B(n_267), .Y(n_262) );
BUFx2_ASAP7_75t_L g381 ( .A(n_263), .Y(n_381) );
INVx1_ASAP7_75t_L g399 ( .A(n_263), .Y(n_399) );
OR2x2_ASAP7_75t_L g500 ( .A(n_263), .B(n_484), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_263), .A2(n_395), .B1(n_564), .B2(n_565), .Y(n_563) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_263), .A2(n_395), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx2_ASAP7_75t_SL g720 ( .A(n_263), .Y(n_720) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_263), .Y(n_1005) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_263), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x4_ASAP7_75t_L g355 ( .A(n_265), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g361 ( .A(n_265), .Y(n_361) );
INVx2_ASAP7_75t_L g369 ( .A(n_265), .Y(n_369) );
INVx1_ASAP7_75t_L g377 ( .A(n_265), .Y(n_377) );
AND2x2_ASAP7_75t_L g416 ( .A(n_265), .B(n_266), .Y(n_416) );
INVx2_ASAP7_75t_L g356 ( .A(n_266), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_266), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g376 ( .A(n_266), .Y(n_376) );
INVx1_ASAP7_75t_L g423 ( .A(n_266), .Y(n_423) );
INVx1_ASAP7_75t_L g434 ( .A(n_266), .Y(n_434) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_700), .Y(n_269) );
BUFx2_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AO22x2_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_618), .B1(n_698), .B2(n_699), .Y(n_271) );
INVx1_ASAP7_75t_L g698 ( .A(n_272), .Y(n_698) );
XNOR2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_456), .Y(n_272) );
NAND4xp75_ASAP7_75t_L g274 ( .A(n_275), .B(n_345), .C(n_437), .D(n_446), .Y(n_274) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_276), .B(n_321), .Y(n_275) );
AOI33xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_285), .A3(n_297), .B1(n_309), .B2(n_310), .B3(n_315), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_278), .Y(n_277) );
OR2x6_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
INVx1_ASAP7_75t_L g903 ( .A(n_279), .Y(n_903) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_SL g520 ( .A(n_280), .Y(n_520) );
BUFx3_ASAP7_75t_L g599 ( .A(n_280), .Y(n_599) );
INVx1_ASAP7_75t_L g778 ( .A(n_280), .Y(n_778) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x4_ASAP7_75t_L g319 ( .A(n_281), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
AND2x2_ASAP7_75t_L g480 ( .A(n_283), .B(n_403), .Y(n_480) );
AND2x4_ASAP7_75t_L g560 ( .A(n_283), .B(n_385), .Y(n_560) );
INVx2_ASAP7_75t_L g613 ( .A(n_283), .Y(n_613) );
AND2x4_ASAP7_75t_L g641 ( .A(n_283), .B(n_385), .Y(n_641) );
OR2x2_ASAP7_75t_L g777 ( .A(n_283), .B(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g911 ( .A(n_283), .Y(n_911) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g436 ( .A(n_284), .Y(n_436) );
OR2x6_ASAP7_75t_L g473 ( .A(n_284), .B(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
INVx1_ASAP7_75t_L g671 ( .A(n_287), .Y(n_671) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_SL g449 ( .A(n_288), .Y(n_449) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_288), .Y(n_505) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_288), .Y(n_519) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_288), .Y(n_663) );
BUFx3_ASAP7_75t_L g789 ( .A(n_288), .Y(n_789) );
BUFx2_ASAP7_75t_L g966 ( .A(n_288), .Y(n_966) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_288), .Y(n_1026) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g455 ( .A(n_289), .Y(n_455) );
INVx2_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_295), .Y(n_308) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x6_ASAP7_75t_L g443 ( .A(n_293), .B(n_440), .Y(n_443) );
OR2x2_ASAP7_75t_L g827 ( .A(n_293), .B(n_440), .Y(n_827) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
INVx2_ASAP7_75t_L g508 ( .A(n_294), .Y(n_508) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_294), .Y(n_673) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
INVx1_ASAP7_75t_L g454 ( .A(n_296), .Y(n_454) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g438 ( .A(n_299), .B(n_439), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_299), .A2(n_536), .B(n_537), .C(n_543), .Y(n_535) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g688 ( .A(n_300), .Y(n_688) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g445 ( .A(n_301), .B(n_328), .Y(n_445) );
INVx6_ASAP7_75t_L g533 ( .A(n_301), .Y(n_533) );
BUFx2_ASAP7_75t_L g876 ( .A(n_301), .Y(n_876) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g689 ( .A(n_306), .B(n_690), .Y(n_689) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_307), .Y(n_607) );
INVx2_ASAP7_75t_L g787 ( .A(n_307), .Y(n_787) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_308), .Y(n_514) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g588 ( .A(n_314), .Y(n_588) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_314), .Y(n_609) );
INVx1_ASAP7_75t_L g747 ( .A(n_314), .Y(n_747) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_314), .Y(n_781) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_314), .Y(n_1021) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx4_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g444 ( .A(n_318), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g790 ( .A(n_318), .B(n_319), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_319), .Y(n_534) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_319), .Y(n_677) );
INVx1_ASAP7_75t_L g764 ( .A(n_319), .Y(n_764) );
INVx2_ASAP7_75t_SL g972 ( .A(n_319), .Y(n_972) );
INVx2_ASAP7_75t_L g1379 ( .A(n_319), .Y(n_1379) );
AND2x4_ASAP7_75t_L g328 ( .A(n_320), .B(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_333), .B1(n_334), .B2(n_340), .C(n_341), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_322), .A2(n_341), .B1(n_792), .B2(n_793), .C(n_794), .Y(n_791) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
OR2x2_ASAP7_75t_L g667 ( .A(n_324), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_325), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_539) );
AND2x4_ASAP7_75t_L g592 ( .A(n_325), .B(n_328), .Y(n_592) );
AND2x2_ASAP7_75t_L g963 ( .A(n_325), .B(n_328), .Y(n_963) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_SL g339 ( .A(n_327), .Y(n_339) );
INVx1_ASAP7_75t_L g344 ( .A(n_327), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_328), .B(n_331), .Y(n_327) );
BUFx2_ASAP7_75t_L g544 ( .A(n_328), .Y(n_544) );
AND2x4_ASAP7_75t_L g591 ( .A(n_328), .B(n_540), .Y(n_591) );
AND2x4_ASAP7_75t_L g666 ( .A(n_328), .B(n_540), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_328), .Y(n_668) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x6_ASAP7_75t_L g653 ( .A(n_331), .B(n_404), .Y(n_653) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g440 ( .A(n_332), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g463 ( .A(n_332), .B(n_351), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_333), .A2(n_340), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g792 ( .A(n_335), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g540 ( .A(n_337), .Y(n_540) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI31xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_362), .A3(n_426), .B(n_435), .Y(n_345) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221x1_ASAP7_75t_L g796 ( .A1(n_348), .A2(n_431), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_796) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_353), .Y(n_348) );
AND2x4_ASAP7_75t_L g358 ( .A(n_349), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g428 ( .A(n_351), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_351), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g405 ( .A(n_352), .Y(n_405) );
INVx1_ASAP7_75t_L g475 ( .A(n_352), .Y(n_475) );
INVx1_ASAP7_75t_L g805 ( .A(n_353), .Y(n_805) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g478 ( .A(n_354), .Y(n_478) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_355), .Y(n_372) );
INVx3_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
AND2x4_ASAP7_75t_L g360 ( .A(n_356), .B(n_361), .Y(n_360) );
INVx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_SL g808 ( .A1(n_358), .A2(n_809), .B1(n_811), .B2(n_814), .C(n_815), .Y(n_808) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_359), .Y(n_813) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_360), .Y(n_472) );
BUFx3_ASAP7_75t_L g487 ( .A(n_360), .Y(n_487) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_360), .Y(n_495) );
BUFx2_ASAP7_75t_L g558 ( .A(n_360), .Y(n_558) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_373), .B1(n_386), .B2(n_394), .C(n_407), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_370), .B2(n_371), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_365), .A2(n_571), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g387 ( .A(n_366), .Y(n_387) );
INVx2_ASAP7_75t_L g712 ( .A(n_366), .Y(n_712) );
BUFx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g570 ( .A(n_367), .Y(n_570) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g466 ( .A(n_368), .Y(n_466) );
BUFx2_ASAP7_75t_L g725 ( .A(n_368), .Y(n_725) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
AND2x4_ASAP7_75t_L g432 ( .A(n_369), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g649 ( .A(n_372), .Y(n_649) );
INVx4_ASAP7_75t_L g714 ( .A(n_372), .Y(n_714) );
INVx2_ASAP7_75t_SL g1357 ( .A(n_372), .Y(n_1357) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_379), .B2(n_382), .C(n_383), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g419 ( .A(n_375), .Y(n_419) );
INVx2_ASAP7_75t_L g717 ( .A(n_375), .Y(n_717) );
BUFx2_ASAP7_75t_L g944 ( .A(n_375), .Y(n_944) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_376), .B(n_377), .Y(n_396) );
INVx1_ASAP7_75t_L g555 ( .A(n_377), .Y(n_555) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g935 ( .A(n_380), .Y(n_935) );
INVx2_ASAP7_75t_SL g942 ( .A(n_380), .Y(n_942) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_389), .B2(n_393), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_388), .A2(n_397), .B1(n_447), .B2(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g810 ( .A(n_391), .Y(n_810) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g469 ( .A(n_392), .Y(n_469) );
INVx3_ASAP7_75t_L g499 ( .A(n_392), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_400), .B1(n_417), .B2(n_438), .C1(n_442), .C2(n_444), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_398), .B2(n_400), .C(n_401), .Y(n_394) );
INVx2_ASAP7_75t_L g732 ( .A(n_395), .Y(n_732) );
BUFx3_ASAP7_75t_L g937 ( .A(n_395), .Y(n_937) );
BUFx3_ASAP7_75t_L g1057 ( .A(n_395), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_398), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_417), .B(n_418), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_411), .A2(n_419), .B(n_420), .Y(n_418) );
OR2x6_ASAP7_75t_L g807 ( .A(n_411), .B(n_717), .Y(n_807) );
INVx1_ASAP7_75t_L g817 ( .A(n_411), .Y(n_817) );
OR2x6_ASAP7_75t_L g818 ( .A(n_411), .B(n_425), .Y(n_818) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g574 ( .A(n_415), .Y(n_574) );
INVx2_ASAP7_75t_L g821 ( .A(n_415), .Y(n_821) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_416), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g800 ( .A1(n_419), .A2(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g1351 ( .A(n_419), .Y(n_1351) );
NAND2x1_ASAP7_75t_SL g482 ( .A(n_421), .B(n_483), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g816 ( .A(n_421), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_423), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_424), .B(n_483), .Y(n_485) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
CKINVDCx6p67_ASAP7_75t_R g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g812 ( .A(n_429), .Y(n_812) );
INVx3_ASAP7_75t_L g1099 ( .A(n_429), .Y(n_1099) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_432), .Y(n_562) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_432), .Y(n_577) );
INVx1_ASAP7_75t_L g842 ( .A(n_432), .Y(n_842) );
INVx1_ASAP7_75t_L g846 ( .A(n_432), .Y(n_846) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g545 ( .A(n_435), .Y(n_545) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g697 ( .A(n_436), .Y(n_697) );
AND2x2_ASAP7_75t_L g447 ( .A(n_439), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g451 ( .A(n_440), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g823 ( .A(n_440), .B(n_824), .Y(n_823) );
OR2x2_ASAP7_75t_L g825 ( .A(n_440), .B(n_745), .Y(n_825) );
INVx2_ASAP7_75t_L g506 ( .A(n_441), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_441), .B(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g510 ( .A(n_441), .B(n_511), .Y(n_510) );
CKINVDCx6p67_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g657 ( .A(n_444), .Y(n_657) );
INVx2_ASAP7_75t_L g611 ( .A(n_445), .Y(n_611) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g595 ( .A(n_449), .Y(n_595) );
INVx2_ASAP7_75t_SL g780 ( .A(n_449), .Y(n_780) );
CKINVDCx6p67_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_452), .A2(n_517), .B(n_518), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_452), .A2(n_631), .B1(n_634), .B2(n_675), .C(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g529 ( .A(n_453), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_453), .Y(n_538) );
BUFx4f_ASAP7_75t_L g1073 ( .A(n_453), .Y(n_1073) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
OR2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_455), .Y(n_511) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_546), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_488), .C(n_501), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_481), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g491 ( .A(n_463), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g494 ( .A(n_463), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g498 ( .A(n_463), .B(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_463), .A2(n_480), .B1(n_569), .B2(n_576), .Y(n_568) );
AND2x4_ASAP7_75t_L g630 ( .A(n_463), .B(n_469), .Y(n_630) );
AND2x6_ASAP7_75t_L g632 ( .A(n_463), .B(n_487), .Y(n_632) );
AND2x4_ASAP7_75t_L g635 ( .A(n_463), .B(n_574), .Y(n_635) );
AND2x2_ASAP7_75t_L g637 ( .A(n_463), .B(n_492), .Y(n_637) );
AND2x2_ASAP7_75t_L g858 ( .A(n_463), .B(n_492), .Y(n_858) );
AND2x2_ASAP7_75t_L g982 ( .A(n_463), .B(n_492), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B1(n_468), .B2(n_470), .C(n_471), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g930 ( .A(n_466), .Y(n_930) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_466), .Y(n_1054) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g571 ( .A(n_469), .Y(n_571) );
BUFx3_ASAP7_75t_L g947 ( .A(n_469), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_470), .A2(n_522), .B1(n_523), .B2(n_525), .Y(n_521) );
BUFx2_ASAP7_75t_L g851 ( .A(n_472), .Y(n_851) );
OAI33xp33_ASAP7_75t_L g927 ( .A1(n_473), .A2(n_928), .A3(n_934), .B1(n_939), .B2(n_941), .B3(n_945), .Y(n_927) );
OAI33xp33_ASAP7_75t_L g987 ( .A1(n_473), .A2(n_939), .A3(n_988), .B1(n_992), .B2(n_1000), .B3(n_1002), .Y(n_987) );
OAI33xp33_ASAP7_75t_L g1041 ( .A1(n_473), .A2(n_733), .A3(n_1042), .B1(n_1049), .B2(n_1052), .B3(n_1056), .Y(n_1041) );
OAI33xp33_ASAP7_75t_L g1346 ( .A1(n_473), .A2(n_733), .A3(n_1347), .B1(n_1353), .B2(n_1358), .B3(n_1361), .Y(n_1346) );
OAI33xp33_ASAP7_75t_L g1423 ( .A1(n_473), .A2(n_653), .A3(n_1424), .B1(n_1427), .B2(n_1430), .B3(n_1431), .Y(n_1423) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .C(n_480), .Y(n_476) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_478), .Y(n_843) );
INVx1_ASAP7_75t_L g932 ( .A(n_478), .Y(n_932) );
INVx1_ASAP7_75t_L g1055 ( .A(n_478), .Y(n_1055) );
AOI33xp33_ASAP7_75t_L g1088 ( .A1(n_480), .A2(n_560), .A3(n_1089), .B1(n_1091), .B2(n_1095), .B3(n_1097), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_482), .Y(n_924) );
INVx2_ASAP7_75t_L g985 ( .A(n_482), .Y(n_985) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_483), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g550 ( .A(n_483), .B(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g553 ( .A(n_483), .B(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g557 ( .A(n_483), .B(n_558), .Y(n_557) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx4f_ASAP7_75t_L g708 ( .A(n_485), .Y(n_708) );
BUFx4f_ASAP7_75t_L g925 ( .A(n_485), .Y(n_925) );
BUFx3_ASAP7_75t_L g926 ( .A(n_486), .Y(n_926) );
BUFx2_ASAP7_75t_L g986 ( .A(n_486), .Y(n_986) );
BUFx2_ASAP7_75t_L g1345 ( .A(n_486), .Y(n_1345) );
NOR2xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_496), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g707 ( .A(n_491), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_491), .A2(n_635), .B1(n_921), .B2(n_922), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_491), .A2(n_635), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_L g734 ( .A(n_494), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_494), .A2(n_498), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
INVx2_ASAP7_75t_SL g645 ( .A(n_495), .Y(n_645) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_495), .Y(n_839) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g579 ( .A(n_499), .Y(n_579) );
INVx1_ASAP7_75t_L g726 ( .A(n_499), .Y(n_726) );
INVx2_ASAP7_75t_L g998 ( .A(n_499), .Y(n_998) );
INVx2_ASAP7_75t_L g1094 ( .A(n_499), .Y(n_1094) );
INVx2_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
AND2x4_ASAP7_75t_L g656 ( .A(n_500), .B(n_657), .Y(n_656) );
OAI31xp33_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_509), .A3(n_515), .B(n_545), .Y(n_501) );
INVx1_ASAP7_75t_L g862 ( .A(n_503), .Y(n_862) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_504), .A2(n_1023), .B1(n_1024), .B2(n_1025), .C(n_1028), .Y(n_1022) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_505), .A2(n_514), .B1(n_582), .B2(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g745 ( .A(n_505), .Y(n_745) );
BUFx4f_ASAP7_75t_L g1408 ( .A(n_505), .Y(n_1408) );
AND2x4_ASAP7_75t_L g513 ( .A(n_506), .B(n_514), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_506), .A2(n_552), .B1(n_556), .B2(n_585), .C1(n_591), .C2(n_592), .Y(n_584) );
AND2x4_ASAP7_75t_L g662 ( .A(n_506), .B(n_663), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_506), .A2(n_513), .B1(n_603), .B2(n_730), .C(n_744), .Y(n_743) );
INVx4_ASAP7_75t_L g695 ( .A(n_507), .Y(n_695) );
INVx1_ASAP7_75t_L g526 ( .A(n_508), .Y(n_526) );
INVx2_ASAP7_75t_L g758 ( .A(n_508), .Y(n_758) );
INVx6_ASAP7_75t_L g693 ( .A(n_510), .Y(n_693) );
INVx1_ASAP7_75t_L g524 ( .A(n_511), .Y(n_524) );
INVx1_ASAP7_75t_L g587 ( .A(n_511), .Y(n_587) );
INVx2_ASAP7_75t_L g676 ( .A(n_511), .Y(n_676) );
BUFx2_ASAP7_75t_L g1377 ( .A(n_511), .Y(n_1377) );
INVx1_ASAP7_75t_L g1017 ( .A(n_512), .Y(n_1017) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_513), .Y(n_679) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_513), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_513), .A2(n_603), .B1(n_900), .B2(n_901), .C(n_904), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_513), .A2(n_603), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_953) );
INVx1_ASAP7_75t_L g1382 ( .A(n_513), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_513), .Y(n_1405) );
INVx2_ASAP7_75t_SL g597 ( .A(n_514), .Y(n_597) );
AND2x4_ASAP7_75t_L g603 ( .A(n_514), .B(n_544), .Y(n_603) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_514), .Y(n_684) );
BUFx4f_ASAP7_75t_L g749 ( .A(n_514), .Y(n_749) );
INVx1_ASAP7_75t_L g762 ( .A(n_514), .Y(n_762) );
INVx1_ASAP7_75t_L g1385 ( .A(n_514), .Y(n_1385) );
OAI211xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_521), .B(n_527), .C(n_535), .Y(n_515) );
BUFx3_ASAP7_75t_L g753 ( .A(n_519), .Y(n_753) );
INVx1_ASAP7_75t_L g686 ( .A(n_520), .Y(n_686) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .C(n_531), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g866 ( .A1(n_529), .A2(n_854), .B(n_867), .C(n_868), .Y(n_866) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
INVx1_ASAP7_75t_L g1388 ( .A(n_532), .Y(n_1388) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g606 ( .A(n_533), .Y(n_606) );
INVx1_ASAP7_75t_L g763 ( .A(n_533), .Y(n_763) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_533), .Y(n_785) );
INVx2_ASAP7_75t_SL g869 ( .A(n_533), .Y(n_869) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
BUFx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_547), .B(n_614), .Y(n_546) );
INVx1_ASAP7_75t_L g616 ( .A(n_548), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g548 ( .A(n_549), .B(n_559), .C(n_568), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_552), .B1(n_553), .B2(n_556), .C(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g625 ( .A(n_550), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_550), .A2(n_557), .B(n_741), .Y(n_770) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_550), .A2(n_553), .B1(n_557), .B2(n_834), .C(n_835), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_550), .A2(n_553), .B1(n_557), .B2(n_1078), .C(n_1079), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_557), .A2(n_622), .B1(n_623), .B2(n_624), .C(n_626), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_558), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_566), .B2(n_567), .Y(n_559) );
BUFx2_ASAP7_75t_L g837 ( .A(n_560), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_566), .A2(n_605), .B1(n_608), .B2(n_610), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_570), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
INVx2_ASAP7_75t_L g994 ( .A(n_570), .Y(n_994) );
INVx1_ASAP7_75t_L g847 ( .A(n_571), .Y(n_847) );
BUFx3_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
INVx1_ASAP7_75t_L g850 ( .A(n_574), .Y(n_850) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_574), .Y(n_1090) );
BUFx3_ASAP7_75t_L g647 ( .A(n_577), .Y(n_647) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g615 ( .A(n_583), .Y(n_615) );
AOI31xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_593), .A3(n_604), .B(n_612), .Y(n_583) );
OAI221xp5_ASAP7_75t_SL g746 ( .A1(n_586), .A2(n_713), .B1(n_718), .B2(n_747), .C(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g602 ( .A(n_588), .Y(n_602) );
INVx1_ASAP7_75t_L g1027 ( .A(n_588), .Y(n_1027) );
INVx4_ASAP7_75t_L g740 ( .A(n_591), .Y(n_740) );
INVx1_ASAP7_75t_SL g1029 ( .A(n_591), .Y(n_1029) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_591), .A2(n_592), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
INVx2_ASAP7_75t_L g1403 ( .A(n_591), .Y(n_1403) );
AOI222xp33_ASAP7_75t_SL g737 ( .A1(n_592), .A2(n_610), .B1(n_738), .B2(n_739), .C1(n_741), .C2(n_742), .Y(n_737) );
INVx2_ASAP7_75t_SL g865 ( .A(n_592), .Y(n_865) );
AOI322xp5_ASAP7_75t_L g893 ( .A1(n_592), .A2(n_666), .A3(n_894), .B1(n_895), .B2(n_896), .C1(n_897), .C2(n_898), .Y(n_893) );
INVx2_ASAP7_75t_L g1402 ( .A(n_592), .Y(n_1402) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_600), .B(n_603), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx3_ASAP7_75t_L g750 ( .A(n_599), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_603), .A2(n_871), .B1(n_872), .B2(n_873), .C(n_875), .Y(n_870) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_603), .A2(n_1017), .B1(n_1018), .B2(n_1019), .C(n_1020), .Y(n_1016) );
INVx1_ASAP7_75t_L g1075 ( .A(n_603), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_603), .A2(n_1405), .B1(n_1406), .B2(n_1407), .C(n_1409), .Y(n_1404) );
INVx1_ASAP7_75t_L g968 ( .A(n_609), .Y(n_968) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g1086 ( .A(n_612), .Y(n_1086) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .C(n_617), .Y(n_614) );
INVx2_ASAP7_75t_L g699 ( .A(n_618), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_654), .Y(n_619) );
AND4x1_ASAP7_75t_L g620 ( .A(n_621), .B(n_627), .C(n_633), .D(n_638), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_631), .B2(n_632), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_629), .A2(n_632), .B1(n_969), .B2(n_979), .Y(n_978) );
BUFx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx2_ASAP7_75t_L g769 ( .A(n_630), .Y(n_769) );
BUFx2_ASAP7_75t_L g918 ( .A(n_630), .Y(n_918) );
BUFx2_ASAP7_75t_L g1339 ( .A(n_630), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_630), .A2(n_632), .B1(n_1417), .B2(n_1418), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_632), .A2(n_769), .B1(n_853), .B2(n_854), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_632), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_632), .A2(n_1338), .B1(n_1339), .B2(n_1340), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_633) );
INVx1_ASAP7_75t_L g767 ( .A(n_635), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_635), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_635), .A2(n_967), .B1(n_981), .B2(n_982), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_635), .A2(n_982), .B1(n_1102), .B2(n_1103), .C(n_1104), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_635), .A2(n_982), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_635), .A2(n_637), .B1(n_1420), .B2(n_1421), .Y(n_1419) );
AOI33xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .A3(n_646), .B1(n_650), .B2(n_651), .B3(n_652), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_649), .A2(n_1355), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
INVx2_ASAP7_75t_L g733 ( .A(n_652), .Y(n_733) );
AOI33xp33_ASAP7_75t_L g836 ( .A1(n_652), .A2(n_837), .A3(n_838), .B1(n_840), .B2(n_844), .B3(n_848), .Y(n_836) );
INVx6_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx5_ASAP7_75t_L g940 ( .A(n_653), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B(n_659), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_655), .A2(n_765), .B1(n_952), .B2(n_975), .Y(n_951) );
INVx5_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g881 ( .A(n_656), .Y(n_881) );
INVx2_ASAP7_75t_SL g913 ( .A(n_656), .Y(n_913) );
INVx1_ASAP7_75t_L g1366 ( .A(n_656), .Y(n_1366) );
AOI31xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_678), .A3(n_691), .B(n_696), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_664), .C(n_669), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_662), .B(n_909), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_662), .B(n_974), .Y(n_973) );
AOI211xp5_ASAP7_75t_L g1369 ( .A1(n_662), .A2(n_1359), .B(n_1370), .C(n_1372), .Y(n_1369) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_662), .A2(n_1398), .B1(n_1399), .B2(n_1400), .C(n_1401), .Y(n_1397) );
BUFx3_ASAP7_75t_L g1373 ( .A(n_663), .Y(n_1373) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_666), .A2(n_961), .B1(n_962), .B2(n_963), .Y(n_960) );
INVx2_ASAP7_75t_SL g1371 ( .A(n_666), .Y(n_1371) );
INVx1_ASAP7_75t_SL g690 ( .A(n_668), .Y(n_690) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g1068 ( .A(n_673), .Y(n_1068) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g824 ( .A(n_676), .Y(n_824) );
INVx2_ASAP7_75t_L g1066 ( .A(n_676), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_681), .B2(n_687), .C(n_689), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_689), .A2(n_1364), .B1(n_1381), .B2(n_1383), .C(n_1386), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_693), .A2(n_695), .B1(n_878), .B2(n_879), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_693), .A2(n_695), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_693), .A2(n_695), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_693), .A2(n_695), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_693), .A2(n_695), .B1(n_1360), .B2(n_1362), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g1410 ( .A1(n_693), .A2(n_695), .B1(n_1411), .B2(n_1412), .Y(n_1410) );
INVx1_ASAP7_75t_L g765 ( .A(n_696), .Y(n_765) );
AOI31xp33_ASAP7_75t_L g1368 ( .A1(n_696), .A2(n_1369), .A3(n_1380), .B(n_1389), .Y(n_1368) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI21x1_ASAP7_75t_L g795 ( .A1(n_697), .A2(n_796), .B(n_808), .Y(n_795) );
XNOR2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_884), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_829), .B1(n_830), .B2(n_883), .Y(n_701) );
INVx1_ASAP7_75t_L g883 ( .A(n_702), .Y(n_883) );
AO22x2_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_771), .B1(n_772), .B2(n_828), .Y(n_702) );
INVx1_ASAP7_75t_L g828 ( .A(n_703), .Y(n_828) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_735), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g1047 ( .A(n_717), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_717), .A2(n_942), .B1(n_1406), .B2(n_1411), .Y(n_1431) );
INVx3_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_726), .B2(n_727), .Y(n_721) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g1355 ( .A(n_725), .Y(n_1355) );
OAI22xp33_ASAP7_75t_L g1002 ( .A1(n_731), .A2(n_954), .B1(n_958), .B2(n_1003), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1424 ( .A1(n_731), .A2(n_942), .B1(n_1425), .B2(n_1426), .Y(n_1424) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_765), .B(n_766), .Y(n_735) );
NAND4xp25_ASAP7_75t_SL g736 ( .A(n_737), .B(n_743), .C(n_746), .D(n_751), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B1(n_755), .B2(n_759), .C(n_760), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_765), .A2(n_860), .B1(n_880), .B2(n_881), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_765), .A2(n_881), .B1(n_1396), .B2(n_1413), .Y(n_1395) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NOR4xp75_ASAP7_75t_L g773 ( .A(n_774), .B(n_795), .C(n_822), .D(n_826), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_791), .Y(n_774) );
AOI33xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .A3(n_782), .B1(n_783), .B2(n_788), .B3(n_790), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g971 ( .A(n_785), .Y(n_971) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g874 ( .A(n_787), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_803), .B(n_807), .Y(n_799) );
INVx1_ASAP7_75t_L g1096 ( .A(n_805), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
XNOR2x1_ASAP7_75t_L g830 ( .A(n_831), .B(n_882), .Y(n_830) );
NAND2x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_859), .Y(n_831) );
AND4x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_836), .C(n_852), .D(n_855), .Y(n_832) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g1092 ( .A(n_842), .Y(n_1092) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_870), .C(n_877), .Y(n_860) );
AOI21xp5_ASAP7_75t_SL g861 ( .A1(n_862), .A2(n_863), .B(n_864), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B1(n_1007), .B2(n_1008), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_948), .B2(n_949), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
XNOR2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_914), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_910), .B1(n_912), .B2(n_913), .Y(n_891) );
NAND4xp25_ASAP7_75t_L g892 ( .A(n_893), .B(n_899), .C(n_905), .D(n_908), .Y(n_892) );
OAI22xp33_ASAP7_75t_L g941 ( .A1(n_900), .A2(n_906), .B1(n_942), .B2(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_907), .A2(n_909), .B1(n_929), .B2(n_946), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g1011 ( .A1(n_910), .A2(n_913), .B1(n_1012), .B2(n_1030), .Y(n_1011) );
CKINVDCx8_ASAP7_75t_R g910 ( .A(n_911), .Y(n_910) );
NOR3xp33_ASAP7_75t_SL g914 ( .A(n_915), .B(n_923), .C(n_927), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_920), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_931), .B1(n_932), .B2(n_933), .Y(n_928) );
BUFx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1427 ( .A1(n_932), .A2(n_993), .B1(n_1428), .B2(n_1429), .Y(n_1427) );
OAI22xp33_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_936), .B1(n_937), .B2(n_938), .Y(n_934) );
CKINVDCx8_ASAP7_75t_R g939 ( .A(n_940), .Y(n_939) );
OAI22xp33_ASAP7_75t_L g988 ( .A1(n_942), .A2(n_989), .B1(n_990), .B2(n_991), .Y(n_988) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g990 ( .A(n_944), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_946), .A2(n_1001), .B1(n_1398), .B2(n_1412), .Y(n_1430) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_SL g948 ( .A(n_949), .Y(n_948) );
XNOR2x1_ASAP7_75t_L g949 ( .A(n_950), .B(n_1006), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_976), .Y(n_950) );
NAND5xp2_ASAP7_75t_L g952 ( .A(n_953), .B(n_957), .C(n_960), .D(n_964), .E(n_973), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_959), .A2(n_974), .B1(n_998), .B2(n_1001), .Y(n_1000) );
OAI221xp5_ASAP7_75t_SL g964 ( .A1(n_965), .A2(n_967), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
NOR3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_983), .C(n_987), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_980), .Y(n_977) );
INVx2_ASAP7_75t_SL g984 ( .A(n_985), .Y(n_984) );
INVx2_ASAP7_75t_L g1040 ( .A(n_985), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_993), .A2(n_995), .B1(n_996), .B2(n_999), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g1001 ( .A(n_994), .Y(n_1001) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx2_ASAP7_75t_SL g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_1005), .A2(n_1014), .B1(n_1018), .B2(n_1057), .Y(n_1056) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
XOR2x2_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1060), .Y(n_1008) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1010), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1031), .Y(n_1010) );
NAND3xp33_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1016), .C(n_1022), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1015), .A2(n_1023), .B1(n_1053), .B2(n_1055), .Y(n_1052) );
NOR3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1039), .C(n_1041), .Y(n_1031) );
NAND2xp5_ASAP7_75t_SL g1032 ( .A(n_1033), .B(n_1036), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1045), .B1(n_1046), .B2(n_1048), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_1043), .Y(n_1348) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1061), .Y(n_1106) );
NAND4xp75_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .C(n_1087), .D(n_1101), .Y(n_1061) );
OAI31xp33_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1076), .A3(n_1085), .B(n_1086), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B1(n_1068), .B2(n_1069), .Y(n_1065) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1068), .Y(n_1374) );
OAI21xp33_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1072), .B(n_1074), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1073), .Y(n_1082) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1073), .Y(n_1376) );
OAI211xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B(n_1083), .C(n_1084), .Y(n_1080) );
AND2x2_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1100), .Y(n_1087) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
OAI21xp33_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1116), .B(n_1331), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
BUFx3_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1110), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1114), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1111), .B(n_1114), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1439 ( .A(n_1111), .Y(n_1439) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_1112), .B(n_1114), .Y(n_1132) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1113), .B(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1115), .Y(n_1125) );
NOR2x1_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1281), .Y(n_1116) );
NAND3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1214), .C(n_1258), .Y(n_1117) );
AOI211xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1140), .B(n_1179), .C(n_1209), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1119), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1119), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1133), .Y(n_1119) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1120), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1120), .B(n_1177), .Y(n_1199) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1120), .Y(n_1213) );
BUFx6f_ASAP7_75t_L g1228 ( .A(n_1120), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1120), .B(n_1172), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1131), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1126), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1124), .B(n_1127), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1438 ( .A(n_1125), .Y(n_1438) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_1126), .B(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1127), .B(n_1130), .Y(n_1171) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1132), .Y(n_1138) );
CKINVDCx6p67_ASAP7_75t_R g1195 ( .A(n_1133), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1133), .B(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1133), .B(n_1213), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1133), .B(n_1249), .Y(n_1248) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_1133), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1133), .B(n_1326), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1133), .B(n_1191), .Y(n_1330) );
OR2x6_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1134), .B(n_1135), .Y(n_1233) );
OAI22xp5_ASAP7_75t_SL g1135 ( .A1(n_1136), .A2(n_1137), .B1(n_1138), .B2(n_1139), .Y(n_1135) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1138), .Y(n_1164) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1138), .Y(n_1202) );
A2O1A1Ixp33_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1155), .B(n_1161), .C(n_1175), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1329 ( .A(n_1141), .B(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1147), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g1157 ( .A(n_1143), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1143), .B(n_1158), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1143), .B(n_1198), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1143), .B(n_1183), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1143), .B(n_1236), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1143), .B(n_1198), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1143), .B(n_1162), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1143), .B(n_1316), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1143), .B(n_1231), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1143), .B(n_1316), .Y(n_1323) );
AND2x4_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1145), .Y(n_1143) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1147), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1147), .B(n_1157), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1151), .Y(n_1147) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1148), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1148), .B(n_1152), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1152), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1152), .B(n_1159), .Y(n_1231) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1152), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1154), .Y(n_1152) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1156), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1156), .B(n_1181), .Y(n_1226) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_1156), .A2(n_1249), .B1(n_1266), .B2(n_1290), .C(n_1292), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1156), .B(n_1223), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1158), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1157), .B(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1157), .B(n_1188), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1157), .B(n_1230), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1157), .B(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1157), .B(n_1231), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1157), .B(n_1163), .Y(n_1272) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1158), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1158), .B(n_1275), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1158), .B(n_1280), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1160), .Y(n_1158) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1159), .Y(n_1198) );
OAI322xp33_ASAP7_75t_L g1234 ( .A1(n_1161), .A2(n_1235), .A3(n_1237), .B1(n_1239), .B2(n_1240), .C1(n_1241), .C2(n_1243), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1172), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1176 ( .A(n_1162), .B(n_1177), .Y(n_1176) );
BUFx3_ASAP7_75t_L g1181 ( .A(n_1162), .Y(n_1181) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_1162), .Y(n_1189) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_1162), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1162), .B(n_1266), .Y(n_1265) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_1163), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1163), .B(n_1177), .Y(n_1249) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1167), .B1(n_1169), .B2(n_1170), .Y(n_1165) );
BUFx3_ASAP7_75t_L g1205 ( .A(n_1167), .Y(n_1205) );
BUFx6f_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1171), .Y(n_1208) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1172), .Y(n_1177) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1172), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1172), .B(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1172), .Y(n_1266) );
NAND3xp33_ASAP7_75t_L g1273 ( .A(n_1172), .B(n_1274), .C(n_1276), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1176), .B(n_1183), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1177), .B(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1177), .B(n_1192), .Y(n_1269) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1178), .Y(n_1218) );
A2O1A1Ixp33_ASAP7_75t_L g1296 ( .A1(n_1178), .A2(n_1233), .B(n_1262), .C(n_1297), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1178), .B(n_1302), .Y(n_1301) );
OAI211xp5_ASAP7_75t_L g1321 ( .A1(n_1178), .A2(n_1322), .B(n_1324), .C(n_1327), .Y(n_1321) );
OAI221xp5_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1184), .B1(n_1186), .B2(n_1191), .C(n_1193), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
NOR3xp33_ASAP7_75t_L g1200 ( .A(n_1181), .B(n_1198), .C(n_1201), .Y(n_1200) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1181), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1181), .B(n_1269), .Y(n_1308) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1183), .Y(n_1244) );
A2O1A1Ixp33_ASAP7_75t_L g1294 ( .A1(n_1184), .A2(n_1235), .B(n_1295), .C(n_1296), .Y(n_1294) );
OAI211xp5_ASAP7_75t_SL g1283 ( .A1(n_1185), .A2(n_1284), .B(n_1286), .C(n_1289), .Y(n_1283) );
INVx3_ASAP7_75t_L g1304 ( .A(n_1185), .Y(n_1304) );
AOI21xp33_ASAP7_75t_L g1209 ( .A1(n_1186), .A2(n_1210), .B(n_1212), .Y(n_1209) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1189), .B(n_1197), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g1211 ( .A(n_1189), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1189), .B(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1189), .B(n_1315), .Y(n_1314) );
INVxp67_ASAP7_75t_L g1326 ( .A(n_1189), .Y(n_1326) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1191), .Y(n_1242) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1191), .Y(n_1327) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1196), .B1(n_1199), .B2(n_1200), .Y(n_1193) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1194), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1195), .B(n_1225), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1195), .B(n_1199), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1195), .B(n_1213), .Y(n_1313) );
NAND2xp5_ASAP7_75t_SL g1318 ( .A(n_1195), .B(n_1269), .Y(n_1318) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1197), .Y(n_1240) );
AOI222xp33_ASAP7_75t_L g1286 ( .A1(n_1198), .A2(n_1231), .B1(n_1261), .B2(n_1269), .C1(n_1287), .C2(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1198), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1199), .B(n_1238), .Y(n_1250) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1199), .Y(n_1311) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1201), .Y(n_1257) );
OAI22xp33_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1205), .B1(n_1206), .B2(n_1207), .Y(n_1203) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1211), .Y(n_1300) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1212), .Y(n_1276) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1213), .Y(n_1239) );
OAI31xp33_ASAP7_75t_SL g1214 ( .A1(n_1215), .A2(n_1224), .A3(n_1227), .B(n_1254), .Y(n_1214) );
OAI222xp33_ASAP7_75t_L g1215 ( .A1(n_1216), .A2(n_1217), .B1(n_1218), .B2(n_1219), .C1(n_1220), .C2(n_1222), .Y(n_1215) );
OAI321xp33_ASAP7_75t_L g1298 ( .A1(n_1217), .A2(n_1245), .A3(n_1295), .B1(n_1299), .B2(n_1300), .C(n_1301), .Y(n_1298) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1220), .A2(n_1260), .B1(n_1263), .B2(n_1264), .Y(n_1259) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1221), .B(n_1285), .Y(n_1328) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1223), .B(n_1237), .Y(n_1285) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
OAI211xp5_ASAP7_75t_SL g1227 ( .A1(n_1228), .A2(n_1229), .B(n_1232), .C(n_1251), .Y(n_1227) );
CKINVDCx14_ASAP7_75t_R g1288 ( .A(n_1228), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1231), .B(n_1272), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1234), .B1(n_1246), .B2(n_1247), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1235), .B(n_1238), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1236), .B(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1236), .Y(n_1291) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1238), .B(n_1262), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1242), .B(n_1280), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1245), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1244), .B(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1246), .Y(n_1263) );
NAND2xp33_ASAP7_75t_SL g1247 ( .A(n_1248), .B(n_1250), .Y(n_1247) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1249), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1253), .Y(n_1251) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1253), .Y(n_1299) );
OAI21xp33_ASAP7_75t_L g1281 ( .A1(n_1254), .A2(n_1282), .B(n_1305), .Y(n_1281) );
INVx3_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
AOI21xp5_ASAP7_75t_L g1258 ( .A1(n_1255), .A2(n_1259), .B(n_1267), .Y(n_1258) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1278 ( .A(n_1263), .B(n_1279), .Y(n_1278) );
OAI211xp5_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1270), .B(n_1273), .C(n_1277), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
AOI211xp5_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1293), .B(n_1294), .C(n_1298), .Y(n_1282) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
NOR3xp33_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1317), .C(n_1329), .Y(n_1305) );
OAI221xp5_ASAP7_75t_SL g1306 ( .A1(n_1307), .A2(n_1308), .B1(n_1309), .B2(n_1311), .C(n_1312), .Y(n_1306) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
OAI211xp5_ASAP7_75t_SL g1317 ( .A1(n_1318), .A2(n_1319), .B(n_1321), .C(n_1328), .Y(n_1317) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx3_ASAP7_75t_SL g1332 ( .A(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1365), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1344), .C(n_1346), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1341), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g1375 ( .A1(n_1340), .A2(n_1342), .B1(n_1376), .B2(n_1377), .C(n_1378), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B1(n_1350), .B2(n_1352), .Y(n_1347) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_1348), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1361) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1351), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1355), .B1(n_1356), .B2(n_1357), .Y(n_1353) );
AOI21xp5_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1367), .B(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
BUFx2_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1393), .Y(n_1433) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1414), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1404), .C(n_1410), .Y(n_1396) );
NOR3xp33_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1422), .C(n_1423), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1419), .Y(n_1415) );
A2O1A1Ixp33_ASAP7_75t_L g1436 ( .A1(n_1435), .A2(n_1437), .B(n_1439), .C(n_1440), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
endmodule