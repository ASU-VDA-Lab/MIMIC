module fake_netlist_6_1918_n_2657 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2657);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2657;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2307;
wire n_2069;
wire n_2362;
wire n_684;
wire n_2539;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_811;
wire n_683;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_1390;
wire n_906;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_1303;
wire n_761;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g577 ( 
.A(n_415),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_48),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_111),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_194),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_568),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_561),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_95),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_311),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_557),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_373),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_492),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_312),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_536),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_176),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_532),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_397),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_527),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_428),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_338),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_241),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_105),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_516),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_325),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_410),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_484),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_376),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_186),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_369),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_269),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_355),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_86),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_21),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_43),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_67),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_258),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_563),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_393),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_368),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_213),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_265),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_472),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_540),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_246),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_26),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_350),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_304),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_178),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_332),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_266),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_330),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_406),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_145),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_68),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_16),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_423),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_411),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_555),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_18),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_467),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_248),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_250),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_84),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_512),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_181),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_33),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_362),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_533),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_111),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_203),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_565),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_232),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_569),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_157),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_58),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_172),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_570),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_293),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_265),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_482),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_376),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_226),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_160),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_298),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_261),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_403),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_164),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_346),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_96),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_268),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_337),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_105),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_258),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_393),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_448),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_115),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_515),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_477),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_163),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_374),
.Y(n_679)
);

INVxp33_ASAP7_75t_SL g680 ( 
.A(n_275),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_172),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_409),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_165),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_168),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_416),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_116),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_85),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_283),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_28),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_146),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_435),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_498),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_289),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_101),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_342),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_391),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_551),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_424),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_23),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_106),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_417),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_439),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_462),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_117),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_66),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_204),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_243),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_330),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_394),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_181),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_449),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_552),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_210),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_575),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_79),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_547),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_7),
.Y(n_717)
);

BUFx10_ASAP7_75t_L g718 ( 
.A(n_207),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_405),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_271),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_152),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_554),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_52),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_356),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_236),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_529),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_50),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_34),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_59),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_107),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_413),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_35),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_441),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_143),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_236),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_125),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_217),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_494),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_161),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_132),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_264),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_108),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_378),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_152),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_333),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_132),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_136),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_537),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_96),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_545),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_344),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_3),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_479),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_151),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_375),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_457),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_440),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_143),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_412),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_20),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_466),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_78),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_574),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_232),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_411),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_89),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_89),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_399),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_359),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_336),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_302),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_471),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_371),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_193),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_507),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_168),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_442),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_451),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_163),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_33),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_212),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_18),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_7),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_289),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_307),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_196),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_446),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_434),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_548),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_511),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_524),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_546),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_207),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_378),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_407),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_175),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_503),
.Y(n_797)
);

BUFx8_ASAP7_75t_SL g798 ( 
.A(n_74),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_387),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_553),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_86),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_307),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_408),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_25),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_126),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_323),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_220),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_120),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_48),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_184),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_305),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_437),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_383),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_58),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_193),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_653),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_653),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_764),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_729),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_620),
.Y(n_820)
);

BUFx5_ASAP7_75t_L g821 ( 
.A(n_577),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_760),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_811),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_770),
.Y(n_827)
);

CKINVDCx16_ASAP7_75t_R g828 ( 
.A(n_701),
.Y(n_828)
);

INVxp33_ASAP7_75t_SL g829 ( 
.A(n_632),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_785),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_785),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_628),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_628),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_798),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_605),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_606),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_611),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_628),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_628),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_628),
.Y(n_840)
);

INVxp33_ASAP7_75t_SL g841 ( 
.A(n_578),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_714),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_610),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_578),
.Y(n_844)
);

CKINVDCx16_ASAP7_75t_R g845 ( 
.A(n_748),
.Y(n_845)
);

INVxp67_ASAP7_75t_SL g846 ( 
.A(n_714),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_700),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_700),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_702),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_637),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_700),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_700),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_612),
.Y(n_853)
);

CKINVDCx16_ASAP7_75t_R g854 ( 
.A(n_605),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_797),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_605),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_700),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_594),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_584),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_590),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_592),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_602),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_596),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_614),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_597),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_598),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_579),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_600),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_660),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_618),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_655),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_622),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_623),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_618),
.Y(n_874)
);

INVxp33_ASAP7_75t_SL g875 ( 
.A(n_579),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_640),
.Y(n_876)
);

INVxp33_ASAP7_75t_SL g877 ( 
.A(n_580),
.Y(n_877)
);

CKINVDCx14_ASAP7_75t_R g878 ( 
.A(n_618),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_646),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_648),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_651),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_655),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_615),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_658),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_661),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_662),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_670),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_683),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_616),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_684),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_688),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_694),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_609),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_667),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_621),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_699),
.Y(n_896)
);

CKINVDCx16_ASAP7_75t_R g897 ( 
.A(n_655),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_691),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_617),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_638),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_602),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_736),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_737),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_580),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_742),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_665),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_583),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_644),
.Y(n_910)
);

INVxp33_ASAP7_75t_L g911 ( 
.A(n_607),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_624),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_665),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_780),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_720),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_839),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_839),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_828),
.B(n_650),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_845),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_858),
.B(n_772),
.Y(n_920)
);

BUFx12f_ASAP7_75t_L g921 ( 
.A(n_834),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_846),
.B(n_772),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_840),
.Y(n_923)
);

CKINVDCx6p67_ASAP7_75t_R g924 ( 
.A(n_854),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_867),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_842),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_840),
.Y(n_927)
);

AND2x6_ASAP7_75t_L g928 ( 
.A(n_898),
.B(n_691),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_836),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_832),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_898),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_849),
.B(n_636),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_898),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_833),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_855),
.B(n_636),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_898),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_898),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_821),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_866),
.B(n_674),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_842),
.B(n_607),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_834),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_838),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_847),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_837),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_821),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_848),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_851),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_820),
.B(n_591),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_857),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_862),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_862),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_816),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_902),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_902),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_870),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_821),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_821),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_911),
.B(n_626),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_870),
.Y(n_960)
);

INVx5_ASAP7_75t_L g961 ( 
.A(n_874),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_821),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_893),
.B(n_703),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_859),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_895),
.B(n_703),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_860),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_821),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_821),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_874),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_817),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_837),
.B(n_680),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_861),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_853),
.B(n_680),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_853),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_864),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_864),
.B(n_581),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_871),
.B(n_897),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_863),
.Y(n_978)
);

NOR2x1_ASAP7_75t_L g979 ( 
.A(n_819),
.B(n_775),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_883),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_920),
.B(n_901),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_933),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_944),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_959),
.B(n_911),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_933),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_926),
.B(n_775),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_919),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_923),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_976),
.B(n_841),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_923),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_952),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_916),
.A2(n_910),
.B(n_790),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_948),
.B(n_841),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_952),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_964),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_952),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_964),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_952),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_952),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_926),
.B(n_790),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_939),
.B(n_652),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_929),
.A2(n_745),
.B1(n_774),
.B2(n_724),
.Y(n_1002)
);

OA21x2_ASAP7_75t_L g1003 ( 
.A1(n_916),
.A2(n_697),
.B(n_677),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_964),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_964),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_953),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_920),
.B(n_878),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_953),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_934),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_945),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_939),
.B(n_965),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_944),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_939),
.B(n_711),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_970),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_933),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_933),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_822),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_920),
.B(n_823),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_940),
.B(n_825),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_939),
.B(n_691),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_964),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_934),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_965),
.B(n_878),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_942),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_965),
.B(n_883),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_965),
.B(n_889),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_942),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_966),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_919),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_940),
.B(n_826),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_933),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_966),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_949),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_949),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_937),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_950),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_966),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_971),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_924),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_967),
.A2(n_726),
.B(n_722),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_937),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_950),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_970),
.B(n_827),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_937),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_966),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_937),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_973),
.B(n_875),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_980),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_966),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_972),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_917),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_972),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_972),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_922),
.B(n_889),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_932),
.B(n_830),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_967),
.A2(n_792),
.B(n_831),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_972),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_972),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_937),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_917),
.Y(n_1060)
);

OAI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_918),
.A2(n_856),
.B1(n_829),
.B2(n_668),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_927),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_943),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_927),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_943),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_975),
.B(n_875),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_930),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1051),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1051),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1011),
.B(n_975),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_984),
.B(n_975),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1038),
.B(n_975),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_984),
.B(n_956),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_993),
.B(n_956),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_1011),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1060),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1047),
.B(n_877),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_989),
.B(n_877),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_1010),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1051),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_1006),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1060),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1011),
.B(n_956),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1067),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1067),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1011),
.Y(n_1086)
);

OAI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_981),
.A2(n_935),
.B1(n_977),
.B2(n_963),
.Y(n_1087)
);

NOR2x1p5_ASAP7_75t_L g1088 ( 
.A(n_983),
.B(n_924),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1066),
.B(n_956),
.Y(n_1089)
);

CKINVDCx6p67_ASAP7_75t_R g1090 ( 
.A(n_987),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1062),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1062),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1048),
.Y(n_1093)
);

NOR2x1p5_ASAP7_75t_L g1094 ( 
.A(n_1012),
.B(n_974),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1064),
.Y(n_1095)
);

INVx8_ASAP7_75t_L g1096 ( 
.A(n_1020),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_1019),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1064),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1022),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1009),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_988),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1025),
.B(n_960),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_1019),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1022),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1006),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1022),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_SL g1107 ( 
.A(n_1026),
.B(n_789),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1007),
.B(n_960),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1043),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1061),
.B(n_960),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1001),
.B(n_967),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_988),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1043),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_987),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_988),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_990),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_990),
.Y(n_1117)
);

INVxp33_ASAP7_75t_L g1118 ( 
.A(n_1030),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1024),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1010),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1009),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1027),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1027),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1033),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1017),
.Y(n_1125)
);

AO22x2_ASAP7_75t_L g1126 ( 
.A1(n_1001),
.A2(n_856),
.B1(n_626),
.B2(n_664),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1033),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1034),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1034),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1001),
.B(n_960),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1024),
.Y(n_1131)
);

OAI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1023),
.A2(n_869),
.B1(n_912),
.B2(n_900),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1024),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1036),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1010),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1008),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1036),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1036),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1008),
.B(n_960),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_1018),
.B(n_1001),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1042),
.Y(n_1141)
);

AND2x2_ASAP7_75t_SL g1142 ( 
.A(n_1013),
.B(n_691),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1008),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1042),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1042),
.Y(n_1145)
);

CKINVDCx6p67_ASAP7_75t_R g1146 ( 
.A(n_1039),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1013),
.B(n_961),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

NOR2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1014),
.B(n_974),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_992),
.A2(n_958),
.B(n_957),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_992),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_1029),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_991),
.Y(n_1153)
);

INVxp33_ASAP7_75t_L g1154 ( 
.A(n_1030),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_991),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1017),
.B(n_867),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1013),
.B(n_961),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_986),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1014),
.B(n_961),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1014),
.B(n_961),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_986),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_994),
.Y(n_1163)
);

NOR2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1018),
.B(n_921),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_994),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_986),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_986),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1000),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_996),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1013),
.B(n_961),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_995),
.A2(n_958),
.B(n_957),
.Y(n_1171)
);

XNOR2xp5_ASAP7_75t_L g1172 ( 
.A(n_1002),
.B(n_836),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_985),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_999),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_985),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_996),
.Y(n_1176)
);

INVxp33_ASAP7_75t_L g1177 ( 
.A(n_1002),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_998),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_912),
.B1(n_900),
.B2(n_909),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_999),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_999),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1003),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1003),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1003),
.Y(n_1185)
);

INVx11_ASAP7_75t_L g1186 ( 
.A(n_1020),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1003),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1000),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_982),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1010),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_995),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1055),
.B(n_824),
.C(n_818),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_1020),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_982),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1000),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1055),
.B(n_905),
.C(n_844),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_985),
.Y(n_1197)
);

AND3x2_ASAP7_75t_L g1198 ( 
.A(n_1049),
.B(n_751),
.C(n_835),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_997),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_982),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_997),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1004),
.B(n_961),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1004),
.Y(n_1203)
);

XNOR2x2_ASAP7_75t_L g1204 ( 
.A(n_1172),
.B(n_599),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1082),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1082),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1091),
.Y(n_1207)
);

INVx4_ASAP7_75t_SL g1208 ( 
.A(n_1140),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1114),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1091),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1095),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1152),
.Y(n_1213)
);

CKINVDCx16_ASAP7_75t_R g1214 ( 
.A(n_1172),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1125),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1068),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_1192),
.B(n_1196),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1068),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1156),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1069),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1078),
.B(n_921),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1077),
.B(n_909),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1090),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1098),
.Y(n_1224)
);

XOR2xp5_ASAP7_75t_L g1225 ( 
.A(n_1180),
.B(n_843),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1098),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1191),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_R g1228 ( 
.A(n_1093),
.B(n_829),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1081),
.B(n_978),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1069),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1086),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1090),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1191),
.Y(n_1233)
);

OR2x6_ASAP7_75t_SL g1234 ( 
.A(n_1156),
.B(n_583),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1093),
.B(n_941),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1097),
.B(n_908),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1076),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1076),
.Y(n_1238)
);

XOR2xp5_ASAP7_75t_L g1239 ( 
.A(n_1177),
.B(n_843),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1092),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1118),
.B(n_913),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1097),
.B(n_882),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1080),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1092),
.B(n_1005),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1084),
.B(n_1057),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1086),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1086),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1100),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1100),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1121),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1075),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1075),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1081),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1085),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1072),
.B(n_925),
.Y(n_1255)
);

XNOR2xp5_ASAP7_75t_L g1256 ( 
.A(n_1164),
.B(n_850),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1118),
.B(n_1154),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1080),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1158),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1146),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1103),
.B(n_1057),
.Y(n_1261)
);

INVxp33_ASAP7_75t_L g1262 ( 
.A(n_1154),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1105),
.B(n_978),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1166),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1103),
.B(n_1021),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1109),
.B(n_850),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1188),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1198),
.Y(n_1268)
);

XOR2xp5_ASAP7_75t_L g1269 ( 
.A(n_1177),
.B(n_894),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1142),
.B(n_941),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1195),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1122),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1122),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1123),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1123),
.Y(n_1275)
);

AND2x2_ASAP7_75t_SL g1276 ( 
.A(n_1142),
.B(n_627),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1146),
.Y(n_1278)
);

XOR2xp5_ASAP7_75t_L g1279 ( 
.A(n_1071),
.B(n_894),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1124),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1127),
.Y(n_1281)
);

XOR2xp5_ASAP7_75t_L g1282 ( 
.A(n_1132),
.B(n_915),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1127),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1116),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1113),
.B(n_915),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1116),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1107),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1105),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1128),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1128),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1117),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1129),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1131),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1136),
.Y(n_1295)
);

AND2x2_ASAP7_75t_SL g1296 ( 
.A(n_1070),
.B(n_627),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1131),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1107),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1087),
.B(n_925),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1136),
.B(n_969),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1143),
.B(n_1162),
.Y(n_1301)
);

CKINVDCx14_ASAP7_75t_R g1302 ( 
.A(n_1140),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1199),
.Y(n_1303)
);

XOR2xp5_ASAP7_75t_L g1304 ( 
.A(n_1126),
.B(n_804),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1201),
.B(n_925),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1149),
.B(n_979),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1162),
.B(n_925),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1135),
.B(n_806),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1133),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1110),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1133),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1134),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1167),
.B(n_979),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1134),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1137),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1137),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1138),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1167),
.B(n_1021),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1141),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1173),
.Y(n_1322)
);

XNOR2xp5_ASAP7_75t_L g1323 ( 
.A(n_1094),
.B(n_581),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1141),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1173),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1144),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1088),
.Y(n_1327)
);

XOR2xp5_ASAP7_75t_L g1328 ( 
.A(n_1126),
.B(n_613),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1135),
.B(n_1063),
.Y(n_1329)
);

CKINVDCx16_ASAP7_75t_R g1330 ( 
.A(n_1140),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1126),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1144),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1145),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1168),
.B(n_1028),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1168),
.B(n_1028),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1101),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1101),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1112),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1148),
.B(n_1032),
.Y(n_1340)
);

XOR2x2_ASAP7_75t_L g1341 ( 
.A(n_1074),
.B(n_673),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1112),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1148),
.B(n_1058),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1115),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1115),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1173),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1153),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1151),
.B(n_1037),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1155),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1126),
.B(n_665),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1099),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1155),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1140),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1159),
.B(n_1045),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1165),
.Y(n_1355)
);

INVxp33_ASAP7_75t_L g1356 ( 
.A(n_1073),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1165),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1140),
.B(n_1037),
.Y(n_1358)
);

AND2x6_ASAP7_75t_L g1359 ( 
.A(n_1159),
.B(n_1050),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1176),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1189),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1104),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1176),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1178),
.Y(n_1364)
);

XOR2xp5_ASAP7_75t_L g1365 ( 
.A(n_1108),
.B(n_619),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1140),
.B(n_718),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1178),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1104),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1104),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1106),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1106),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1106),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1163),
.B(n_718),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1163),
.B(n_718),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1111),
.B(n_1119),
.Y(n_1375)
);

XOR2xp5_ASAP7_75t_L g1376 ( 
.A(n_1102),
.B(n_634),
.Y(n_1376)
);

XOR2xp5_ASAP7_75t_L g1377 ( 
.A(n_1083),
.B(n_642),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1119),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1173),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1119),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1173),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1169),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1169),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1179),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_1175),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1181),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1179),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1135),
.B(n_1052),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1189),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1182),
.B(n_1052),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1183),
.B(n_773),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1309),
.B(n_1079),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1257),
.B(n_773),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1213),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1227),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1216),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1322),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1219),
.B(n_1183),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1218),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1233),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1222),
.B(n_1214),
.C(n_1305),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1309),
.B(n_1079),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1237),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1238),
.B(n_1190),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1219),
.B(n_1184),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1240),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1231),
.B(n_1200),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1231),
.B(n_1200),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1222),
.B(n_1200),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1205),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1375),
.B(n_1174),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1262),
.B(n_1174),
.Y(n_1412)
);

AND2x6_ASAP7_75t_SL g1413 ( 
.A(n_1235),
.B(n_781),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1270),
.B(n_1120),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1215),
.B(n_1174),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1215),
.B(n_1194),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1270),
.B(n_1120),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1242),
.B(n_1266),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1276),
.A2(n_1185),
.B1(n_1187),
.B2(n_1184),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_SL g1420 ( 
.A(n_1235),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1285),
.B(n_1241),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1236),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1279),
.B(n_1253),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1254),
.B(n_1276),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1217),
.A2(n_754),
.B1(n_769),
.B2(n_749),
.C(n_746),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1206),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1288),
.B(n_1120),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1207),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1288),
.B(n_1120),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1255),
.B(n_1194),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1210),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1303),
.B(n_1120),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1385),
.B(n_1193),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1373),
.B(n_773),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1228),
.B(n_629),
.C(n_625),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1306),
.B(n_1185),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1261),
.B(n_1187),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1311),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1228),
.Y(n_1439)
);

AND2x4_ASAP7_75t_SL g1440 ( 
.A(n_1301),
.B(n_1175),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_SL g1441 ( 
.A(n_1235),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1261),
.B(n_1020),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1220),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1230),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1255),
.A2(n_1299),
.B1(n_1298),
.B2(n_1287),
.Y(n_1445)
);

INVx8_ASAP7_75t_L g1446 ( 
.A(n_1358),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1211),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1375),
.B(n_1175),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1299),
.A2(n_1130),
.B1(n_1157),
.B2(n_1147),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1243),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1338),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1305),
.B(n_1089),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1340),
.A2(n_1096),
.B(n_1193),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1295),
.Y(n_1454)
);

NOR2xp67_ASAP7_75t_L g1455 ( 
.A(n_1223),
.B(n_1139),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1308),
.B(n_1193),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1265),
.B(n_1020),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1265),
.B(n_1020),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1391),
.B(n_1053),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1239),
.B(n_786),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1229),
.B(n_1175),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1212),
.B(n_1053),
.Y(n_1462)
);

NOR2xp67_ASAP7_75t_SL g1463 ( 
.A(n_1330),
.B(n_1175),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1229),
.B(n_1197),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1344),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1263),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1224),
.B(n_1197),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1296),
.A2(n_1096),
.B1(n_1161),
.B2(n_1160),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1226),
.B(n_1197),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1374),
.B(n_801),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1294),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1244),
.B(n_1197),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_SL g1473 ( 
.A(n_1268),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1331),
.A2(n_1096),
.B1(n_1170),
.B2(n_1202),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1353),
.B(n_1197),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1263),
.B(n_582),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1341),
.B(n_865),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1297),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1244),
.B(n_1248),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1345),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1234),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1322),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1259),
.B(n_982),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1264),
.B(n_1267),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1347),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_SL g1486 ( 
.A(n_1322),
.B(n_582),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1389),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1269),
.B(n_1171),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1249),
.B(n_1150),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1221),
.B(n_1356),
.Y(n_1490)
);

BUFx12f_ASAP7_75t_L g1491 ( 
.A(n_1232),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1350),
.B(n_868),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1366),
.A2(n_656),
.B1(n_659),
.B2(n_647),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1349),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1307),
.B(n_872),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1250),
.B(n_1150),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1352),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1325),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1282),
.B(n_1186),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_SL g1500 ( 
.A(n_1358),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1271),
.B(n_1059),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1377),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1221),
.B(n_585),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1355),
.Y(n_1504)
);

NOR2xp67_ASAP7_75t_L g1505 ( 
.A(n_1260),
.B(n_676),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1304),
.B(n_1186),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_L g1507 ( 
.A(n_1325),
.B(n_685),
.Y(n_1507)
);

AO22x1_ASAP7_75t_L g1508 ( 
.A1(n_1327),
.A2(n_586),
.B1(n_603),
.B2(n_588),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1225),
.B(n_630),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1386),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1357),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1346),
.B(n_585),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1251),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1252),
.A2(n_1040),
.B(n_1056),
.C(n_795),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1284),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1314),
.B(n_1059),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1208),
.B(n_587),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1246),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1208),
.B(n_587),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1360),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1363),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1328),
.B(n_631),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1376),
.B(n_633),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1245),
.B(n_1063),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1346),
.B(n_1065),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1379),
.B(n_1065),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1286),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1204),
.B(n_873),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1379),
.B(n_930),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1336),
.B(n_955),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1319),
.B(n_955),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1325),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1365),
.B(n_1256),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1247),
.A2(n_593),
.B1(n_601),
.B2(n_589),
.Y(n_1534)
);

INVx8_ASAP7_75t_L g1535 ( 
.A(n_1381),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1208),
.B(n_589),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1323),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1381),
.B(n_593),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1291),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1381),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1258),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1310),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1312),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1364),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1343),
.B(n_985),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1319),
.B(n_601),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1367),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1313),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1334),
.B(n_639),
.C(n_635),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1334),
.B(n_876),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1388),
.B(n_777),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1388),
.B(n_777),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1302),
.B(n_879),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1315),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1361),
.B(n_641),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1343),
.B(n_985),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1272),
.B(n_880),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1273),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1351),
.B(n_778),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1274),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1275),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1277),
.B(n_881),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1348),
.B(n_1015),
.Y(n_1563)
);

INVxp33_ASAP7_75t_L g1564 ( 
.A(n_1209),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1278),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1316),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1329),
.Y(n_1567)
);

BUFx8_ASAP7_75t_L g1568 ( 
.A(n_1280),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1281),
.A2(n_787),
.B1(n_788),
.B2(n_778),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1283),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1317),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1289),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1318),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1362),
.B(n_787),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1368),
.B(n_788),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1290),
.Y(n_1576)
);

AO22x1_ASAP7_75t_L g1577 ( 
.A1(n_1359),
.A2(n_588),
.B1(n_595),
.B2(n_586),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1372),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1292),
.B(n_955),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1359),
.A2(n_698),
.B1(n_712),
.B2(n_692),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1320),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1354),
.B(n_1015),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1321),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1394),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1418),
.B(n_1300),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1439),
.B(n_1293),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1409),
.A2(n_1390),
.B(n_1383),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1470),
.B(n_1324),
.Y(n_1588)
);

BUFx12f_ASAP7_75t_L g1589 ( 
.A(n_1491),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1523),
.A2(n_733),
.B1(n_738),
.B2(n_716),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1495),
.B(n_1492),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1434),
.B(n_1382),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1466),
.B(n_1384),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1445),
.A2(n_1370),
.B1(n_1371),
.B2(n_1369),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1401),
.B(n_1378),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1456),
.A2(n_968),
.B(n_938),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1421),
.B(n_1326),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1393),
.B(n_1387),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1395),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1535),
.Y(n_1600)
);

AND2x2_ASAP7_75t_SL g1601 ( 
.A(n_1522),
.B(n_1533),
.Y(n_1601)
);

NAND2x1_ASAP7_75t_L g1602 ( 
.A(n_1475),
.B(n_1359),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1509),
.A2(n_753),
.B1(n_756),
.B2(n_750),
.Y(n_1603)
);

NOR3xp33_ASAP7_75t_L g1604 ( 
.A(n_1425),
.B(n_885),
.C(n_884),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1477),
.B(n_1553),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1490),
.A2(n_796),
.B(n_802),
.C(n_794),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1423),
.B(n_1380),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1409),
.A2(n_1333),
.B(n_1332),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1488),
.B(n_1335),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1479),
.A2(n_938),
.B(n_945),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1412),
.B(n_1337),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1472),
.A2(n_938),
.B(n_945),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1419),
.A2(n_1342),
.B(n_1339),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1397),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1454),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1503),
.A2(n_1528),
.B(n_1452),
.C(n_1422),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1562),
.B(n_1359),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1424),
.B(n_791),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1430),
.A2(n_1016),
.B(n_1015),
.Y(n_1619)
);

INVx5_ASAP7_75t_L g1620 ( 
.A(n_1535),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1437),
.A2(n_1031),
.B(n_1016),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1397),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1550),
.B(n_791),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1400),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1550),
.B(n_886),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1484),
.B(n_800),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1448),
.A2(n_1031),
.B(n_1016),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1392),
.A2(n_1402),
.B(n_1411),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1438),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1487),
.B(n_887),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1544),
.B(n_800),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1502),
.B(n_812),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1546),
.B(n_812),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1512),
.B(n_595),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1506),
.A2(n_761),
.B1(n_763),
.B2(n_757),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1404),
.A2(n_1031),
.B(n_1016),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1416),
.B(n_803),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1404),
.A2(n_1031),
.B(n_1016),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1555),
.B(n_810),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1499),
.B(n_888),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1459),
.A2(n_1041),
.B(n_1035),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1512),
.B(n_603),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1403),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1406),
.B(n_813),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1541),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1460),
.B(n_643),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1476),
.A2(n_814),
.B(n_689),
.C(n_707),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1500),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1565),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1473),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1485),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1449),
.A2(n_962),
.B(n_891),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1494),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1551),
.A2(n_689),
.B(n_707),
.C(n_664),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1398),
.B(n_890),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1435),
.B(n_645),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1513),
.B(n_604),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1453),
.A2(n_1035),
.B(n_1031),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1405),
.B(n_892),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1564),
.B(n_649),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1415),
.B(n_1557),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1505),
.B(n_604),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1411),
.A2(n_1035),
.B(n_1031),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1537),
.B(n_654),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1545),
.A2(n_1041),
.B(n_1035),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1552),
.B(n_657),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1497),
.B(n_896),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1545),
.A2(n_1035),
.B(n_1044),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1556),
.A2(n_1035),
.B(n_1044),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1504),
.B(n_899),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1549),
.B(n_608),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1511),
.B(n_1520),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1521),
.B(n_903),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1547),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1471),
.B(n_904),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1455),
.B(n_906),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1518),
.B(n_663),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1397),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1493),
.B(n_608),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1478),
.B(n_907),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1432),
.A2(n_771),
.B(n_779),
.C(n_747),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1475),
.B(n_914),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1442),
.A2(n_771),
.B(n_747),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1556),
.A2(n_1044),
.B(n_1041),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1563),
.A2(n_1044),
.B(n_1041),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1558),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1410),
.B(n_666),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1426),
.B(n_669),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1535),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1538),
.A2(n_779),
.B(n_672),
.C(n_675),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1428),
.B(n_671),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1481),
.A2(n_679),
.B1(n_681),
.B2(n_678),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1542),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1560),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1446),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1431),
.B(n_682),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1543),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1548),
.Y(n_1698)
);

AND2x6_ASAP7_75t_L g1699 ( 
.A(n_1567),
.B(n_1046),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1457),
.A2(n_928),
.B(n_687),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1414),
.A2(n_690),
.B(n_693),
.C(n_686),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1582),
.A2(n_1408),
.B(n_1407),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1482),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1568),
.B(n_782),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1447),
.B(n_695),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1500),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1554),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1408),
.A2(n_1046),
.B(n_936),
.Y(n_1708)
);

INVxp33_ASAP7_75t_SL g1709 ( 
.A(n_1486),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1566),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1561),
.A2(n_783),
.B(n_784),
.C(n_782),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1570),
.B(n_696),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1524),
.A2(n_1046),
.B(n_936),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1572),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1571),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1482),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1576),
.Y(n_1717)
);

O2A1O1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1417),
.A2(n_1559),
.B(n_1575),
.C(n_1574),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1573),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1581),
.B(n_704),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1583),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1508),
.B(n_705),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1489),
.A2(n_931),
.B(n_951),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1396),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1568),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1475),
.A2(n_784),
.B1(n_793),
.B2(n_783),
.Y(n_1726)
);

AOI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1530),
.A2(n_946),
.B(n_943),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1489),
.A2(n_1496),
.B(n_1458),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1516),
.B(n_706),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1496),
.A2(n_931),
.B(n_951),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1514),
.A2(n_1436),
.B(n_1529),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1534),
.A2(n_709),
.B1(n_710),
.B2(n_708),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1569),
.B(n_793),
.Y(n_1733)
);

CKINVDCx10_ASAP7_75t_R g1734 ( 
.A(n_1420),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1515),
.B(n_713),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1525),
.A2(n_931),
.B(n_951),
.Y(n_1736)
);

O2A1O1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1461),
.A2(n_717),
.B(n_719),
.C(n_715),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1527),
.B(n_721),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1526),
.A2(n_931),
.B(n_951),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1577),
.B(n_799),
.C(n_805),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1427),
.A2(n_954),
.B(n_951),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1429),
.A2(n_954),
.B(n_946),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1580),
.A2(n_805),
.B(n_807),
.C(n_799),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1473),
.Y(n_1744)
);

INVxp33_ASAP7_75t_L g1745 ( 
.A(n_1531),
.Y(n_1745)
);

NOR2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1540),
.B(n_807),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1539),
.B(n_723),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1399),
.B(n_725),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1443),
.B(n_727),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1578),
.B(n_1464),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1467),
.A2(n_954),
.B(n_946),
.Y(n_1751)
);

AND2x2_ASAP7_75t_SL g1752 ( 
.A(n_1440),
.B(n_0),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1444),
.B(n_728),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1450),
.B(n_730),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1467),
.A2(n_954),
.B(n_946),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1451),
.B(n_731),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1465),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1480),
.B(n_1510),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1446),
.B(n_732),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_L g1760 ( 
.A(n_1446),
.B(n_808),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1517),
.A2(n_739),
.B(n_740),
.C(n_735),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1614),
.Y(n_1762)
);

INVx3_ASAP7_75t_SL g1763 ( 
.A(n_1649),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1591),
.B(n_1519),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1616),
.A2(n_1536),
.B(n_1507),
.C(n_1433),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1661),
.A2(n_1474),
.B1(n_1468),
.B2(n_1441),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1609),
.B(n_1463),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1597),
.B(n_1469),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1645),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1588),
.B(n_1579),
.Y(n_1770)
);

BUFx12f_ASAP7_75t_L g1771 ( 
.A(n_1589),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1640),
.B(n_1462),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1615),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1605),
.B(n_1598),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1639),
.A2(n_1501),
.B(n_1483),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1592),
.B(n_1498),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1646),
.B(n_1413),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1601),
.A2(n_1441),
.B1(n_1420),
.B2(n_1482),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1702),
.A2(n_1532),
.B(n_1498),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1740),
.A2(n_809),
.B1(n_808),
.B2(n_743),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_SL g1781 ( 
.A1(n_1743),
.A2(n_1532),
.B(n_1498),
.C(n_2),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1748),
.B(n_1532),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1584),
.B(n_741),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1693),
.Y(n_1784)
);

AO21x1_ASAP7_75t_L g1785 ( 
.A1(n_1595),
.A2(n_0),
.B(n_1),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1620),
.B(n_943),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1697),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1695),
.B(n_947),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1600),
.Y(n_1789)
);

AOI22x1_ASAP7_75t_L g1790 ( 
.A1(n_1608),
.A2(n_809),
.B1(n_755),
.B2(n_758),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1698),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1745),
.B(n_744),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1629),
.B(n_759),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1731),
.A2(n_954),
.B(n_947),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1618),
.B(n_762),
.Y(n_1795)
);

AOI21x1_ASAP7_75t_L g1796 ( 
.A1(n_1727),
.A2(n_947),
.B(n_928),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1630),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1731),
.A2(n_928),
.B(n_576),
.Y(n_1798)
);

OAI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1666),
.A2(n_766),
.B(n_765),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1633),
.A2(n_768),
.B1(n_776),
.B2(n_767),
.Y(n_1800)
);

BUFx8_ASAP7_75t_L g1801 ( 
.A(n_1725),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1585),
.A2(n_815),
.B1(n_3),
.B2(n_1),
.Y(n_1802)
);

OR2x6_ASAP7_75t_SL g1803 ( 
.A(n_1759),
.B(n_2),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1586),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1656),
.B(n_4),
.C(n_5),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1625),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1655),
.B(n_6),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1659),
.B(n_8),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1664),
.B(n_414),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1637),
.B(n_8),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1625),
.B(n_9),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1610),
.A2(n_928),
.B(n_571),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1672),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1626),
.B(n_9),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1611),
.B(n_10),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1709),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1587),
.A2(n_1728),
.B(n_1619),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1718),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1683),
.A2(n_419),
.B(n_418),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1593),
.Y(n_1820)
);

O2A1O1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1679),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1607),
.B(n_14),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1660),
.B(n_420),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1590),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1636),
.A2(n_573),
.B(n_422),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1677),
.B(n_17),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1706),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1603),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1729),
.A2(n_19),
.B(n_22),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1631),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1758),
.B(n_24),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1638),
.A2(n_425),
.B(n_421),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1667),
.B(n_25),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1635),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1676),
.B(n_27),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1750),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1670),
.B(n_29),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1722),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_SL g1839 ( 
.A(n_1648),
.B(n_1620),
.Y(n_1839)
);

A2O1A1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1690),
.A2(n_35),
.B(n_32),
.C(n_34),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1593),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1707),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1612),
.A2(n_427),
.B(n_426),
.Y(n_1843)
);

BUFx12f_ASAP7_75t_L g1844 ( 
.A(n_1746),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1634),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_SL g1846 ( 
.A1(n_1602),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1734),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1641),
.A2(n_572),
.B(n_430),
.Y(n_1848)
);

INVx4_ASAP7_75t_L g1849 ( 
.A(n_1600),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1596),
.A2(n_567),
.B(n_431),
.Y(n_1850)
);

INVx4_ASAP7_75t_L g1851 ( 
.A(n_1614),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1676),
.B(n_39),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1614),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1621),
.A2(n_566),
.B(n_432),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1622),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1682),
.B(n_39),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1632),
.B(n_1671),
.Y(n_1857)
);

AO32x1_ASAP7_75t_L g1858 ( 
.A1(n_1594),
.A2(n_42),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1710),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1617),
.B(n_40),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1700),
.A2(n_433),
.B(n_429),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1599),
.Y(n_1862)
);

OR2x6_ASAP7_75t_SL g1863 ( 
.A(n_1726),
.B(n_41),
.Y(n_1863)
);

NAND2x1_ASAP7_75t_L g1864 ( 
.A(n_1699),
.B(n_436),
.Y(n_1864)
);

BUFx8_ASAP7_75t_L g1865 ( 
.A(n_1622),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1682),
.B(n_42),
.Y(n_1866)
);

INVxp33_ASAP7_75t_L g1867 ( 
.A(n_1623),
.Y(n_1867)
);

INVx3_ASAP7_75t_SL g1868 ( 
.A(n_1752),
.Y(n_1868)
);

BUFx2_ASAP7_75t_SL g1869 ( 
.A(n_1689),
.Y(n_1869)
);

INVx4_ASAP7_75t_L g1870 ( 
.A(n_1622),
.Y(n_1870)
);

INVx4_ASAP7_75t_L g1871 ( 
.A(n_1678),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1673),
.B(n_44),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1700),
.A2(n_562),
.B(n_443),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1624),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1658),
.A2(n_560),
.B(n_444),
.Y(n_1875)
);

O2A1O1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1642),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1675),
.B(n_45),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1715),
.B(n_1721),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1701),
.A2(n_1652),
.B(n_1737),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1663),
.A2(n_559),
.B(n_445),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1643),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1761),
.A2(n_49),
.B(n_46),
.C(n_47),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1686),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1657),
.B(n_438),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1724),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1651),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1680),
.B(n_51),
.Y(n_1887)
);

O2A1O1Ixp5_ASAP7_75t_L g1888 ( 
.A1(n_1628),
.A2(n_1627),
.B(n_1662),
.C(n_1681),
.Y(n_1888)
);

INVx5_ASAP7_75t_L g1889 ( 
.A(n_1699),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1678),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1613),
.A2(n_450),
.B(n_447),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1719),
.B(n_1757),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1733),
.B(n_452),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1665),
.A2(n_558),
.B(n_454),
.Y(n_1894)
);

OAI21xp33_ASAP7_75t_L g1895 ( 
.A1(n_1604),
.A2(n_51),
.B(n_52),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1644),
.B(n_53),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_L g1897 ( 
.A(n_1732),
.B(n_53),
.C(n_54),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1695),
.B(n_54),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1653),
.Y(n_1899)
);

AOI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1668),
.A2(n_455),
.B(n_453),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1674),
.B(n_55),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1687),
.B(n_55),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1694),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1688),
.B(n_56),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1669),
.A2(n_458),
.B(n_456),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1691),
.B(n_56),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1696),
.B(n_1705),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1712),
.B(n_57),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1714),
.B(n_57),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1678),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_SL g1911 ( 
.A1(n_1711),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1703),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1717),
.B(n_60),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1689),
.B(n_459),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1720),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1684),
.A2(n_461),
.B(n_460),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1692),
.B(n_62),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1760),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1735),
.B(n_64),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1654),
.B(n_1647),
.C(n_1606),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1738),
.B(n_65),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_L g1922 ( 
.A1(n_1685),
.A2(n_464),
.B(n_463),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1716),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1703),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1886),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1817),
.A2(n_1794),
.A3(n_1873),
.B(n_1861),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1862),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1813),
.B(n_1716),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_L g1929 ( 
.A(n_1805),
.B(n_1704),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1767),
.A2(n_1650),
.B1(n_1744),
.B2(n_1747),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1874),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1772),
.B(n_1749),
.Y(n_1932)
);

AOI21xp33_ASAP7_75t_L g1933 ( 
.A1(n_1879),
.A2(n_1754),
.B(n_1753),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_R g1934 ( 
.A(n_1771),
.B(n_1844),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1867),
.B(n_1756),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1797),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1907),
.B(n_1703),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1798),
.A2(n_1742),
.B(n_1751),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1777),
.A2(n_1708),
.B1(n_1713),
.B2(n_1755),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1773),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1881),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_SL g1942 ( 
.A1(n_1785),
.A2(n_1730),
.B(n_1723),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1768),
.B(n_1699),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1903),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1770),
.B(n_1699),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1774),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1899),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1920),
.A2(n_1799),
.B(n_1897),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1892),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1763),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1776),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1815),
.B(n_66),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1920),
.A2(n_1741),
.B(n_1739),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1923),
.B(n_465),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1764),
.B(n_67),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1895),
.A2(n_1809),
.B(n_1829),
.C(n_1823),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1819),
.A2(n_1736),
.B(n_469),
.Y(n_1957)
);

OAI21x1_ASAP7_75t_L g1958 ( 
.A1(n_1796),
.A2(n_470),
.B(n_468),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1820),
.B(n_68),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1799),
.A2(n_69),
.B(n_70),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1779),
.A2(n_474),
.B(n_473),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1841),
.B(n_69),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1900),
.A2(n_476),
.B(n_475),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1766),
.B(n_478),
.Y(n_1964)
);

NAND2x1p5_ASAP7_75t_L g1965 ( 
.A(n_1889),
.B(n_1839),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1769),
.B(n_70),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1784),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1787),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1791),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1917),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1842),
.B(n_71),
.Y(n_1971)
);

AOI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1850),
.A2(n_481),
.B(n_480),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1859),
.B(n_72),
.Y(n_1973)
);

OAI21x1_ASAP7_75t_L g1974 ( 
.A1(n_1922),
.A2(n_1888),
.B(n_1854),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1853),
.Y(n_1975)
);

NAND3xp33_ASAP7_75t_SL g1976 ( 
.A(n_1816),
.B(n_73),
.C(n_74),
.Y(n_1976)
);

AO31x2_ASAP7_75t_L g1977 ( 
.A1(n_1818),
.A2(n_485),
.A3(n_487),
.B(n_483),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1885),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1775),
.A2(n_489),
.B(n_488),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1868),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1810),
.B(n_75),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1782),
.B(n_76),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1762),
.Y(n_1983)
);

OAI21x1_ASAP7_75t_L g1984 ( 
.A1(n_1880),
.A2(n_491),
.B(n_490),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1848),
.A2(n_495),
.B(n_493),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1875),
.A2(n_497),
.B(n_496),
.Y(n_1986)
);

AOI21x1_ASAP7_75t_L g1987 ( 
.A1(n_1843),
.A2(n_500),
.B(n_499),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1889),
.A2(n_502),
.B(n_501),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1889),
.A2(n_505),
.B(n_504),
.Y(n_1989)
);

INVxp67_ASAP7_75t_SL g1990 ( 
.A(n_1878),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1891),
.A2(n_508),
.B(n_506),
.Y(n_1991)
);

AOI21xp33_ASAP7_75t_L g1992 ( 
.A1(n_1765),
.A2(n_1895),
.B(n_1790),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1807),
.B(n_77),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1792),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1812),
.A2(n_510),
.B(n_509),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1825),
.A2(n_1832),
.B(n_1894),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1789),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1808),
.B(n_1822),
.Y(n_1998)
);

AND3x4_ASAP7_75t_L g1999 ( 
.A(n_1914),
.B(n_78),
.C(n_79),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1762),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1827),
.Y(n_2001)
);

NAND2x1p5_ASAP7_75t_L g2002 ( 
.A(n_1789),
.B(n_513),
.Y(n_2002)
);

AOI221x1_ASAP7_75t_L g2003 ( 
.A1(n_1805),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1856),
.B(n_514),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1860),
.B(n_80),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1806),
.B(n_517),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1901),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1840),
.A2(n_81),
.B(n_82),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1882),
.A2(n_83),
.B(n_84),
.Y(n_2009)
);

OAI21x1_ASAP7_75t_L g2010 ( 
.A1(n_1905),
.A2(n_1916),
.B(n_1864),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1913),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1814),
.B(n_1833),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1837),
.B(n_85),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1855),
.Y(n_2014)
);

OAI22x1_ASAP7_75t_L g2015 ( 
.A1(n_1816),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_2015)
);

INVx4_ASAP7_75t_SL g2016 ( 
.A(n_1847),
.Y(n_2016)
);

OAI21x1_ASAP7_75t_L g2017 ( 
.A1(n_1786),
.A2(n_519),
.B(n_518),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1865),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1858),
.A2(n_521),
.B(n_520),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1858),
.A2(n_1893),
.B(n_1781),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1858),
.A2(n_523),
.B(n_522),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1846),
.A2(n_528),
.B(n_525),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1831),
.B(n_1896),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1909),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1865),
.Y(n_2025)
);

AO21x2_ASAP7_75t_L g2026 ( 
.A1(n_1921),
.A2(n_87),
.B(n_88),
.Y(n_2026)
);

AO22x2_ASAP7_75t_L g2027 ( 
.A1(n_1824),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1795),
.A2(n_531),
.B(n_530),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1911),
.A2(n_538),
.B(n_535),
.Y(n_2029)
);

AOI21xp33_ASAP7_75t_L g2030 ( 
.A1(n_1821),
.A2(n_91),
.B(n_92),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1857),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1778),
.B(n_539),
.Y(n_2032)
);

OAI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_1826),
.A2(n_97),
.B1(n_93),
.B2(n_94),
.C(n_98),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1912),
.A2(n_1876),
.B(n_1845),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1912),
.A2(n_542),
.B(n_541),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1918),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1872),
.B(n_99),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1877),
.B(n_100),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1940),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1951),
.B(n_1811),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1927),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1931),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1936),
.B(n_1866),
.Y(n_2043)
);

BUFx2_ASAP7_75t_SL g2044 ( 
.A(n_1950),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1946),
.B(n_1924),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1941),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1947),
.B(n_1838),
.Y(n_2047)
);

NOR2x1_ASAP7_75t_L g2048 ( 
.A(n_1929),
.B(n_1869),
.Y(n_2048)
);

A2O1A1Ixp33_ASAP7_75t_L g2049 ( 
.A1(n_1956),
.A2(n_1838),
.B(n_1884),
.C(n_1902),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1940),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1932),
.B(n_1904),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1925),
.Y(n_2052)
);

INVxp67_ASAP7_75t_L g2053 ( 
.A(n_2001),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1975),
.B(n_1914),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1949),
.B(n_1908),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_2016),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1996),
.A2(n_1919),
.B(n_1887),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_2018),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1944),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1940),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1978),
.Y(n_2061)
);

BUFx2_ASAP7_75t_SL g2062 ( 
.A(n_2025),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1978),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1957),
.A2(n_1828),
.B(n_1834),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2014),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1976),
.A2(n_1830),
.B1(n_1915),
.B2(n_1802),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_1948),
.A2(n_1836),
.B1(n_1804),
.B2(n_1835),
.Y(n_2067)
);

OAI21xp33_ASAP7_75t_L g2068 ( 
.A1(n_1960),
.A2(n_1883),
.B(n_1906),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_2000),
.Y(n_2069)
);

NAND2x1_ASAP7_75t_L g2070 ( 
.A(n_1967),
.B(n_1788),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_2000),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2007),
.B(n_1852),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2024),
.B(n_1803),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2011),
.B(n_1863),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2023),
.B(n_1890),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1968),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_1935),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1933),
.A2(n_1898),
.B(n_1800),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1990),
.B(n_1793),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_2000),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2012),
.B(n_1937),
.Y(n_2081)
);

OR2x6_ASAP7_75t_L g2082 ( 
.A(n_1965),
.B(n_1849),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2009),
.A2(n_1801),
.B1(n_1783),
.B2(n_1780),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1997),
.B(n_1851),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1969),
.B(n_1851),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1928),
.Y(n_2086)
);

A2O1A1Ixp33_ASAP7_75t_SL g2087 ( 
.A1(n_2033),
.A2(n_1801),
.B(n_1788),
.C(n_1849),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1979),
.A2(n_1871),
.B(n_1870),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1992),
.A2(n_1871),
.B(n_1870),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_1983),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1983),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1991),
.A2(n_1910),
.B(n_1788),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_1938),
.A2(n_1910),
.B(n_1788),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1966),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1971),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_1943),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1998),
.B(n_1762),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_1954),
.B(n_543),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1994),
.B(n_100),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_1954),
.Y(n_2100)
);

OAI21xp33_ASAP7_75t_L g2101 ( 
.A1(n_2008),
.A2(n_101),
.B(n_102),
.Y(n_2101)
);

OAI22xp33_ASAP7_75t_SL g2102 ( 
.A1(n_2031),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2102)
);

O2A1O1Ixp5_ASAP7_75t_SL g2103 ( 
.A1(n_1939),
.A2(n_106),
.B(n_103),
.C(n_104),
.Y(n_2103)
);

INVx3_ASAP7_75t_SL g2104 ( 
.A(n_2016),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1959),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1973),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1945),
.B(n_556),
.Y(n_2107)
);

AND2x2_ASAP7_75t_SL g2108 ( 
.A(n_1970),
.B(n_107),
.Y(n_2108)
);

OR2x6_ASAP7_75t_L g2109 ( 
.A(n_1942),
.B(n_544),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_2034),
.Y(n_2110)
);

NAND2xp33_ASAP7_75t_L g2111 ( 
.A(n_2015),
.B(n_108),
.Y(n_2111)
);

INVx5_ASAP7_75t_L g2112 ( 
.A(n_2004),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_1982),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2029),
.A2(n_550),
.B(n_549),
.Y(n_2114)
);

INVx3_ASAP7_75t_SL g2115 ( 
.A(n_2032),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1962),
.Y(n_2116)
);

INVx8_ASAP7_75t_L g2117 ( 
.A(n_2098),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2041),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2042),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_2060),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_SL g2121 ( 
.A1(n_2108),
.A2(n_2027),
.B1(n_2020),
.B2(n_1980),
.Y(n_2121)
);

BUFx8_ASAP7_75t_L g2122 ( 
.A(n_2098),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2101),
.A2(n_2027),
.B1(n_1999),
.B2(n_2030),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_SL g2124 ( 
.A1(n_2111),
.A2(n_2036),
.B1(n_2026),
.B2(n_2019),
.Y(n_2124)
);

AOI22xp33_ASAP7_75t_L g2125 ( 
.A1(n_2101),
.A2(n_1964),
.B1(n_2005),
.B2(n_1952),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2046),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_2044),
.Y(n_2127)
);

BUFx12f_ASAP7_75t_L g2128 ( 
.A(n_2107),
.Y(n_2128)
);

BUFx2_ASAP7_75t_L g2129 ( 
.A(n_2065),
.Y(n_2129)
);

CKINVDCx6p67_ASAP7_75t_R g2130 ( 
.A(n_2104),
.Y(n_2130)
);

INVx6_ASAP7_75t_SL g2131 ( 
.A(n_2082),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2083),
.A2(n_1930),
.B1(n_2022),
.B2(n_1981),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2061),
.Y(n_2133)
);

INVx6_ASAP7_75t_L g2134 ( 
.A(n_2112),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_2068),
.A2(n_1993),
.B1(n_2037),
.B2(n_2013),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2063),
.Y(n_2136)
);

CKINVDCx20_ASAP7_75t_R g2137 ( 
.A(n_2058),
.Y(n_2137)
);

INVx3_ASAP7_75t_SL g2138 ( 
.A(n_2056),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2068),
.A2(n_2038),
.B1(n_1955),
.B2(n_2021),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2096),
.B(n_1926),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2064),
.A2(n_2028),
.B1(n_2006),
.B2(n_1995),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2076),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_2066),
.A2(n_1961),
.B1(n_1953),
.B2(n_1988),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_SL g2144 ( 
.A1(n_2102),
.A2(n_2003),
.B1(n_2002),
.B2(n_1984),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2052),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2066),
.A2(n_1989),
.B1(n_1985),
.B2(n_1986),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_2062),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2059),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2053),
.B(n_1926),
.Y(n_2149)
);

INVx6_ASAP7_75t_L g2150 ( 
.A(n_2112),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2067),
.A2(n_2102),
.B1(n_2078),
.B2(n_2099),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_2090),
.Y(n_2152)
);

AOI21xp33_ASAP7_75t_L g2153 ( 
.A1(n_2087),
.A2(n_2035),
.B(n_1963),
.Y(n_2153)
);

INVx5_ASAP7_75t_L g2154 ( 
.A(n_2109),
.Y(n_2154)
);

AOI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_2049),
.A2(n_2010),
.B1(n_2017),
.B2(n_1974),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_2100),
.Y(n_2156)
);

OAI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2047),
.A2(n_1987),
.B1(n_1972),
.B2(n_1977),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2086),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2045),
.Y(n_2159)
);

CKINVDCx20_ASAP7_75t_R g2160 ( 
.A(n_2075),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_2084),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2110),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_2084),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_2140),
.B(n_2047),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_2057),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2152),
.B(n_2129),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2159),
.B(n_2073),
.Y(n_2167)
);

O2A1O1Ixp5_ASAP7_75t_L g2168 ( 
.A1(n_2132),
.A2(n_2157),
.B(n_2153),
.C(n_2114),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2161),
.B(n_2163),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2137),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2161),
.B(n_2105),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2163),
.B(n_2043),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2133),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2149),
.B(n_2074),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_2134),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2162),
.B(n_2074),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2136),
.Y(n_2177)
);

AOI21x1_ASAP7_75t_SL g2178 ( 
.A1(n_2130),
.A2(n_2055),
.B(n_2079),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2123),
.A2(n_2077),
.B1(n_2112),
.B2(n_2079),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_2154),
.B(n_2082),
.Y(n_2180)
);

AOI21x1_ASAP7_75t_SL g2181 ( 
.A1(n_2121),
.A2(n_2055),
.B(n_2072),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2148),
.B(n_2081),
.Y(n_2182)
);

O2A1O1Ixp33_ASAP7_75t_L g2183 ( 
.A1(n_2123),
.A2(n_2072),
.B(n_2051),
.C(n_2094),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2154),
.B(n_2082),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2121),
.A2(n_2048),
.B1(n_2115),
.B2(n_2113),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_2154),
.B(n_2085),
.Y(n_2186)
);

A2O1A1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_2151),
.A2(n_2093),
.B(n_2088),
.C(n_2092),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2118),
.B(n_2119),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_2145),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_2138),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_R g2191 ( 
.A(n_2190),
.B(n_2138),
.Y(n_2191)
);

CKINVDCx16_ASAP7_75t_R g2192 ( 
.A(n_2166),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2164),
.B(n_2126),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2164),
.B(n_2142),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2174),
.B(n_2116),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2173),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2187),
.A2(n_2141),
.B(n_2143),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2165),
.Y(n_2198)
);

NAND2xp33_ASAP7_75t_R g2199 ( 
.A(n_2170),
.B(n_2109),
.Y(n_2199)
);

HB1xp67_ASAP7_75t_L g2200 ( 
.A(n_2165),
.Y(n_2200)
);

INVx5_ASAP7_75t_SL g2201 ( 
.A(n_2180),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2198),
.B(n_2175),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2200),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_2201),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2196),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2194),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2192),
.B(n_2175),
.Y(n_2207)
);

AO21x2_ASAP7_75t_L g2208 ( 
.A1(n_2197),
.A2(n_2185),
.B(n_2179),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_2201),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2202),
.B(n_2174),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2202),
.B(n_2193),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2203),
.B(n_2206),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_2207),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2203),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_2207),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_2202),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2205),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2205),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_2208),
.A2(n_2179),
.B1(n_2151),
.B2(n_2185),
.Y(n_2219)
);

AOI221x1_ASAP7_75t_L g2220 ( 
.A1(n_2214),
.A2(n_2204),
.B1(n_2209),
.B2(n_2207),
.C(n_2206),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_2216),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_L g2222 ( 
.A(n_2219),
.B(n_2168),
.C(n_2135),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2213),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2219),
.A2(n_2208),
.B1(n_2204),
.B2(n_2209),
.Y(n_2224)
);

OAI211xp5_ASAP7_75t_L g2225 ( 
.A1(n_2215),
.A2(n_2135),
.B(n_2183),
.C(n_2144),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2212),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2215),
.B(n_2204),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_SL g2228 ( 
.A1(n_2210),
.A2(n_2208),
.B1(n_2191),
.B2(n_2204),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2211),
.B(n_2204),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2212),
.A2(n_2208),
.B1(n_2209),
.B2(n_2154),
.Y(n_2230)
);

NAND3xp33_ASAP7_75t_L g2231 ( 
.A(n_2217),
.B(n_2168),
.C(n_2183),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2221),
.B(n_2218),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_SL g2233 ( 
.A(n_2227),
.B(n_2209),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2226),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2223),
.B(n_2209),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2229),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2228),
.B(n_2166),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2220),
.Y(n_2238)
);

NAND2x1_ASAP7_75t_L g2239 ( 
.A(n_2224),
.B(n_2205),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_2231),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2236),
.B(n_2222),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2238),
.B(n_2228),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2240),
.B(n_2225),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2237),
.B(n_2230),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2244),
.B(n_2234),
.Y(n_2245)
);

OAI21xp33_ASAP7_75t_L g2246 ( 
.A1(n_2243),
.A2(n_2233),
.B(n_2235),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_2241),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2242),
.Y(n_2248)
);

OAI211xp5_ASAP7_75t_L g2249 ( 
.A1(n_2246),
.A2(n_2239),
.B(n_2232),
.C(n_2225),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_2245),
.Y(n_2250)
);

NOR3xp33_ASAP7_75t_L g2251 ( 
.A(n_2247),
.B(n_2232),
.C(n_1934),
.Y(n_2251)
);

AOI211xp5_ASAP7_75t_L g2252 ( 
.A1(n_2248),
.A2(n_2147),
.B(n_2127),
.C(n_2180),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2246),
.B(n_2160),
.Y(n_2253)
);

INVxp67_ASAP7_75t_SL g2254 ( 
.A(n_2247),
.Y(n_2254)
);

CKINVDCx14_ASAP7_75t_R g2255 ( 
.A(n_2253),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2254),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_2250),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2251),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2249),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2252),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2254),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2254),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2254),
.B(n_2167),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2250),
.Y(n_2264)
);

A2O1A1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_2259),
.A2(n_2175),
.B(n_2176),
.C(n_2180),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2264),
.B(n_2176),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2263),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2256),
.B(n_2171),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2257),
.B(n_2167),
.Y(n_2269)
);

AOI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2255),
.A2(n_2199),
.B1(n_2039),
.B2(n_2050),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2261),
.B(n_2180),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2262),
.B(n_2116),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2255),
.B(n_2171),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2260),
.Y(n_2274)
);

A2O1A1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2260),
.A2(n_2184),
.B(n_2125),
.C(n_2143),
.Y(n_2275)
);

AO21x1_ASAP7_75t_L g2276 ( 
.A1(n_2258),
.A2(n_2195),
.B(n_2184),
.Y(n_2276)
);

NAND3x1_ASAP7_75t_L g2277 ( 
.A(n_2259),
.B(n_2089),
.C(n_2097),
.Y(n_2277)
);

OAI221xp5_ASAP7_75t_SL g2278 ( 
.A1(n_2265),
.A2(n_2274),
.B1(n_2273),
.B2(n_2266),
.C(n_2268),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2269),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2270),
.A2(n_2184),
.B1(n_2116),
.B2(n_2156),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2267),
.Y(n_2281)
);

OAI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2275),
.A2(n_2125),
.B1(n_2124),
.B2(n_2144),
.C(n_2139),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2271),
.B(n_2172),
.Y(n_2283)
);

AOI222xp33_ASAP7_75t_L g2284 ( 
.A1(n_2272),
.A2(n_2276),
.B1(n_2277),
.B2(n_2139),
.C1(n_2157),
.C2(n_2181),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2274),
.A2(n_2184),
.B1(n_2128),
.B2(n_2150),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2269),
.B(n_2172),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2269),
.B(n_2169),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2269),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2269),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_2267),
.B(n_2120),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2267),
.B(n_2095),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2269),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2279),
.B(n_2169),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2288),
.B(n_2186),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2289),
.B(n_2292),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2281),
.B(n_109),
.Y(n_2296)
);

INVxp67_ASAP7_75t_L g2297 ( 
.A(n_2290),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2291),
.Y(n_2298)
);

OAI221xp5_ASAP7_75t_L g2299 ( 
.A1(n_2285),
.A2(n_2124),
.B1(n_2150),
.B2(n_2134),
.C(n_2109),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2283),
.Y(n_2300)
);

CKINVDCx14_ASAP7_75t_R g2301 ( 
.A(n_2278),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2286),
.B(n_2182),
.Y(n_2302)
);

INVx1_ASAP7_75t_SL g2303 ( 
.A(n_2287),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2280),
.B(n_2186),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2284),
.B(n_2186),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2282),
.B(n_2186),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2305),
.B(n_2106),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_2305),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2293),
.Y(n_2309)
);

NAND3xp33_ASAP7_75t_L g2310 ( 
.A(n_2301),
.B(n_2103),
.C(n_109),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2294),
.Y(n_2311)
);

NAND3xp33_ASAP7_75t_L g2312 ( 
.A(n_2295),
.B(n_110),
.C(n_112),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2303),
.B(n_2182),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2296),
.Y(n_2314)
);

NAND3xp33_ASAP7_75t_SL g2315 ( 
.A(n_2303),
.B(n_110),
.C(n_112),
.Y(n_2315)
);

NOR3xp33_ASAP7_75t_L g2316 ( 
.A(n_2297),
.B(n_2107),
.C(n_2097),
.Y(n_2316)
);

INVx1_ASAP7_75t_SL g2317 ( 
.A(n_2298),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2306),
.B(n_2091),
.Y(n_2318)
);

NOR3x1_ASAP7_75t_L g2319 ( 
.A(n_2300),
.B(n_113),
.C(n_114),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2302),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2304),
.B(n_2299),
.Y(n_2321)
);

NAND4xp25_ASAP7_75t_L g2322 ( 
.A(n_2303),
.B(n_2146),
.C(n_115),
.D(n_113),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2293),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2303),
.B(n_114),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2305),
.B(n_2040),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2293),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2293),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2293),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2308),
.B(n_2188),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2317),
.B(n_116),
.C(n_117),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_L g2331 ( 
.A(n_2321),
.B(n_2146),
.C(n_120),
.D(n_118),
.Y(n_2331)
);

INVxp67_ASAP7_75t_L g2332 ( 
.A(n_2324),
.Y(n_2332)
);

OAI21xp33_ASAP7_75t_SL g2333 ( 
.A1(n_2325),
.A2(n_2181),
.B(n_2188),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2311),
.Y(n_2334)
);

OAI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2312),
.A2(n_2131),
.B1(n_2150),
.B2(n_2134),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2309),
.B(n_2189),
.Y(n_2336)
);

NOR3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2315),
.B(n_118),
.C(n_119),
.Y(n_2337)
);

NAND2xp33_ASAP7_75t_SL g2338 ( 
.A(n_2307),
.B(n_2070),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2323),
.B(n_119),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2326),
.B(n_121),
.Y(n_2340)
);

NOR4xp25_ASAP7_75t_L g2341 ( 
.A(n_2327),
.B(n_123),
.C(n_121),
.D(n_122),
.Y(n_2341)
);

INVxp67_ASAP7_75t_L g2342 ( 
.A(n_2328),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2319),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2313),
.Y(n_2344)
);

OAI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2322),
.A2(n_2131),
.B1(n_2117),
.B2(n_2173),
.Y(n_2345)
);

NOR2x1_ASAP7_75t_L g2346 ( 
.A(n_2314),
.B(n_122),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2320),
.Y(n_2347)
);

AOI221xp5_ASAP7_75t_L g2348 ( 
.A1(n_2318),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2322),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2316),
.B(n_124),
.Y(n_2350)
);

NOR3xp33_ASAP7_75t_L g2351 ( 
.A(n_2310),
.B(n_127),
.C(n_128),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2308),
.B(n_127),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2308),
.B(n_128),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2308),
.B(n_2122),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2308),
.B(n_129),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_L g2356 ( 
.A1(n_2308),
.A2(n_131),
.B(n_129),
.C(n_130),
.Y(n_2356)
);

NAND4xp25_ASAP7_75t_L g2357 ( 
.A(n_2321),
.B(n_133),
.C(n_130),
.D(n_131),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2308),
.A2(n_2122),
.B1(n_2071),
.B2(n_2080),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2308),
.B(n_133),
.Y(n_2359)
);

NOR3x1_ASAP7_75t_L g2360 ( 
.A(n_2308),
.B(n_134),
.C(n_135),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_2308),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_L g2362 ( 
.A(n_2308),
.B(n_134),
.C(n_135),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2308),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2308),
.B(n_136),
.Y(n_2364)
);

NOR2xp67_ASAP7_75t_SL g2365 ( 
.A(n_2308),
.B(n_137),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2361),
.A2(n_137),
.B(n_138),
.Y(n_2366)
);

NAND3xp33_ASAP7_75t_SL g2367 ( 
.A(n_2362),
.B(n_2356),
.C(n_2363),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2365),
.B(n_138),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2354),
.B(n_2091),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2334),
.A2(n_2071),
.B1(n_2080),
.B2(n_2069),
.Y(n_2370)
);

NOR3xp33_ASAP7_75t_L g2371 ( 
.A(n_2357),
.B(n_139),
.C(n_140),
.Y(n_2371)
);

OAI221xp5_ASAP7_75t_L g2372 ( 
.A1(n_2358),
.A2(n_2155),
.B1(n_141),
.B2(n_139),
.C(n_140),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2352),
.B(n_141),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_L g2374 ( 
.A(n_2342),
.B(n_142),
.C(n_144),
.Y(n_2374)
);

INVxp33_ASAP7_75t_L g2375 ( 
.A(n_2353),
.Y(n_2375)
);

NAND4xp25_ASAP7_75t_L g2376 ( 
.A(n_2331),
.B(n_145),
.C(n_142),
.D(n_144),
.Y(n_2376)
);

NOR2x1_ASAP7_75t_L g2377 ( 
.A(n_2346),
.B(n_146),
.Y(n_2377)
);

NAND4xp25_ASAP7_75t_SL g2378 ( 
.A(n_2351),
.B(n_2178),
.C(n_149),
.D(n_147),
.Y(n_2378)
);

NAND5xp2_ASAP7_75t_L g2379 ( 
.A(n_2343),
.B(n_149),
.C(n_147),
.D(n_148),
.E(n_150),
.Y(n_2379)
);

O2A1O1Ixp5_ASAP7_75t_SL g2380 ( 
.A1(n_2347),
.A2(n_151),
.B(n_148),
.C(n_150),
.Y(n_2380)
);

NAND4xp75_ASAP7_75t_L g2381 ( 
.A(n_2360),
.B(n_155),
.C(n_153),
.D(n_154),
.Y(n_2381)
);

AOI211xp5_ASAP7_75t_L g2382 ( 
.A1(n_2341),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_2382)
);

AOI211xp5_ASAP7_75t_SL g2383 ( 
.A1(n_2355),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_2383)
);

AOI211xp5_ASAP7_75t_L g2384 ( 
.A1(n_2359),
.A2(n_159),
.B(n_156),
.C(n_158),
.Y(n_2384)
);

NOR4xp25_ASAP7_75t_SL g2385 ( 
.A(n_2349),
.B(n_161),
.C(n_159),
.D(n_160),
.Y(n_2385)
);

NAND5xp2_ASAP7_75t_L g2386 ( 
.A(n_2344),
.B(n_165),
.C(n_162),
.D(n_164),
.E(n_166),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2364),
.B(n_162),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_SL g2388 ( 
.A(n_2337),
.B(n_2091),
.Y(n_2388)
);

NOR2x1_ASAP7_75t_L g2389 ( 
.A(n_2339),
.B(n_166),
.Y(n_2389)
);

AO21x1_ASAP7_75t_L g2390 ( 
.A1(n_2340),
.A2(n_167),
.B(n_169),
.Y(n_2390)
);

NAND3xp33_ASAP7_75t_L g2391 ( 
.A(n_2348),
.B(n_167),
.C(n_169),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2329),
.B(n_170),
.Y(n_2392)
);

NOR3xp33_ASAP7_75t_L g2393 ( 
.A(n_2347),
.B(n_170),
.C(n_171),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2330),
.B(n_171),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2336),
.A2(n_2069),
.B1(n_2177),
.B2(n_2173),
.Y(n_2395)
);

OA211x2_ASAP7_75t_L g2396 ( 
.A1(n_2350),
.A2(n_2332),
.B(n_2345),
.C(n_2338),
.Y(n_2396)
);

NAND4xp75_ASAP7_75t_L g2397 ( 
.A(n_2333),
.B(n_2335),
.C(n_175),
.D(n_173),
.Y(n_2397)
);

AOI221xp5_ASAP7_75t_L g2398 ( 
.A1(n_2361),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.C(n_177),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2361),
.B(n_2177),
.Y(n_2399)
);

NOR3xp33_ASAP7_75t_L g2400 ( 
.A(n_2363),
.B(n_174),
.C(n_177),
.Y(n_2400)
);

NOR3xp33_ASAP7_75t_L g2401 ( 
.A(n_2363),
.B(n_178),
.C(n_179),
.Y(n_2401)
);

OAI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2391),
.A2(n_1958),
.B(n_2054),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2379),
.B(n_179),
.Y(n_2403)
);

OAI211xp5_ASAP7_75t_L g2404 ( 
.A1(n_2382),
.A2(n_183),
.B(n_180),
.C(n_182),
.Y(n_2404)
);

NAND3xp33_ASAP7_75t_L g2405 ( 
.A(n_2377),
.B(n_180),
.C(n_182),
.Y(n_2405)
);

NAND4xp25_ASAP7_75t_L g2406 ( 
.A(n_2396),
.B(n_185),
.C(n_183),
.D(n_184),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2390),
.Y(n_2407)
);

AOI211xp5_ASAP7_75t_L g2408 ( 
.A1(n_2376),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_2387),
.B(n_187),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2386),
.B(n_188),
.Y(n_2410)
);

NOR3x2_ASAP7_75t_L g2411 ( 
.A(n_2381),
.B(n_188),
.C(n_189),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2368),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_L g2413 ( 
.A(n_2383),
.B(n_2371),
.C(n_2366),
.Y(n_2413)
);

XNOR2xp5_ASAP7_75t_L g2414 ( 
.A(n_2384),
.B(n_189),
.Y(n_2414)
);

NAND4xp25_ASAP7_75t_L g2415 ( 
.A(n_2367),
.B(n_192),
.C(n_190),
.D(n_191),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_SL g2416 ( 
.A(n_2385),
.B(n_190),
.C(n_191),
.Y(n_2416)
);

OAI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_2370),
.A2(n_2177),
.B1(n_2117),
.B2(n_2178),
.Y(n_2417)
);

OAI21xp5_ASAP7_75t_SL g2418 ( 
.A1(n_2375),
.A2(n_192),
.B(n_194),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2389),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2373),
.Y(n_2420)
);

NAND4xp25_ASAP7_75t_L g2421 ( 
.A(n_2388),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_2421)
);

NAND4xp25_ASAP7_75t_L g2422 ( 
.A(n_2369),
.B(n_198),
.C(n_195),
.D(n_197),
.Y(n_2422)
);

AND4x1_ASAP7_75t_L g2423 ( 
.A(n_2392),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2393),
.B(n_2400),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2401),
.B(n_199),
.Y(n_2425)
);

NAND3x1_ASAP7_75t_L g2426 ( 
.A(n_2394),
.B(n_200),
.C(n_201),
.Y(n_2426)
);

NOR3xp33_ASAP7_75t_L g2427 ( 
.A(n_2397),
.B(n_201),
.C(n_202),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2398),
.A2(n_202),
.B(n_203),
.Y(n_2428)
);

OAI211xp5_ASAP7_75t_SL g2429 ( 
.A1(n_2372),
.A2(n_2374),
.B(n_2399),
.C(n_2395),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_2378),
.B(n_204),
.C(n_205),
.Y(n_2430)
);

NAND3xp33_ASAP7_75t_SL g2431 ( 
.A(n_2380),
.B(n_205),
.C(n_206),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2383),
.B(n_206),
.Y(n_2432)
);

NAND4xp25_ASAP7_75t_L g2433 ( 
.A(n_2396),
.B(n_210),
.C(n_208),
.D(n_209),
.Y(n_2433)
);

OAI211xp5_ASAP7_75t_SL g2434 ( 
.A1(n_2377),
.A2(n_211),
.B(n_208),
.C(n_209),
.Y(n_2434)
);

OAI211xp5_ASAP7_75t_SL g2435 ( 
.A1(n_2377),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_2435)
);

OAI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2382),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2436)
);

NOR2xp67_ASAP7_75t_L g2437 ( 
.A(n_2379),
.B(n_214),
.Y(n_2437)
);

NAND4xp25_ASAP7_75t_L g2438 ( 
.A(n_2396),
.B(n_217),
.C(n_215),
.D(n_216),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2370),
.A2(n_2117),
.B1(n_2085),
.B2(n_220),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2377),
.Y(n_2440)
);

NOR3xp33_ASAP7_75t_L g2441 ( 
.A(n_2367),
.B(n_218),
.C(n_219),
.Y(n_2441)
);

INVxp67_ASAP7_75t_L g2442 ( 
.A(n_2379),
.Y(n_2442)
);

OAI221xp5_ASAP7_75t_L g2443 ( 
.A1(n_2382),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.C(n_222),
.Y(n_2443)
);

OR3x1_ASAP7_75t_L g2444 ( 
.A(n_2367),
.B(n_221),
.C(n_222),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_SL g2445 ( 
.A(n_2385),
.B(n_223),
.C(n_224),
.Y(n_2445)
);

OAI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2382),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2388),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.C(n_228),
.Y(n_2447)
);

NAND3xp33_ASAP7_75t_SL g2448 ( 
.A(n_2385),
.B(n_227),
.C(n_228),
.Y(n_2448)
);

NOR3xp33_ASAP7_75t_L g2449 ( 
.A(n_2367),
.B(n_229),
.C(n_230),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2388),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.C(n_233),
.Y(n_2450)
);

OAI211xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2377),
.A2(n_234),
.B(n_231),
.C(n_233),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_2377),
.Y(n_2452)
);

NOR2xp67_ASAP7_75t_L g2453 ( 
.A(n_2379),
.B(n_234),
.Y(n_2453)
);

AOI211x1_ASAP7_75t_L g2454 ( 
.A1(n_2369),
.A2(n_238),
.B(n_235),
.C(n_237),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2383),
.B(n_235),
.Y(n_2455)
);

AOI211xp5_ASAP7_75t_L g2456 ( 
.A1(n_2416),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_2409),
.B(n_239),
.Y(n_2457)
);

HB1xp67_ASAP7_75t_L g2458 ( 
.A(n_2409),
.Y(n_2458)
);

NOR4xp25_ASAP7_75t_SL g2459 ( 
.A(n_2407),
.B(n_242),
.C(n_240),
.D(n_241),
.Y(n_2459)
);

OAI211xp5_ASAP7_75t_L g2460 ( 
.A1(n_2406),
.A2(n_243),
.B(n_240),
.C(n_242),
.Y(n_2460)
);

XOR2x2_ASAP7_75t_L g2461 ( 
.A(n_2437),
.B(n_244),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2427),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2462)
);

HB1xp67_ASAP7_75t_L g2463 ( 
.A(n_2423),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2411),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2445),
.B(n_245),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2432),
.Y(n_2466)
);

INVxp67_ASAP7_75t_L g2467 ( 
.A(n_2403),
.Y(n_2467)
);

INVx1_ASAP7_75t_SL g2468 ( 
.A(n_2444),
.Y(n_2468)
);

INVx4_ASAP7_75t_SL g2469 ( 
.A(n_2452),
.Y(n_2469)
);

NOR2x1_ASAP7_75t_L g2470 ( 
.A(n_2433),
.B(n_247),
.Y(n_2470)
);

OAI22xp33_ASAP7_75t_L g2471 ( 
.A1(n_2438),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2453),
.B(n_249),
.Y(n_2472)
);

INVx1_ASAP7_75t_SL g2473 ( 
.A(n_2455),
.Y(n_2473)
);

OAI211xp5_ASAP7_75t_SL g2474 ( 
.A1(n_2442),
.A2(n_2424),
.B(n_2440),
.C(n_2419),
.Y(n_2474)
);

NOR2x1_ASAP7_75t_L g2475 ( 
.A(n_2448),
.B(n_2405),
.Y(n_2475)
);

INVxp33_ASAP7_75t_L g2476 ( 
.A(n_2410),
.Y(n_2476)
);

BUFx12f_ASAP7_75t_L g2477 ( 
.A(n_2413),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2426),
.Y(n_2478)
);

NOR4xp25_ASAP7_75t_L g2479 ( 
.A(n_2431),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2441),
.B(n_2449),
.Y(n_2480)
);

CKINVDCx16_ASAP7_75t_R g2481 ( 
.A(n_2414),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2430),
.B(n_251),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2415),
.B(n_252),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_R g2484 ( 
.A(n_2425),
.B(n_253),
.Y(n_2484)
);

NOR3xp33_ASAP7_75t_SL g2485 ( 
.A(n_2404),
.B(n_253),
.C(n_254),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2454),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2434),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2443),
.A2(n_254),
.B(n_255),
.Y(n_2488)
);

INVxp67_ASAP7_75t_L g2489 ( 
.A(n_2421),
.Y(n_2489)
);

AND3x1_ASAP7_75t_L g2490 ( 
.A(n_2408),
.B(n_255),
.C(n_256),
.Y(n_2490)
);

NAND2xp33_ASAP7_75t_R g2491 ( 
.A(n_2412),
.B(n_256),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2447),
.B(n_257),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2420),
.B(n_257),
.Y(n_2493)
);

NAND4xp25_ASAP7_75t_L g2494 ( 
.A(n_2428),
.B(n_259),
.C(n_260),
.D(n_261),
.Y(n_2494)
);

OAI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2436),
.A2(n_259),
.B(n_260),
.Y(n_2495)
);

XNOR2xp5_ASAP7_75t_L g2496 ( 
.A(n_2422),
.B(n_262),
.Y(n_2496)
);

AOI22xp5_ASAP7_75t_L g2497 ( 
.A1(n_2435),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2418),
.B(n_263),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2450),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_2499)
);

INVx1_ASAP7_75t_SL g2500 ( 
.A(n_2439),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2446),
.B(n_267),
.Y(n_2501)
);

HB1xp67_ASAP7_75t_L g2502 ( 
.A(n_2402),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2451),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2429),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2417),
.B(n_269),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2403),
.B(n_270),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2406),
.B(n_270),
.Y(n_2507)
);

OAI221xp5_ASAP7_75t_L g2508 ( 
.A1(n_2406),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.C(n_274),
.Y(n_2508)
);

AOI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2403),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2493),
.Y(n_2510)
);

NOR2x1_ASAP7_75t_L g2511 ( 
.A(n_2457),
.B(n_2478),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2469),
.Y(n_2512)
);

AOI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2483),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_2513)
);

AOI22x1_ASAP7_75t_L g2514 ( 
.A1(n_2458),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2461),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2469),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2479),
.B(n_278),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2506),
.B(n_279),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2472),
.Y(n_2519)
);

NOR2x1_ASAP7_75t_L g2520 ( 
.A(n_2475),
.B(n_279),
.Y(n_2520)
);

NAND4xp75_ASAP7_75t_L g2521 ( 
.A(n_2470),
.B(n_280),
.C(n_281),
.D(n_282),
.Y(n_2521)
);

XNOR2xp5_ASAP7_75t_L g2522 ( 
.A(n_2496),
.B(n_2490),
.Y(n_2522)
);

AOI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2468),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_2494),
.B(n_283),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2507),
.B(n_284),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_L g2526 ( 
.A(n_2464),
.B(n_284),
.Y(n_2526)
);

XNOR2xp5_ASAP7_75t_L g2527 ( 
.A(n_2476),
.B(n_2509),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2482),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2501),
.Y(n_2529)
);

NOR2x1_ASAP7_75t_L g2530 ( 
.A(n_2474),
.B(n_285),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2463),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2485),
.B(n_285),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2471),
.B(n_286),
.Y(n_2533)
);

NAND4xp75_ASAP7_75t_L g2534 ( 
.A(n_2504),
.B(n_2466),
.C(n_2498),
.D(n_2495),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2497),
.Y(n_2535)
);

INVx2_ASAP7_75t_SL g2536 ( 
.A(n_2465),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2487),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2486),
.B(n_286),
.Y(n_2538)
);

NOR2x1_ASAP7_75t_L g2539 ( 
.A(n_2460),
.B(n_287),
.Y(n_2539)
);

NOR2x1_ASAP7_75t_L g2540 ( 
.A(n_2503),
.B(n_287),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2508),
.Y(n_2541)
);

NOR2x1_ASAP7_75t_L g2542 ( 
.A(n_2480),
.B(n_288),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2456),
.B(n_288),
.Y(n_2543)
);

AND2x4_ASAP7_75t_L g2544 ( 
.A(n_2489),
.B(n_290),
.Y(n_2544)
);

NOR2xp67_ASAP7_75t_L g2545 ( 
.A(n_2467),
.B(n_290),
.Y(n_2545)
);

NOR2x1_ASAP7_75t_L g2546 ( 
.A(n_2480),
.B(n_291),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2473),
.Y(n_2547)
);

AO22x2_ASAP7_75t_L g2548 ( 
.A1(n_2500),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2505),
.Y(n_2549)
);

NAND4xp75_ASAP7_75t_L g2550 ( 
.A(n_2488),
.B(n_292),
.C(n_294),
.D(n_295),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2477),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2499),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2491),
.Y(n_2553)
);

OAI211xp5_ASAP7_75t_L g2554 ( 
.A1(n_2462),
.A2(n_296),
.B(n_297),
.C(n_298),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_L g2555 ( 
.A1(n_2481),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_2555)
);

AND3x2_ASAP7_75t_L g2556 ( 
.A(n_2553),
.B(n_2502),
.C(n_2459),
.Y(n_2556)
);

NOR3xp33_ASAP7_75t_SL g2557 ( 
.A(n_2512),
.B(n_2492),
.C(n_2484),
.Y(n_2557)
);

NOR2x1p5_ASAP7_75t_L g2558 ( 
.A(n_2521),
.B(n_299),
.Y(n_2558)
);

NAND4xp25_ASAP7_75t_SL g2559 ( 
.A(n_2554),
.B(n_300),
.C(n_301),
.D(n_302),
.Y(n_2559)
);

AND5x1_ASAP7_75t_L g2560 ( 
.A(n_2513),
.B(n_301),
.C(n_303),
.D(n_304),
.E(n_305),
.Y(n_2560)
);

AND2x2_ASAP7_75t_SL g2561 ( 
.A(n_2538),
.B(n_303),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2545),
.B(n_306),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2542),
.Y(n_2563)
);

OAI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2516),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2520),
.B(n_308),
.Y(n_2565)
);

NOR4xp25_ASAP7_75t_L g2566 ( 
.A(n_2531),
.B(n_309),
.C(n_310),
.D(n_311),
.Y(n_2566)
);

NAND5xp2_ASAP7_75t_L g2567 ( 
.A(n_2541),
.B(n_310),
.C(n_312),
.D(n_313),
.E(n_314),
.Y(n_2567)
);

NAND5xp2_ASAP7_75t_L g2568 ( 
.A(n_2535),
.B(n_313),
.C(n_314),
.D(n_315),
.E(n_316),
.Y(n_2568)
);

OAI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2524),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_2569)
);

BUFx2_ASAP7_75t_L g2570 ( 
.A(n_2548),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2532),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_2571)
);

NAND5xp2_ASAP7_75t_L g2572 ( 
.A(n_2552),
.B(n_318),
.C(n_319),
.D(n_320),
.E(n_321),
.Y(n_2572)
);

NAND4xp25_ASAP7_75t_L g2573 ( 
.A(n_2530),
.B(n_320),
.C(n_321),
.D(n_322),
.Y(n_2573)
);

NOR3xp33_ASAP7_75t_SL g2574 ( 
.A(n_2534),
.B(n_322),
.C(n_323),
.Y(n_2574)
);

NOR3xp33_ASAP7_75t_SL g2575 ( 
.A(n_2533),
.B(n_324),
.C(n_325),
.Y(n_2575)
);

AND4x1_ASAP7_75t_L g2576 ( 
.A(n_2511),
.B(n_324),
.C(n_326),
.D(n_327),
.Y(n_2576)
);

O2A1O1Ixp33_ASAP7_75t_L g2577 ( 
.A1(n_2518),
.A2(n_326),
.B(n_327),
.C(n_328),
.Y(n_2577)
);

OAI22x1_ASAP7_75t_L g2578 ( 
.A1(n_2514),
.A2(n_328),
.B1(n_329),
.B2(n_331),
.Y(n_2578)
);

NAND4xp75_ASAP7_75t_L g2579 ( 
.A(n_2526),
.B(n_329),
.C(n_331),
.D(n_332),
.Y(n_2579)
);

NOR4xp25_ASAP7_75t_L g2580 ( 
.A(n_2525),
.B(n_333),
.C(n_334),
.D(n_335),
.Y(n_2580)
);

NAND5xp2_ASAP7_75t_L g2581 ( 
.A(n_2528),
.B(n_334),
.C(n_335),
.D(n_336),
.E(n_337),
.Y(n_2581)
);

NOR3xp33_ASAP7_75t_L g2582 ( 
.A(n_2537),
.B(n_338),
.C(n_339),
.Y(n_2582)
);

NAND4xp25_ASAP7_75t_L g2583 ( 
.A(n_2539),
.B(n_339),
.C(n_340),
.D(n_341),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2561),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2557),
.Y(n_2585)
);

O2A1O1Ixp33_ASAP7_75t_L g2586 ( 
.A1(n_2565),
.A2(n_2562),
.B(n_2570),
.C(n_2563),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2579),
.Y(n_2587)
);

BUFx12f_ASAP7_75t_L g2588 ( 
.A(n_2558),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2580),
.B(n_2546),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_2574),
.Y(n_2590)
);

NOR4xp25_ASAP7_75t_L g2591 ( 
.A(n_2559),
.B(n_2536),
.C(n_2547),
.D(n_2519),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2575),
.B(n_2510),
.Y(n_2592)
);

AOI221xp5_ASAP7_75t_SL g2593 ( 
.A1(n_2573),
.A2(n_2522),
.B1(n_2517),
.B2(n_2515),
.C(n_2549),
.Y(n_2593)
);

BUFx2_ASAP7_75t_L g2594 ( 
.A(n_2578),
.Y(n_2594)
);

OAI221xp5_ASAP7_75t_SL g2595 ( 
.A1(n_2560),
.A2(n_2543),
.B1(n_2527),
.B2(n_2529),
.C(n_2551),
.Y(n_2595)
);

AOI221xp5_ASAP7_75t_L g2596 ( 
.A1(n_2583),
.A2(n_2548),
.B1(n_2523),
.B2(n_2555),
.C(n_2544),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2576),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2571),
.Y(n_2598)
);

INVx2_ASAP7_75t_SL g2599 ( 
.A(n_2556),
.Y(n_2599)
);

OAI22xp5_ASAP7_75t_SL g2600 ( 
.A1(n_2566),
.A2(n_2540),
.B1(n_2569),
.B2(n_2564),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2567),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_R g2602 ( 
.A(n_2572),
.B(n_2568),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_2581),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2582),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2577),
.Y(n_2605)
);

NAND3xp33_ASAP7_75t_SL g2606 ( 
.A(n_2585),
.B(n_2550),
.C(n_341),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2599),
.A2(n_340),
.B1(n_342),
.B2(n_343),
.Y(n_2607)
);

AOI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2588),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2603),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_2609)
);

OAI221xp5_ASAP7_75t_SL g2610 ( 
.A1(n_2596),
.A2(n_2591),
.B1(n_2586),
.B2(n_2587),
.C(n_2589),
.Y(n_2610)
);

AOI32xp33_ASAP7_75t_L g2611 ( 
.A1(n_2592),
.A2(n_2601),
.A3(n_2590),
.B1(n_2594),
.B2(n_2584),
.Y(n_2611)
);

AOI322xp5_ASAP7_75t_L g2612 ( 
.A1(n_2593),
.A2(n_2597),
.A3(n_2605),
.B1(n_2598),
.B2(n_2604),
.C1(n_2595),
.C2(n_2602),
.Y(n_2612)
);

AOI22x1_ASAP7_75t_L g2613 ( 
.A1(n_2600),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2600),
.Y(n_2614)
);

OAI22xp33_ASAP7_75t_SL g2615 ( 
.A1(n_2599),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_2615)
);

O2A1O1Ixp5_ASAP7_75t_L g2616 ( 
.A1(n_2589),
.A2(n_351),
.B(n_352),
.C(n_353),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2599),
.B(n_351),
.Y(n_2617)
);

OAI322xp33_ASAP7_75t_L g2618 ( 
.A1(n_2599),
.A2(n_352),
.A3(n_353),
.B1(n_354),
.B2(n_355),
.C1(n_356),
.C2(n_357),
.Y(n_2618)
);

AOI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_2599),
.A2(n_354),
.B1(n_357),
.B2(n_358),
.C(n_359),
.Y(n_2619)
);

AOI322xp5_ASAP7_75t_L g2620 ( 
.A1(n_2599),
.A2(n_358),
.A3(n_360),
.B1(n_361),
.B2(n_362),
.C1(n_363),
.C2(n_364),
.Y(n_2620)
);

OAI221xp5_ASAP7_75t_L g2621 ( 
.A1(n_2599),
.A2(n_360),
.B1(n_361),
.B2(n_363),
.C(n_364),
.Y(n_2621)
);

AOI221xp5_ASAP7_75t_SL g2622 ( 
.A1(n_2586),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.C(n_368),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_2589),
.Y(n_2623)
);

AOI322xp5_ASAP7_75t_L g2624 ( 
.A1(n_2599),
.A2(n_365),
.A3(n_366),
.B1(n_367),
.B2(n_369),
.C1(n_370),
.C2(n_371),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2617),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2615),
.Y(n_2626)
);

AOI22x1_ASAP7_75t_L g2627 ( 
.A1(n_2614),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_2627)
);

AO22x1_ASAP7_75t_SL g2628 ( 
.A1(n_2623),
.A2(n_372),
.B1(n_374),
.B2(n_375),
.Y(n_2628)
);

OAI22x1_ASAP7_75t_L g2629 ( 
.A1(n_2613),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2606),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2621),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2622),
.B(n_381),
.Y(n_2632)
);

OAI22xp33_ASAP7_75t_SL g2633 ( 
.A1(n_2610),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_2633)
);

AO22x2_ASAP7_75t_L g2634 ( 
.A1(n_2612),
.A2(n_2611),
.B1(n_2616),
.B2(n_2619),
.Y(n_2634)
);

AOI211xp5_ASAP7_75t_SL g2635 ( 
.A1(n_2633),
.A2(n_2618),
.B(n_2607),
.C(n_2609),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2628),
.Y(n_2636)
);

NAND4xp25_ASAP7_75t_SL g2637 ( 
.A(n_2630),
.B(n_2608),
.C(n_2624),
.D(n_2620),
.Y(n_2637)
);

OAI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2631),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.C(n_387),
.Y(n_2638)
);

NAND5xp2_ASAP7_75t_L g2639 ( 
.A(n_2625),
.B(n_2626),
.C(n_2632),
.D(n_2634),
.E(n_2629),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2636),
.Y(n_2640)
);

OAI22x1_ASAP7_75t_L g2641 ( 
.A1(n_2637),
.A2(n_2627),
.B1(n_2634),
.B2(n_389),
.Y(n_2641)
);

OA21x2_ASAP7_75t_L g2642 ( 
.A1(n_2638),
.A2(n_386),
.B(n_388),
.Y(n_2642)
);

AO22x2_ASAP7_75t_L g2643 ( 
.A1(n_2640),
.A2(n_2639),
.B1(n_2635),
.B2(n_390),
.Y(n_2643)
);

XOR2xp5_ASAP7_75t_L g2644 ( 
.A(n_2641),
.B(n_388),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2642),
.Y(n_2645)
);

OAI31xp33_ASAP7_75t_L g2646 ( 
.A1(n_2640),
.A2(n_389),
.A3(n_390),
.B(n_391),
.Y(n_2646)
);

OAI21x1_ASAP7_75t_SL g2647 ( 
.A1(n_2644),
.A2(n_392),
.B(n_394),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2643),
.Y(n_2648)
);

AOI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2645),
.A2(n_392),
.B(n_395),
.Y(n_2649)
);

OAI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2648),
.A2(n_2646),
.B(n_396),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2650),
.A2(n_2649),
.B1(n_2647),
.B2(n_397),
.Y(n_2651)
);

OAI21xp5_ASAP7_75t_L g2652 ( 
.A1(n_2651),
.A2(n_395),
.B(n_396),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2651),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_2653)
);

HB1xp67_ASAP7_75t_L g2654 ( 
.A(n_2652),
.Y(n_2654)
);

AOI221xp5_ASAP7_75t_L g2655 ( 
.A1(n_2654),
.A2(n_2653),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2655),
.A2(n_398),
.B(n_401),
.Y(n_2656)
);

AOI211xp5_ASAP7_75t_L g2657 ( 
.A1(n_2656),
.A2(n_402),
.B(n_403),
.C(n_404),
.Y(n_2657)
);


endmodule