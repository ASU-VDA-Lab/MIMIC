module fake_jpeg_10387_n_60 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_20),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_42)
);

OR2x4_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_2),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_29),
.B(n_33),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_40),
.C(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_38),
.B1(n_36),
.B2(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_50),
.B(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_7),
.C(n_8),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_51),
.C(n_47),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_54),
.B1(n_49),
.B2(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_9),
.Y(n_58)
);

AOI321xp33_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_21),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_19),
.Y(n_60)
);


endmodule