module fake_jpeg_5056_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_36),
.Y(n_72)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_17),
.B1(n_27),
.B2(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_49),
.B(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_57),
.B1(n_37),
.B2(n_21),
.Y(n_85)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_32),
.CON(n_57),
.SN(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_46),
.B1(n_29),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_37),
.B1(n_17),
.B2(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_18),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_19),
.C(n_28),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_91),
.B1(n_50),
.B2(n_42),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_80),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_38),
.B1(n_44),
.B2(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_85),
.B1(n_44),
.B2(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_26),
.B(n_24),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_25),
.B(n_26),
.C(n_19),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_24),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_53),
.B(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_19),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_99),
.C(n_90),
.Y(n_119)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_55),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_122),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_35),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_68),
.B1(n_63),
.B2(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_109),
.B1(n_86),
.B2(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_63),
.B1(n_70),
.B2(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_73),
.B1(n_44),
.B2(n_35),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_113),
.B1(n_123),
.B2(n_90),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_125),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_73),
.B(n_51),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_55),
.B(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_127),
.B1(n_89),
.B2(n_80),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_35),
.B1(n_60),
.B2(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_54),
.C(n_43),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_54),
.B1(n_14),
.B2(n_15),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_98),
.B1(n_93),
.B2(n_97),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_129),
.B(n_135),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_154),
.B1(n_118),
.B2(n_50),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_140),
.B1(n_145),
.B2(n_113),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_91),
.B1(n_74),
.B2(n_79),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_102),
.B1(n_104),
.B2(n_124),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_137),
.B(n_139),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_90),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_96),
.B1(n_81),
.B2(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_87),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_149),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_100),
.B(n_0),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_156),
.B(n_26),
.Y(n_165)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_153),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_76),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_76),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_83),
.B1(n_54),
.B2(n_14),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_54),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_26),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_164),
.C(n_172),
.Y(n_199)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_108),
.B1(n_103),
.B2(n_115),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_171),
.B1(n_179),
.B2(n_183),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_115),
.C(n_113),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_176),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_166),
.B(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_102),
.B1(n_104),
.B2(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_178),
.B1(n_135),
.B2(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_120),
.C(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_148),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_106),
.C(n_83),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_180),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_106),
.B(n_25),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_118),
.B1(n_43),
.B2(n_42),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_129),
.B(n_25),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_182),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_28),
.B1(n_23),
.B2(n_25),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_28),
.B1(n_23),
.B2(n_2),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_132),
.B1(n_153),
.B2(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_145),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_196),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_197),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_150),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_208),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_205),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_179),
.B1(n_161),
.B2(n_163),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_150),
.B1(n_136),
.B2(n_147),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_144),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_158),
.B(n_150),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_158),
.C(n_164),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_230),
.C(n_235),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_175),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_239),
.B(n_186),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_162),
.B(n_176),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_231),
.B1(n_238),
.B2(n_193),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_172),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_227),
.B1(n_194),
.B2(n_198),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_163),
.B1(n_136),
.B2(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_187),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_167),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_165),
.B(n_168),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_142),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_178),
.C(n_170),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_144),
.C(n_23),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_192),
.C(n_208),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_204),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_188),
.A2(n_16),
.B(n_15),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_262),
.B1(n_264),
.B2(n_220),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_256),
.B1(n_263),
.B2(n_216),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_218),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_237),
.CI(n_227),
.CON(n_272),
.SN(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_219),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_215),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_234),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_236),
.C(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_195),
.B1(n_194),
.B2(n_209),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_210),
.B1(n_212),
.B2(n_5),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_266),
.C(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_255),
.C(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_217),
.C(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_272),
.B(n_264),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_12),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_224),
.B1(n_214),
.B2(n_222),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_247),
.B(n_13),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_13),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_244),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_285),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_296),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_267),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_290),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_259),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_294),
.C(n_265),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_260),
.C(n_243),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_241),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_11),
.B1(n_3),
.B2(n_5),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_243),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_270),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_277),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_272),
.B(n_11),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_276),
.B1(n_11),
.B2(n_5),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_269),
.C(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_302),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_273),
.C(n_282),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_297),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_277),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_0),
.B(n_3),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_291),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_287),
.B1(n_292),
.B2(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_289),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_321),
.B(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_305),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_0),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_6),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_330),
.C(n_319),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_303),
.B(n_310),
.C(n_302),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_328),
.A2(n_331),
.B(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_300),
.Y(n_330)
);

OAI31xp33_ASAP7_75t_L g331 ( 
.A1(n_314),
.A2(n_301),
.A3(n_307),
.B(n_9),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_322),
.B(n_315),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_333),
.A2(n_334),
.B(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_7),
.C(n_8),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_336),
.A2(n_7),
.B(n_8),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.C(n_337),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_7),
.B(n_8),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_8),
.B(n_9),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_9),
.B(n_336),
.Y(n_343)
);


endmodule