module fake_jpeg_1058_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_20),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_37),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_22),
.B(n_20),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_13),
.B(n_14),
.C(n_23),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_39),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_14),
.B1(n_13),
.B2(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_29),
.B1(n_37),
.B2(n_18),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_48),
.B1(n_36),
.B2(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_26),
.B(n_34),
.C(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_49),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_36),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_64),
.B1(n_36),
.B2(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_11),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_26),
.B(n_17),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_48),
.C(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_7),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_81),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_82),
.B1(n_83),
.B2(n_68),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_49),
.B1(n_16),
.B2(n_3),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_49),
.B1(n_16),
.B2(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_61),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_68),
.B1(n_65),
.B2(n_60),
.C(n_82),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_73),
.C(n_77),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_103),
.C(n_60),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_72),
.B(n_81),
.C(n_87),
.D(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_52),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_72),
.B1(n_80),
.B2(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_105),
.B1(n_93),
.B2(n_90),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_60),
.C(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_78),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_106),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_99),
.B(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_100),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

OAI211xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_103),
.B(n_98),
.C(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_116),
.B(n_6),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_97),
.C(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_59),
.C(n_67),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_111),
.A3(n_110),
.B1(n_85),
.B2(n_84),
.C1(n_88),
.C2(n_67),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_1),
.C(n_4),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_115),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_125),
.B(n_5),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_122),
.B(n_5),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_126),
.Y(n_129)
);


endmodule