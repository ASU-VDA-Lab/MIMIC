module fake_jpeg_23786_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_0),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_16),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_10),
.B1(n_8),
.B2(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

NAND2x1_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_4),
.Y(n_18)
);

AOI222xp33_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_19),
.B1(n_6),
.B2(n_17),
.C1(n_14),
.C2(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_21),
.C(n_24),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_29),
.B(n_31),
.Y(n_36)
);

AOI321xp33_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_37),
.A3(n_34),
.B1(n_9),
.B2(n_5),
.C(n_4),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_19),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_5),
.B(n_9),
.Y(n_39)
);


endmodule