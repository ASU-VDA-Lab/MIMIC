module real_aes_15693_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_0), .Y(n_237) );
AND2x4_ASAP7_75t_L g110 ( .A(n_1), .B(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g178 ( .A(n_2), .Y(n_178) );
INVx1_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_4), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g867 ( .A(n_4), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_5), .B(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g106 ( .A(n_6), .B(n_20), .Y(n_106) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_7), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_8), .B(n_172), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_9), .B(n_172), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_10), .B(n_197), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_11), .A2(n_78), .B1(n_147), .B2(n_172), .Y(n_246) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_12), .A2(n_33), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_13), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_14), .B(n_187), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_15), .Y(n_533) );
AO32x2_ASAP7_75t_L g243 ( .A1(n_16), .A2(n_164), .A3(n_165), .B1(n_244), .B2(n_247), .Y(n_243) );
AO32x1_ASAP7_75t_L g281 ( .A1(n_16), .A2(n_164), .A3(n_165), .B1(n_244), .B2(n_247), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_17), .B(n_518), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_18), .B(n_164), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_19), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_21), .A2(n_39), .B1(n_175), .B2(n_187), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_22), .A2(n_87), .B1(n_147), .B2(n_155), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_23), .B(n_154), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_24), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_25), .B(n_210), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_26), .A2(n_58), .B1(n_155), .B2(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_27), .B(n_172), .Y(n_588) );
INVx2_ASAP7_75t_L g853 ( .A(n_28), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_29), .B(n_151), .Y(n_619) );
BUFx3_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
INVx1_ASAP7_75t_L g118 ( .A(n_30), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_31), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_32), .B(n_524), .Y(n_625) );
AND2x2_ASAP7_75t_L g539 ( .A(n_34), .B(n_524), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_35), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_36), .B(n_209), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_37), .B(n_518), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_38), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_40), .B(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_41), .A2(n_72), .B1(n_209), .B2(n_210), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_42), .B(n_252), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_43), .A2(n_188), .B(n_235), .C(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_44), .A2(n_74), .B1(n_147), .B2(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g143 ( .A(n_45), .Y(n_143) );
AND2x4_ASAP7_75t_L g161 ( .A(n_46), .B(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_47), .A2(n_48), .B1(n_155), .B2(n_175), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_49), .B(n_164), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_50), .B(n_524), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_51), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_52), .B(n_155), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_53), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g162 ( .A(n_54), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_55), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_56), .A2(n_235), .B(n_236), .C(n_238), .Y(n_234) );
NAND3xp33_ASAP7_75t_L g159 ( .A(n_57), .B(n_147), .C(n_157), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_59), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_60), .B(n_164), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_61), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g240 ( .A(n_62), .B(n_241), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_63), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_64), .B(n_151), .C(n_187), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_65), .A2(n_91), .B1(n_172), .B2(n_209), .Y(n_213) );
INVx2_ASAP7_75t_L g152 ( .A(n_66), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_67), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_68), .B(n_516), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_69), .B(n_172), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_70), .B(n_212), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_71), .A2(n_857), .B1(n_868), .B2(n_872), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_73), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_75), .B(n_191), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_76), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_77), .A2(n_86), .B1(n_518), .B2(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_79), .B(n_172), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_80), .B(n_157), .Y(n_156) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_81), .B(n_150), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_82), .A2(n_100), .B1(n_112), .B2(n_876), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_83), .B(n_185), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_84), .A2(n_98), .B1(n_155), .B2(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_85), .B(n_210), .Y(n_267) );
AOI22xp33_ASAP7_75t_SL g121 ( .A1(n_88), .A2(n_122), .B1(n_847), .B2(n_848), .Y(n_121) );
INVx1_ASAP7_75t_SL g848 ( .A(n_88), .Y(n_848) );
INVx1_ASAP7_75t_L g109 ( .A(n_89), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_89), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_90), .B(n_197), .Y(n_273) );
NAND2xp33_ASAP7_75t_L g571 ( .A(n_92), .B(n_150), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_93), .B(n_524), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_94), .B(n_150), .C(n_212), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_95), .B(n_516), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_96), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_97), .B(n_518), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
BUFx12f_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_SL g876 ( .A(n_102), .Y(n_876) );
OR2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g875 ( .A(n_104), .B(n_126), .Y(n_875) );
NOR2x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g855 ( .A(n_105), .Y(n_855) );
INVx1_ASAP7_75t_L g119 ( .A(n_106), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND3x2_ASAP7_75t_L g116 ( .A(n_108), .B(n_117), .C(n_119), .Y(n_116) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g126 ( .A(n_109), .Y(n_126) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_120), .Y(n_112) );
AOI31xp33_ASAP7_75t_L g866 ( .A1(n_113), .A2(n_128), .A3(n_859), .B(n_867), .Y(n_866) );
NOR2x1_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g863 ( .A(n_118), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_119), .B(n_855), .Y(n_854) );
AND2x6_ASAP7_75t_SL g861 ( .A(n_119), .B(n_862), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_849), .B(n_856), .Y(n_120) );
INVx1_ASAP7_75t_L g847 ( .A(n_122), .Y(n_847) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_127), .B(n_503), .Y(n_122) );
INVx8_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
BUFx8_ASAP7_75t_SL g846 ( .A(n_126), .Y(n_846) );
BUFx2_ASAP7_75t_L g865 ( .A(n_127), .Y(n_865) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_413), .Y(n_128) );
NAND4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_318), .C(n_345), .D(n_381), .Y(n_129) );
AOI221x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_223), .B1(n_257), .B2(n_293), .C(n_297), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_199), .C(n_221), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_166), .Y(n_134) );
INVx2_ASAP7_75t_L g258 ( .A(n_135), .Y(n_258) );
AND2x2_ASAP7_75t_L g431 ( .A(n_135), .B(n_375), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_135), .B(n_222), .Y(n_440) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g446 ( .A(n_136), .Y(n_446) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g291 ( .A(n_137), .Y(n_291) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g374 ( .A(n_138), .B(n_220), .Y(n_374) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B(n_163), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_139), .A2(n_144), .B(n_163), .Y(n_303) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_139), .A2(n_513), .B(n_523), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_139), .A2(n_544), .B(n_552), .Y(n_543) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_139), .A2(n_544), .B(n_552), .Y(n_642) );
OAI21xp33_ASAP7_75t_SL g733 ( .A1(n_139), .A2(n_513), .B(n_523), .Y(n_733) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g524 ( .A(n_140), .Y(n_524) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVx2_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_142), .Y(n_165) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_153), .B(n_160), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_SL g210 ( .A(n_147), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_147), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_148), .Y(n_150) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx1_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx1_ASAP7_75t_L g235 ( .A(n_148), .Y(n_235) );
INVx3_ASAP7_75t_L g516 ( .A(n_148), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_148), .Y(n_519) );
INVx2_ASAP7_75t_L g551 ( .A(n_150), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_171), .B1(n_173), .B2(n_174), .Y(n_170) );
INVx6_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_151), .A2(n_188), .B1(n_245), .B2(n_246), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g545 ( .A1(n_151), .A2(n_184), .B(n_546), .C(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_151), .A2(n_590), .B(n_591), .Y(n_589) );
BUFx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
INVx2_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx1_ASAP7_75t_L g212 ( .A(n_152), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_159), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp33_ASAP7_75t_L g536 ( .A1(n_155), .A2(n_516), .B1(n_537), .B2(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g596 ( .A(n_155), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_155), .A2(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
AOI31xp67_ASAP7_75t_L g168 ( .A1(n_160), .A2(n_169), .A3(n_170), .B(n_176), .Y(n_168) );
OAI21x1_ASAP7_75t_L g181 ( .A1(n_160), .A2(n_182), .B(n_189), .Y(n_181) );
OAI21x1_ASAP7_75t_L g513 ( .A1(n_160), .A2(n_514), .B(n_520), .Y(n_513) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_160), .A2(n_545), .B(n_548), .Y(n_544) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_160), .A2(n_557), .B(n_560), .Y(n_556) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_160), .B(n_165), .Y(n_576) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_160), .A2(n_586), .B(n_589), .Y(n_585) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_160), .A2(n_618), .B(n_621), .Y(n_617) );
BUFx10_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
INVx1_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
AO31x2_ASAP7_75t_L g249 ( .A1(n_161), .A2(n_206), .A3(n_250), .B(n_255), .Y(n_249) );
BUFx10_ASAP7_75t_L g529 ( .A(n_161), .Y(n_529) );
INVx2_ASAP7_75t_L g169 ( .A(n_164), .Y(n_169) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_165), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
BUFx3_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_165), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_SL g264 ( .A(n_165), .Y(n_264) );
INVx1_ASAP7_75t_SL g555 ( .A(n_165), .Y(n_555) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_166), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_166), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g444 ( .A(n_166), .Y(n_444) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
AND2x2_ASAP7_75t_L g222 ( .A(n_167), .B(n_205), .Y(n_222) );
INVx2_ASAP7_75t_L g300 ( .A(n_167), .Y(n_300) );
AND2x2_ASAP7_75t_L g365 ( .A(n_167), .B(n_303), .Y(n_365) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g220 ( .A(n_168), .Y(n_220) );
INVx3_ASAP7_75t_L g272 ( .A(n_172), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_172), .A2(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g624 ( .A(n_172), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_173), .A2(n_208), .B1(n_211), .B2(n_213), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_173), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_173), .A2(n_270), .B(n_271), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_173), .A2(n_535), .B1(n_595), .B2(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_175), .A2(n_187), .B1(n_231), .B2(n_232), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g292 ( .A(n_179), .Y(n_292) );
AND2x2_ASAP7_75t_L g302 ( .A(n_179), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g364 ( .A(n_179), .B(n_205), .Y(n_364) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_196), .Y(n_179) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_180), .A2(n_181), .B(n_196), .Y(n_202) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_180), .A2(n_585), .B(n_592), .Y(n_584) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_180), .A2(n_617), .B(n_625), .Y(n_616) );
OA21x2_ASAP7_75t_L g628 ( .A1(n_180), .A2(n_617), .B(n_625), .Y(n_628) );
OAI21x1_ASAP7_75t_L g631 ( .A1(n_180), .A2(n_585), .B(n_592), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_188), .Y(n_182) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g252 ( .A(n_187), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_188), .A2(n_515), .B(n_517), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_188), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_188), .A2(n_570), .B(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_188), .A2(n_587), .B(n_588), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B1(n_194), .B2(n_195), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_191), .A2(n_549), .B(n_550), .Y(n_548) );
INVx2_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_192), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx3_ASAP7_75t_L g238 ( .A(n_193), .Y(n_238) );
INVx2_ASAP7_75t_L g227 ( .A(n_197), .Y(n_227) );
NOR2xp67_ASAP7_75t_SL g527 ( .A(n_197), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_198), .A2(n_529), .A3(n_594), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g329 ( .A(n_199), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_203), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_201), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_201), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_201), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_201), .B(n_399), .Y(n_406) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g375 ( .A(n_202), .B(n_350), .Y(n_375) );
OR2x2_ASAP7_75t_L g377 ( .A(n_202), .B(n_303), .Y(n_377) );
INVx1_ASAP7_75t_L g436 ( .A(n_202), .Y(n_436) );
BUFx2_ASAP7_75t_L g450 ( .A(n_202), .Y(n_450) );
OR2x2_ASAP7_75t_L g478 ( .A(n_202), .B(n_205), .Y(n_478) );
INVx1_ASAP7_75t_L g497 ( .A(n_203), .Y(n_497) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g344 ( .A(n_204), .Y(n_344) );
OR2x2_ASAP7_75t_L g357 ( .A(n_204), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g376 ( .A(n_204), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_219), .Y(n_204) );
INVx2_ASAP7_75t_L g296 ( .A(n_205), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_205), .B(n_219), .Y(n_312) );
INVx1_ASAP7_75t_L g350 ( .A(n_205), .Y(n_350) );
INVx1_ASAP7_75t_L g393 ( .A(n_205), .Y(n_393) );
AND2x2_ASAP7_75t_L g435 ( .A(n_205), .B(n_436), .Y(n_435) );
AO31x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .A3(n_214), .B(n_216), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_209), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_SL g247 ( .A(n_215), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g241 ( .A(n_218), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_218), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g491 ( .A(n_221), .Y(n_491) );
AND2x4_ASAP7_75t_L g429 ( .A(n_222), .B(n_289), .Y(n_429) );
INVx2_ASAP7_75t_L g458 ( .A(n_222), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_222), .B(n_450), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_223), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_242), .Y(n_223) );
AND2x2_ASAP7_75t_L g369 ( .A(n_224), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g390 ( .A(n_224), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g261 ( .A(n_225), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g285 ( .A(n_225), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g316 ( .A(n_225), .Y(n_316) );
AND2x2_ASAP7_75t_L g356 ( .A(n_225), .B(n_248), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_225), .B(n_340), .Y(n_397) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g309 ( .A(n_226), .Y(n_309) );
AOI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_240), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_234), .B(n_239), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_230), .B(n_233), .Y(n_229) );
AOI21x1_ASAP7_75t_L g621 ( .A1(n_233), .A2(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g574 ( .A(n_235), .Y(n_574) );
INVx2_ASAP7_75t_L g254 ( .A(n_238), .Y(n_254) );
INVx2_ASAP7_75t_L g535 ( .A(n_238), .Y(n_535) );
INVx3_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
AND2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_315), .Y(n_320) );
AND2x2_ASAP7_75t_L g475 ( .A(n_242), .B(n_279), .Y(n_475) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_248), .Y(n_242) );
INVx1_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
AND2x2_ASAP7_75t_L g354 ( .A(n_243), .B(n_262), .Y(n_354) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_247), .A2(n_266), .B(n_269), .Y(n_265) );
AND2x4_ASAP7_75t_L g307 ( .A(n_248), .B(n_308), .Y(n_307) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g280 ( .A(n_249), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g317 ( .A(n_249), .B(n_281), .Y(n_317) );
AND2x2_ASAP7_75t_L g327 ( .A(n_249), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_249), .B(n_262), .Y(n_379) );
AND2x2_ASAP7_75t_L g385 ( .A(n_249), .B(n_309), .Y(n_385) );
AOI21x1_ASAP7_75t_L g266 ( .A1(n_254), .A2(n_267), .B(n_268), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_254), .A2(n_521), .B(n_522), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_276), .Y(n_257) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_258), .A2(n_419), .B(n_423), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_258), .B(n_449), .Y(n_496) );
NAND2x1_ASAP7_75t_SL g259 ( .A(n_260), .B(n_274), .Y(n_259) );
INVx1_ASAP7_75t_L g502 ( .A(n_260), .Y(n_502) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx2_ASAP7_75t_L g279 ( .A(n_262), .Y(n_279) );
INVx2_ASAP7_75t_L g284 ( .A(n_262), .Y(n_284) );
INVxp67_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
AND2x2_ASAP7_75t_L g325 ( .A(n_262), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g336 ( .A(n_262), .B(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g340 ( .A(n_262), .Y(n_340) );
INVx1_ASAP7_75t_L g358 ( .A(n_262), .Y(n_358) );
OR2x2_ASAP7_75t_L g391 ( .A(n_262), .B(n_326), .Y(n_391) );
INVx1_ASAP7_75t_L g462 ( .A(n_262), .Y(n_462) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_273), .Y(n_263) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI21xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_282), .B(n_287), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_278), .A2(n_401), .B1(n_403), .B2(n_406), .Y(n_400) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_279), .B(n_327), .Y(n_361) );
BUFx2_ASAP7_75t_L g420 ( .A(n_279), .Y(n_420) );
INVx2_ASAP7_75t_L g370 ( .A(n_280), .Y(n_370) );
OR2x2_ASAP7_75t_L g454 ( .A(n_280), .B(n_284), .Y(n_454) );
INVx1_ASAP7_75t_L g286 ( .A(n_281), .Y(n_286) );
INVx1_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
NOR2x1p5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_284), .Y(n_405) );
OR2x2_ASAP7_75t_L g489 ( .A(n_284), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g492 ( .A(n_284), .B(n_327), .Y(n_492) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_285), .Y(n_455) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_289), .B(n_349), .Y(n_411) );
AND2x2_ASAP7_75t_L g501 ( .A(n_289), .B(n_299), .Y(n_501) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g410 ( .A(n_290), .B(n_299), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g367 ( .A(n_291), .B(n_300), .Y(n_367) );
AND2x2_ASAP7_75t_L g402 ( .A(n_291), .B(n_296), .Y(n_402) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g321 ( .A(n_294), .B(n_302), .Y(n_321) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g461 ( .A(n_296), .B(n_462), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_310), .B2(n_313), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_298), .A2(n_499), .B(n_500), .C(n_502), .Y(n_498) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g349 ( .A(n_300), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g417 ( .A(n_300), .Y(n_417) );
OR2x2_ASAP7_75t_L g464 ( .A(n_301), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g319 ( .A(n_305), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g422 ( .A(n_308), .Y(n_422) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
INVx1_ASAP7_75t_L g409 ( .A(n_309), .Y(n_409) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g465 ( .A(n_312), .Y(n_465) );
AND2x2_ASAP7_75t_L g487 ( .A(n_312), .B(n_450), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_313), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g339 ( .A(n_317), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g395 ( .A(n_317), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g490 ( .A(n_317), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B1(n_322), .B2(n_329), .C(n_330), .Y(n_318) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx2_ASAP7_75t_L g412 ( .A(n_325), .Y(n_412) );
BUFx2_ASAP7_75t_L g432 ( .A(n_327), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_338), .B(n_341), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
AND2x2_ASAP7_75t_L g474 ( .A(n_333), .B(n_396), .Y(n_474) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
AND2x2_ASAP7_75t_L g470 ( .A(n_335), .B(n_340), .Y(n_470) );
INVx1_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B(n_359), .C(n_371), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .B1(n_355), .B2(n_357), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
BUFx2_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
AND2x2_ASAP7_75t_L g480 ( .A(n_354), .B(n_422), .Y(n_480) );
OAI21xp33_ASAP7_75t_L g483 ( .A1(n_355), .A2(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B1(n_366), .B2(n_368), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_362), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g434 ( .A(n_367), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g421 ( .A(n_370), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_370), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_376), .B(n_378), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
AND2x2_ASAP7_75t_L g448 ( .A(n_373), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g485 ( .A(n_373), .B(n_450), .Y(n_485) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
OR2x2_ASAP7_75t_L g477 ( .A(n_374), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g392 ( .A(n_377), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g424 ( .A(n_377), .Y(n_424) );
OR2x2_ASAP7_75t_L g457 ( .A(n_377), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_400), .C(n_407), .Y(n_381) );
OAI322xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .A3(n_388), .B1(n_390), .B2(n_392), .C1(n_394), .C2(n_398), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_384), .A2(n_424), .B(n_460), .C(n_463), .Y(n_459) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g404 ( .A(n_385), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
AND2x4_ASAP7_75t_L g469 ( .A(n_385), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_387), .A2(n_425), .A3(n_439), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_393), .B(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_411), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_471), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_418), .B(n_426), .C(n_451), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_419), .A2(n_494), .B(n_495), .C(n_497), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_421), .A2(n_474), .A3(n_475), .B(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx2_ASAP7_75t_L g433 ( .A(n_425), .Y(n_433) );
NAND4xp25_ASAP7_75t_SL g426 ( .A(n_427), .B(n_430), .C(n_438), .D(n_447), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI32xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .A3(n_433), .B1(n_434), .B2(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
INVx1_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_459), .C(n_466), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_455), .B(n_456), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_460), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_483), .C(n_493), .D(n_498), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_479), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_474), .A2(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_491), .B2(n_492), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_490), .Y(n_499) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_846), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_505), .B(n_741), .Y(n_504) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_676), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_600), .C(n_649), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_540), .B(n_564), .C(n_581), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g815 ( .A(n_509), .B(n_734), .Y(n_815) );
OR2x2_ASAP7_75t_L g826 ( .A(n_509), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_510), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g717 ( .A(n_510), .B(n_607), .Y(n_717) );
AND2x2_ASAP7_75t_L g838 ( .A(n_510), .B(n_648), .Y(n_838) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_525), .Y(n_510) );
INVx2_ASAP7_75t_L g668 ( .A(n_511), .Y(n_668) );
AND2x2_ASAP7_75t_L g683 ( .A(n_511), .B(n_635), .Y(n_683) );
AND2x2_ASAP7_75t_L g692 ( .A(n_511), .B(n_566), .Y(n_692) );
AND2x2_ASAP7_75t_L g761 ( .A(n_511), .B(n_647), .Y(n_761) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g579 ( .A(n_512), .Y(n_579) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g732 ( .A(n_525), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g580 ( .A(n_526), .B(n_554), .Y(n_580) );
INVx2_ASAP7_75t_L g605 ( .A(n_526), .Y(n_605) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_530), .B(n_539), .Y(n_526) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g769 ( .A(n_540), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_553), .Y(n_541) );
INVx1_ASAP7_75t_L g789 ( .A(n_542), .Y(n_789) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g627 ( .A(n_543), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g710 ( .A(n_543), .B(n_616), .Y(n_710) );
AND2x2_ASAP7_75t_L g636 ( .A(n_553), .B(n_579), .Y(n_636) );
INVxp67_ASAP7_75t_L g785 ( .A(n_553), .Y(n_785) );
OR2x2_ASAP7_75t_L g827 ( .A(n_553), .B(n_566), .Y(n_827) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_563), .Y(n_554) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_577), .Y(n_564) );
INVx1_ASAP7_75t_L g682 ( .A(n_565), .Y(n_682) );
AND2x2_ASAP7_75t_L g836 ( .A(n_565), .B(n_732), .Y(n_836) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g608 ( .A(n_566), .Y(n_608) );
INVx4_ASAP7_75t_L g647 ( .A(n_566), .Y(n_647) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B(n_576), .Y(n_568) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g663 ( .A(n_578), .B(n_646), .Y(n_663) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g700 ( .A(n_579), .B(n_648), .Y(n_700) );
INVx2_ASAP7_75t_L g666 ( .A(n_580), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_580), .B(n_671), .Y(n_834) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_583), .B(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g819 ( .A(n_583), .Y(n_819) );
AND2x2_ASAP7_75t_L g833 ( .A(n_583), .B(n_655), .Y(n_833) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
AND2x2_ASAP7_75t_L g768 ( .A(n_584), .B(n_675), .Y(n_768) );
OR2x2_ASAP7_75t_L g805 ( .A(n_584), .B(n_593), .Y(n_805) );
AND2x2_ASAP7_75t_L g615 ( .A(n_593), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g629 ( .A(n_593), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g675 ( .A(n_593), .Y(n_675) );
OR2x2_ASAP7_75t_L g688 ( .A(n_593), .B(n_628), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_593), .B(n_628), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_610), .B(n_632), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI31xp33_ASAP7_75t_L g678 ( .A1(n_602), .A2(n_679), .A3(n_681), .B(n_684), .Y(n_678) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
AND2x2_ASAP7_75t_L g691 ( .A(n_603), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g701 ( .A(n_604), .Y(n_701) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_604), .Y(n_707) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g635 ( .A(n_605), .Y(n_635) );
AND2x2_ASAP7_75t_L g664 ( .A(n_605), .B(n_648), .Y(n_664) );
INVx2_ASAP7_75t_L g714 ( .A(n_605), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_606), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g739 ( .A(n_607), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g788 ( .A(n_607), .B(n_789), .Y(n_788) );
AOI33xp33_ASAP7_75t_L g843 ( .A1(n_607), .A2(n_673), .A3(n_683), .B1(n_710), .B2(n_819), .B3(n_844), .Y(n_843) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g648 ( .A(n_609), .Y(n_648) );
INVx1_ASAP7_75t_L g735 ( .A(n_609), .Y(n_735) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_626), .Y(n_611) );
INVx2_ASAP7_75t_L g643 ( .A(n_612), .Y(n_643) );
AND2x2_ASAP7_75t_L g724 ( .A(n_612), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g686 ( .A(n_613), .Y(n_686) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g754 ( .A(n_614), .B(n_641), .Y(n_754) );
AND2x2_ASAP7_75t_L g704 ( .A(n_615), .B(n_698), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_615), .B(n_722), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_615), .B(n_754), .Y(n_803) );
AND2x2_ASAP7_75t_L g640 ( .A(n_616), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g659 ( .A(n_616), .B(n_654), .Y(n_659) );
INVx1_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g729 ( .A(n_627), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_627), .B(n_822), .Y(n_824) );
AND2x2_ASAP7_75t_L g837 ( .A(n_627), .B(n_653), .Y(n_837) );
AND2x2_ASAP7_75t_L g655 ( .A(n_628), .B(n_641), .Y(n_655) );
INVx2_ASAP7_75t_L g637 ( .A(n_629), .Y(n_637) );
AND2x2_ASAP7_75t_L g751 ( .A(n_629), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g810 ( .A(n_629), .B(n_722), .Y(n_810) );
BUFx2_ASAP7_75t_L g792 ( .A(n_630), .Y(n_792) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g654 ( .A(n_631), .Y(n_654) );
OAI32xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .A3(n_638), .B1(n_643), .B2(n_644), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx2_ASAP7_75t_L g740 ( .A(n_635), .Y(n_740) );
AND2x2_ASAP7_75t_L g770 ( .A(n_635), .B(n_692), .Y(n_770) );
AND2x2_ASAP7_75t_L g712 ( .A(n_636), .B(n_713), .Y(n_712) );
AND3x2_ASAP7_75t_L g719 ( .A(n_636), .B(n_646), .C(n_714), .Y(n_719) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_639), .A2(n_661), .B1(n_670), .B2(n_672), .Y(n_669) );
OAI322xp33_ASAP7_75t_L g817 ( .A1(n_639), .A2(n_738), .A3(n_818), .B1(n_819), .B2(n_820), .C1(n_821), .C2(n_824), .Y(n_817) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g839 ( .A(n_640), .B(n_822), .Y(n_839) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_641), .Y(n_658) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_641), .Y(n_698) );
BUFx3_ASAP7_75t_L g722 ( .A(n_641), .Y(n_722) );
INVx1_ASAP7_75t_L g748 ( .A(n_641), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_641), .Y(n_752) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g706 ( .A(n_645), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g757 ( .A(n_646), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_646), .B(n_714), .Y(n_808) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2x1_ASAP7_75t_L g667 ( .A(n_647), .B(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g671 ( .A(n_647), .Y(n_671) );
AND2x2_ASAP7_75t_L g713 ( .A(n_647), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g734 ( .A(n_647), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_648), .B(n_761), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_656), .B(n_660), .C(n_669), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI31xp33_ASAP7_75t_L g811 ( .A1(n_651), .A2(n_812), .A3(n_814), .B(n_815), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .Y(n_651) );
AND2x4_ASAP7_75t_L g764 ( .A(n_652), .B(n_673), .Y(n_764) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_653), .Y(n_696) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g780 ( .A(n_654), .B(n_674), .Y(n_780) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .Y(n_660) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g820 ( .A(n_663), .Y(n_820) );
AND2x2_ASAP7_75t_L g680 ( .A(n_664), .B(n_671), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g749 ( .A1(n_665), .A2(n_750), .B1(n_753), .B2(n_755), .Y(n_749) );
OR2x6_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_SL g807 ( .A(n_668), .Y(n_807) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g777 ( .A(n_673), .B(n_722), .Y(n_777) );
INVx2_ASAP7_75t_L g823 ( .A(n_673), .Y(n_823) );
AND2x4_ASAP7_75t_L g831 ( .A(n_673), .B(n_752), .Y(n_831) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_693), .C(n_723), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_689), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_680), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AND2x4_ASAP7_75t_L g744 ( .A(n_682), .B(n_699), .Y(n_744) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_685), .B(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
AND2x2_ASAP7_75t_L g775 ( .A(n_687), .B(n_754), .Y(n_775) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_688), .Y(n_695) );
INVx1_ASAP7_75t_L g813 ( .A(n_688), .Y(n_813) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g842 ( .A(n_691), .Y(n_842) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_692), .Y(n_727) );
AOI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B(n_702), .C(n_715), .Y(n_693) );
NOR3x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .C(n_697), .Y(n_694) );
NAND2x1_ASAP7_75t_L g763 ( .A(n_697), .B(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NOR2x1p5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B1(n_708), .B2(n_711), .Y(n_702) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g796 ( .A(n_707), .Y(n_796) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g791 ( .A(n_710), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g845 ( .A(n_713), .Y(n_845) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g799 ( .A(n_720), .Y(n_799) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g726 ( .A(n_722), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_722), .B(n_780), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B(n_728), .Y(n_723) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_726), .B(n_813), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_736), .B2(n_738), .Y(n_728) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g781 ( .A(n_731), .Y(n_781) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g756 ( .A(n_732), .B(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g773 ( .A(n_733), .Y(n_773) );
INVx1_ASAP7_75t_L g793 ( .A(n_734), .Y(n_793) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_797), .Y(n_741) );
NAND3xp33_ASAP7_75t_SL g742 ( .A(n_743), .B(n_758), .C(n_771), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_749), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g804 ( .A(n_747), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g801 ( .A(n_756), .B(n_784), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B1(n_765), .B2(n_769), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g814 ( .A(n_764), .Y(n_814) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_766), .A2(n_787), .B(n_790), .Y(n_786) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_782), .B1(n_786), .B2(n_794), .Y(n_771) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B(n_776), .Y(n_772) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g841 ( .A(n_777), .Y(n_841) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g830 ( .A(n_780), .Y(n_830) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx2_ASAP7_75t_L g822 ( .A(n_792), .Y(n_822) );
INVxp67_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_816), .Y(n_797) );
AOI211xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B(n_802), .C(n_811), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .B(n_806), .C(n_809), .Y(n_802) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_825), .C(n_840), .Y(n_816) );
OR2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_828), .B1(n_832), .B2(n_834), .C(n_835), .Y(n_825) );
NOR2xp67_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_835) );
OAI21xp33_ASAP7_75t_SL g840 ( .A1(n_841), .A2(n_842), .B(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
BUFx12f_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AND2x6_ASAP7_75t_SL g851 ( .A(n_852), .B(n_854), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx3_ASAP7_75t_L g871 ( .A(n_853), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_853), .B(n_874), .Y(n_873) );
OAI21x1_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_864), .B(n_866), .Y(n_857) );
INVx5_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
CKINVDCx11_ASAP7_75t_R g869 ( .A(n_870), .Y(n_869) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
BUFx10_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
endmodule