module fake_jpeg_26802_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_40),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_64),
.Y(n_81)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_58),
.B1(n_63),
.B2(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_86),
.B1(n_54),
.B2(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_56),
.B1(n_63),
.B2(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_90),
.B1(n_59),
.B2(n_66),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_56),
.B1(n_61),
.B2(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_51),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_55),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_1),
.B(n_3),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_61),
.B1(n_68),
.B2(n_65),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_60),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_78),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_88),
.B(n_50),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_14),
.B(n_16),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_62),
.B1(n_79),
.B2(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_97),
.B1(n_103),
.B2(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_120),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_24),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_123),
.C(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_12),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_109),
.C(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_13),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_108),
.B(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_17),
.C(n_19),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_33),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_21),
.B(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_26),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_140),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_142),
.B1(n_138),
.B2(n_131),
.C(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_128),
.B1(n_127),
.B2(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

OAI31xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_143),
.A3(n_39),
.B(n_41),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_46),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_38),
.Y(n_154)
);


endmodule