module real_aes_7615_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
AOI21xp5_ASAP7_75t_L g9 ( .A1(n_0), .A2(n_10), .B(n_22), .Y(n_9) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g27 ( .A(n_2), .Y(n_27) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_3), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_4), .B(n_29), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g31 ( .A(n_6), .Y(n_31) );
INVx1_ASAP7_75t_L g30 ( .A(n_7), .Y(n_30) );
INVx1_ASAP7_75t_L g21 ( .A(n_8), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_11), .B(n_16), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g11 ( .A(n_12), .B(n_13), .Y(n_11) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_17), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_18), .B(n_20), .Y(n_17) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_19), .B(n_25), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_23), .Y(n_22) );
OR2x2_ASAP7_75t_SL g23 ( .A(n_24), .B(n_26), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_27), .B(n_28), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_30), .B(n_31), .Y(n_29) );
endmodule