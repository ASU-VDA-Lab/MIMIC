module fake_jpeg_17614_n_83 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_12),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_30),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_13),
.C(n_15),
.Y(n_30)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_22),
.Y(n_31)
);

FAx1_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_42),
.CI(n_21),
.CON(n_52),
.SN(n_52)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_36),
.B1(n_41),
.B2(n_17),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_22),
.B(n_17),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_39),
.B(n_43),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_40),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_20),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_22),
.B1(n_18),
.B2(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_11),
.B1(n_17),
.B2(n_19),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_21),
.B1(n_19),
.B2(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_9),
.B1(n_16),
.B2(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.C(n_1),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_14),
.C(n_15),
.Y(n_54)
);

OAI322xp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_31),
.A3(n_42),
.B1(n_35),
.B2(n_34),
.C1(n_39),
.C2(n_33),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_47),
.B(n_48),
.Y(n_64)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_38),
.B(n_36),
.C(n_39),
.D(n_3),
.Y(n_57)
);

XOR2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_54),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_7),
.C(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_57),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_47),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

AO221x1_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_78),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_80),
.B(n_51),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_69),
.B(n_49),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_2),
.C(n_4),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_4),
.Y(n_83)
);


endmodule