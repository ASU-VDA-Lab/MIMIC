module fake_jpeg_1973_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx12f_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_0),
.CON(n_53),
.SN(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_50),
.B1(n_40),
.B2(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_50),
.B1(n_47),
.B2(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_42),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_53),
.B(n_44),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_4),
.C(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_77),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_45),
.B1(n_39),
.B2(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_81),
.B1(n_61),
.B2(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_79),
.B1(n_66),
.B2(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

BUFx2_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_65),
.B1(n_66),
.B2(n_6),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_91),
.B1(n_9),
.B2(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_8),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_80),
.B1(n_73),
.B2(n_72),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_81),
.B(n_70),
.C(n_82),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_18),
.B(n_29),
.C(n_28),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_22),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_71),
.B1(n_66),
.B2(n_10),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_89),
.B1(n_13),
.B2(n_14),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_21),
.C(n_31),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_20),
.C(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_108),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_11),
.B1(n_17),
.B2(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_8),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_9),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_89),
.B1(n_14),
.B2(n_16),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_102),
.B1(n_98),
.B2(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_11),
.B(n_16),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_23),
.B(n_121),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_124),
.A3(n_117),
.B1(n_113),
.B2(n_115),
.C1(n_114),
.C2(n_122),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_103),
.A3(n_104),
.B1(n_17),
.B2(n_25),
.C1(n_27),
.C2(n_24),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_129),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_131),
.B(n_125),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_119),
.C(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_126),
.B(n_130),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_128),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_125),
.Y(n_143)
);


endmodule