module fake_ariane_1907_n_1680 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1680);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1680;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_737;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_380;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_677;
wire n_439;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_266),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_365),
.Y(n_369)
);

INVxp33_ASAP7_75t_R g370 ( 
.A(n_331),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_65),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_257),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_159),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_232),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_41),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_45),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_16),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_127),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_46),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_244),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_108),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_45),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_243),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_55),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_205),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_229),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_175),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_116),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_190),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_267),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_292),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_126),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_29),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_224),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_132),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_101),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_245),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_3),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_288),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_319),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_146),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_153),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_265),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_152),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_143),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_88),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_183),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_66),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_223),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_131),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_76),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_258),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_141),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_114),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_164),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_125),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_147),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_311),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_57),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_203),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_113),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_343),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_249),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_196),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_71),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_66),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_24),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_34),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_333),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_344),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_320),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_149),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_120),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_324),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_80),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_192),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_254),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_75),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_182),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_202),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_33),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_285),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_7),
.Y(n_448)
);

BUFx8_ASAP7_75t_SL g449 ( 
.A(n_34),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_184),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_9),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_276),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_6),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_51),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_130),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_129),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_111),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_291),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_67),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_300),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_51),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_94),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_16),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_151),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_329),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_119),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_49),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_339),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_247),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_123),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_72),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_363),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_359),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_90),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_49),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_133),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_156),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_142),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_23),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_271),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_235),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_294),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_209),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_81),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_335),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_253),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_74),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_342),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_318),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_345),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_358),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_268),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_214),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_352),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_77),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_118),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_264),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_240),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_50),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_40),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_100),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_86),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_315),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_193),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_112),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_137),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_33),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_91),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_36),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_63),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_30),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_5),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_304),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_31),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_15),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_138),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_124),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_367),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_115),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_325),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_134),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_168),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_360),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_155),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_56),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_144),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_89),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_12),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_39),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_165),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_93),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_280),
.Y(n_533)
);

BUFx8_ASAP7_75t_SL g534 ( 
.A(n_173),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_27),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_176),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_12),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_279),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_77),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_82),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_219),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_208),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_44),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_356),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_261),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_273),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_204),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_256),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_323),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_70),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_269),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_166),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_54),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_139),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_92),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_8),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_349),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_295),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_362),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_69),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_178),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_0),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_15),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_332),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_296),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_272),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_74),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_23),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_305),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_361),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_20),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_56),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_87),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_284),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_105),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_61),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_246),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_41),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_10),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_58),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_8),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_180),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_0),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_9),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_250),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_201),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_237),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_46),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_263),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_117),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g591 ( 
.A(n_42),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_35),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_299),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_73),
.Y(n_594)
);

BUFx8_ASAP7_75t_SL g595 ( 
.A(n_65),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_218),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_110),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_25),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_99),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_109),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_334),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_76),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_57),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_171),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_400),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_385),
.B(n_1),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_585),
.B(n_1),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_384),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_384),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_512),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_400),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_2),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_488),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_579),
.B(n_2),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_400),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_455),
.B(n_3),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_455),
.B(n_4),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_400),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_4),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_591),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_449),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_567),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_534),
.B(n_5),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_384),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_567),
.B(n_6),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_450),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_412),
.B(n_7),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_488),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_557),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_449),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_568),
.B(n_10),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_485),
.B(n_11),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_557),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_485),
.B(n_454),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_595),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_488),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_568),
.B(n_11),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_398),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_450),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_398),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_421),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_383),
.B(n_13),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_375),
.B(n_13),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_450),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_421),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_463),
.B(n_14),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_595),
.Y(n_650)
);

BUFx12f_ASAP7_75t_L g651 ( 
.A(n_481),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_562),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_389),
.B(n_14),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_457),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_568),
.B(n_458),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_481),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_458),
.B(n_17),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_405),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_371),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_405),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_562),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_457),
.B(n_17),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_368),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_369),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_393),
.B(n_18),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_394),
.B(n_18),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_534),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_505),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_505),
.B(n_19),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

INVx6_ASAP7_75t_L g675 ( 
.A(n_536),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_527),
.B(n_19),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_392),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_580),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_536),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_527),
.B(n_20),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_396),
.B(n_21),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_406),
.B(n_21),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_580),
.Y(n_684)
);

BUFx8_ASAP7_75t_SL g685 ( 
.A(n_452),
.Y(n_685)
);

INVx6_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_580),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_593),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_593),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_377),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_558),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_377),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_425),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_381),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_387),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_372),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_408),
.B(n_22),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_425),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_483),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_483),
.Y(n_701)
);

BUFx12f_ASAP7_75t_L g702 ( 
.A(n_423),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_376),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_419),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_466),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_466),
.B(n_22),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_420),
.B(n_24),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_378),
.B(n_25),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_379),
.B(n_26),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_397),
.Y(n_710)
);

BUFx8_ASAP7_75t_L g711 ( 
.A(n_370),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_402),
.B(n_26),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_427),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_428),
.B(n_27),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_429),
.B(n_28),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_434),
.B(n_28),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_441),
.B(n_29),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_456),
.B(n_470),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_415),
.B(n_30),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_486),
.Y(n_720)
);

BUFx8_ASAP7_75t_SL g721 ( 
.A(n_594),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_430),
.B(n_31),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_464),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_486),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_471),
.B(n_32),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_477),
.B(n_32),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_504),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_504),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_525),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_468),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_482),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_476),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_490),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_487),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_497),
.B(n_35),
.Y(n_736)
);

INVx5_ASAP7_75t_L g737 ( 
.A(n_545),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_501),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_508),
.B(n_36),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_503),
.B(n_37),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_401),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_431),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_SL g743 ( 
.A(n_492),
.B(n_37),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_522),
.B(n_38),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_524),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_38),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_511),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_432),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_546),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_537),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_551),
.B(n_555),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_401),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_556),
.B(n_39),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_564),
.B(n_40),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_433),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_566),
.B(n_42),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_560),
.B(n_572),
.Y(n_757)
);

INVx6_ASAP7_75t_L g758 ( 
.A(n_401),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_573),
.Y(n_759)
);

CKINVDCx6p67_ASAP7_75t_R g760 ( 
.A(n_492),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_574),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_575),
.B(n_43),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_404),
.Y(n_763)
);

BUFx8_ASAP7_75t_SL g764 ( 
.A(n_414),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_588),
.B(n_43),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_706),
.A2(n_416),
.B1(n_484),
.B2(n_445),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_659),
.A2(n_603),
.B1(n_602),
.B2(n_447),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_621),
.B(n_440),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_633),
.A2(n_461),
.B1(n_413),
.B2(n_577),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_706),
.A2(n_533),
.B1(n_446),
.B2(n_448),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_SL g771 ( 
.A1(n_743),
.A2(n_460),
.B1(n_462),
.B2(n_443),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_619),
.A2(n_480),
.B1(n_496),
.B2(n_472),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_743),
.A2(n_510),
.B1(n_513),
.B2(n_500),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_608),
.B(n_582),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_744),
.A2(n_705),
.B1(n_677),
.B2(n_612),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_641),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_623),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_624),
.A2(n_516),
.B1(n_526),
.B2(n_515),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_632),
.B(n_638),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_R g780 ( 
.A1(n_606),
.A2(n_535),
.B1(n_539),
.B2(n_529),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_610),
.A2(n_550),
.B1(n_553),
.B2(n_543),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_661),
.B(n_637),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_687),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_640),
.A2(n_599),
.B1(n_601),
.B2(n_597),
.Y(n_784)
);

AO22x2_ASAP7_75t_L g785 ( 
.A1(n_614),
.A2(n_646),
.B1(n_649),
.B2(n_619),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_641),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_624),
.A2(n_571),
.B1(n_576),
.B2(n_563),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_655),
.B(n_578),
.Y(n_788)
);

AO22x2_ASAP7_75t_L g789 ( 
.A1(n_665),
.A2(n_583),
.B1(n_584),
.B2(n_581),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_675),
.B(n_592),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_608),
.B(n_373),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_679),
.A2(n_598),
.B1(n_380),
.B2(n_382),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_687),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_692),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_692),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_675),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_692),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_607),
.A2(n_386),
.B1(n_388),
.B2(n_374),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_665),
.A2(n_48),
.B1(n_44),
.B2(n_47),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_630),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_693),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_705),
.A2(n_391),
.B1(n_395),
.B2(n_390),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_SL g805 ( 
.A1(n_607),
.A2(n_403),
.B1(n_407),
.B2(n_399),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_691),
.A2(n_409),
.B1(n_411),
.B2(n_410),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_686),
.B(n_417),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_686),
.B(n_691),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_658),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_751),
.A2(n_422),
.B1(n_424),
.B2(n_418),
.Y(n_811)
);

AO22x2_ASAP7_75t_L g812 ( 
.A1(n_673),
.A2(n_680),
.B1(n_676),
.B2(n_616),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_673),
.A2(n_435),
.B1(n_436),
.B2(n_426),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_698),
.B(n_437),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_693),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_748),
.A2(n_755),
.B1(n_629),
.B2(n_680),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_698),
.B(n_438),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_699),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_699),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_699),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_608),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_751),
.A2(n_653),
.B1(n_669),
.B2(n_645),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_SL g823 ( 
.A1(n_645),
.A2(n_442),
.B1(n_444),
.B2(n_439),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_698),
.B(n_451),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_653),
.A2(n_459),
.B1(n_465),
.B2(n_453),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_676),
.A2(n_467),
.B1(n_473),
.B2(n_469),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_622),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_669),
.A2(n_475),
.B1(n_478),
.B2(n_474),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_650),
.A2(n_760),
.B1(n_671),
.B2(n_656),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_625),
.B(n_479),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_628),
.A2(n_491),
.B1(n_493),
.B2(n_489),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_664),
.Y(n_833)
);

OAI22xp33_ASAP7_75t_R g834 ( 
.A1(n_670),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_628),
.A2(n_604),
.B1(n_600),
.B2(n_596),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_494),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_609),
.A2(n_590),
.B1(n_589),
.B2(n_587),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_605),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_666),
.B(n_667),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_666),
.B(n_495),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_668),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_700),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_684),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_642),
.B(n_498),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_656),
.A2(n_586),
.B1(n_570),
.B2(n_569),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_667),
.B(n_499),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_635),
.B(n_616),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_651),
.A2(n_565),
.B1(n_561),
.B2(n_559),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_696),
.B(n_502),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_681),
.A2(n_552),
.B1(n_549),
.B2(n_548),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_506),
.Y(n_851)
);

OA22x2_ASAP7_75t_L g852 ( 
.A1(n_637),
.A2(n_547),
.B1(n_542),
.B2(n_541),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_605),
.Y(n_853)
);

AO22x2_ASAP7_75t_L g854 ( 
.A1(n_617),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_647),
.B(n_507),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_656),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_52),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_700),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_695),
.A2(n_540),
.B1(n_538),
.B2(n_532),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_697),
.A2(n_531),
.B1(n_528),
.B2(n_523),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_SL g862 ( 
.A1(n_685),
.A2(n_521),
.B1(n_520),
.B2(n_519),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_674),
.B(n_509),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_717),
.A2(n_518),
.B1(n_517),
.B2(n_514),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_617),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_865)
);

INVx3_ASAP7_75t_SL g866 ( 
.A(n_627),
.Y(n_866)
);

OAI22xp33_ASAP7_75t_L g867 ( 
.A1(n_674),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_635),
.A2(n_627),
.B1(n_719),
.B2(n_712),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_681),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_611),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_777),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_793),
.Y(n_872)
);

XNOR2x2_ASAP7_75t_L g873 ( 
.A(n_769),
.B(n_721),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_783),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_847),
.B(n_712),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_809),
.B(n_790),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_794),
.Y(n_877)
);

XOR2xp5_ASAP7_75t_L g878 ( 
.A(n_862),
.B(n_711),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_796),
.B(n_674),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_782),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_776),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_786),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_795),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_822),
.B(n_682),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_801),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_797),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_808),
.B(n_682),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_804),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_827),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_779),
.Y(n_890)
);

INVxp33_ASAP7_75t_L g891 ( 
.A(n_768),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_799),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_802),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_815),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_812),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_821),
.B(n_682),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_818),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_819),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_820),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_842),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_788),
.B(n_704),
.Y(n_901)
);

XOR2xp5_ASAP7_75t_L g902 ( 
.A(n_766),
.B(n_711),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_831),
.B(n_757),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_856),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_859),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_807),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_779),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_810),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_833),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_868),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_866),
.B(n_683),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_841),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_839),
.B(n_660),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_844),
.B(n_735),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_870),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_855),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_812),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_816),
.B(n_694),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_829),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_857),
.B(n_702),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_829),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_840),
.B(n_846),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_863),
.B(n_719),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_829),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_838),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_849),
.B(n_660),
.Y(n_927)
);

AND2x6_ASAP7_75t_L g928 ( 
.A(n_826),
.B(n_722),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_838),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_851),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_781),
.B(n_742),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_838),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_791),
.A2(n_718),
.B(n_707),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_861),
.A2(n_707),
.B(n_683),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_792),
.B(n_688),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_814),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_824),
.B(n_722),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_853),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_854),
.B(n_739),
.Y(n_940)
);

INVx4_ASAP7_75t_SL g941 ( 
.A(n_853),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_785),
.Y(n_942)
);

INVxp33_ASAP7_75t_L g943 ( 
.A(n_775),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_785),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_813),
.B(n_662),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_852),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_836),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_837),
.B(n_689),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_817),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_848),
.B(n_784),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_784),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_767),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_767),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_770),
.B(n_764),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_806),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_774),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_800),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_798),
.B(n_662),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_800),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_860),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_864),
.B(n_713),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_772),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_SL g963 ( 
.A(n_773),
.B(n_787),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_854),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_949),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_885),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_963),
.B(n_803),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_930),
.B(n_811),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_923),
.B(n_769),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_930),
.B(n_771),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_888),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_908),
.Y(n_972)
);

AND2x2_ASAP7_75t_SL g973 ( 
.A(n_875),
.B(n_739),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_875),
.B(n_865),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_895),
.B(n_765),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_895),
.B(n_765),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_880),
.B(n_918),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_903),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_880),
.B(n_865),
.Y(n_979)
);

AND2x6_ASAP7_75t_L g980 ( 
.A(n_957),
.B(n_708),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_889),
.Y(n_981)
);

AND2x6_ASAP7_75t_SL g982 ( 
.A(n_940),
.B(n_858),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_918),
.B(n_789),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_909),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_949),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_964),
.B(n_714),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_940),
.B(n_858),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_910),
.B(n_789),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_912),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_901),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_910),
.B(n_709),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_903),
.B(n_753),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_915),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_872),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_940),
.B(n_750),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_949),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_876),
.B(n_750),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_871),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_942),
.B(n_731),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_934),
.B(n_731),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_923),
.B(n_701),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_949),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_906),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_914),
.B(n_938),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_917),
.B(n_805),
.Y(n_1005)
);

AND2x4_ASAP7_75t_SL g1006 ( 
.A(n_938),
.B(n_701),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_933),
.B(n_701),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_906),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_937),
.B(n_823),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_874),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_877),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_883),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_924),
.B(n_703),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_948),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_924),
.B(n_710),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_935),
.B(n_723),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_944),
.B(n_733),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_962),
.B(n_738),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_892),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_933),
.B(n_720),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_945),
.B(n_937),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_959),
.B(n_747),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_913),
.B(n_720),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_946),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_920),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_884),
.B(n_690),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_884),
.B(n_690),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_893),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_894),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_959),
.B(n_728),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_922),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_897),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_928),
.B(n_951),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_887),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_891),
.B(n_728),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_928),
.B(n_729),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_898),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_899),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_891),
.B(n_825),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_900),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_947),
.B(n_828),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_945),
.B(n_729),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_887),
.B(n_732),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_904),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_931),
.B(n_732),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_958),
.B(n_850),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_919),
.B(n_950),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_943),
.B(n_732),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_921),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_958),
.B(n_745),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_890),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_905),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_927),
.B(n_832),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_961),
.B(n_913),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_916),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_927),
.B(n_720),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_961),
.B(n_745),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_952),
.B(n_745),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_953),
.B(n_749),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_911),
.A2(n_715),
.B(n_714),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_925),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_956),
.B(n_749),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_907),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_926),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1034),
.B(n_928),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1055),
.B(n_928),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_994),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_966),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_985),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_981),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_SL g1072 ( 
.A(n_985),
.B(n_929),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1055),
.B(n_1000),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_994),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_1034),
.B(n_954),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_966),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_977),
.B(n_763),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1034),
.B(n_928),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_1034),
.B(n_985),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_973),
.B(n_778),
.Y(n_1080)
);

BUFx2_ASAP7_75t_SL g1081 ( 
.A(n_987),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1000),
.B(n_960),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_987),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1043),
.B(n_955),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_987),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_987),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1043),
.B(n_879),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_981),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_973),
.B(n_869),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1022),
.B(n_830),
.Y(n_1090)
);

CKINVDCx6p67_ASAP7_75t_R g1091 ( 
.A(n_1052),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_998),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_973),
.B(n_867),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_985),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_977),
.B(n_1049),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_995),
.B(n_881),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_1052),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_998),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1049),
.B(n_902),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_982),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_SL g1101 ( 
.A(n_974),
.B(n_834),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_995),
.B(n_882),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_L g1103 ( 
.A(n_965),
.B(n_996),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_991),
.B(n_932),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_991),
.B(n_936),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_985),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1064),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_985),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1001),
.B(n_939),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1001),
.B(n_896),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_966),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_982),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_978),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_971),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1064),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_998),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1025),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1023),
.B(n_941),
.Y(n_1119)
);

NAND2x1_ASAP7_75t_L g1120 ( 
.A(n_1026),
.B(n_758),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_R g1121 ( 
.A(n_979),
.B(n_780),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_SL g1122 ( 
.A(n_967),
.B(n_715),
.Y(n_1122)
);

BUFx4f_ASAP7_75t_L g1123 ( 
.A(n_980),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1023),
.B(n_941),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_971),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_1050),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1004),
.B(n_878),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1027),
.B(n_724),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1025),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1012),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_978),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1004),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1023),
.B(n_1031),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1012),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1035),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_971),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1015),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_965),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_965),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1023),
.B(n_941),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1015),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1031),
.B(n_749),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1030),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_975),
.B(n_759),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_996),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1046),
.B(n_641),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_990),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_972),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1073),
.B(n_974),
.Y(n_1149)
);

BUFx12f_ASAP7_75t_L g1150 ( 
.A(n_1071),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_SL g1151 ( 
.A(n_1091),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_1088),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1083),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1073),
.B(n_1028),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1100),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1097),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1119),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1119),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1124),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1124),
.B(n_996),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1107),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_1116),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1135),
.Y(n_1163)
);

INVx3_ASAP7_75t_SL g1164 ( 
.A(n_1126),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1082),
.B(n_1084),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1092),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_1066),
.B(n_1037),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1140),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1140),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1133),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1098),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1083),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1085),
.Y(n_1173)
);

CKINVDCx16_ASAP7_75t_R g1174 ( 
.A(n_1101),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1068),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_1132),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1070),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1074),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1130),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1086),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1112),
.Y(n_1182)
);

BUFx5_ASAP7_75t_L g1183 ( 
.A(n_1117),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1134),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1086),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1093),
.A2(n_969),
.B1(n_780),
.B2(n_834),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1093),
.A2(n_970),
.B1(n_968),
.B2(n_1047),
.Y(n_1187)
);

INVx6_ASAP7_75t_L g1188 ( 
.A(n_1138),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1095),
.A2(n_969),
.B1(n_988),
.B2(n_1047),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1141),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1143),
.Y(n_1192)
);

CKINVDCx8_ASAP7_75t_R g1193 ( 
.A(n_1081),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1077),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1133),
.Y(n_1195)
);

CKINVDCx6p67_ASAP7_75t_R g1196 ( 
.A(n_1127),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1069),
.Y(n_1197)
);

INVx5_ASAP7_75t_SL g1198 ( 
.A(n_1075),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1118),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1070),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1070),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1129),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1142),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_1101),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1113),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1138),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1131),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1142),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1106),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1106),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1147),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1138),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1114),
.B(n_1014),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1147),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1104),
.Y(n_1215)
);

INVx6_ASAP7_75t_L g1216 ( 
.A(n_1139),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1076),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1106),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1174),
.A2(n_873),
.B1(n_1089),
.B2(n_1082),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1151),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1150),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1199),
.Y(n_1222)
);

INVx6_ASAP7_75t_L g1223 ( 
.A(n_1194),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1186),
.A2(n_1084),
.B1(n_1099),
.B2(n_1048),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1202),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1186),
.A2(n_1048),
.B1(n_1089),
.B2(n_1014),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1166),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1175),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1157),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1171),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1209),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1152),
.Y(n_1232)
);

NAND2x1p5_ASAP7_75t_L g1233 ( 
.A(n_1172),
.B(n_1123),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_1157),
.Y(n_1234)
);

CKINVDCx14_ASAP7_75t_R g1235 ( 
.A(n_1155),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1172),
.B(n_1123),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1197),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1217),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1165),
.A2(n_1046),
.B1(n_1075),
.B2(n_988),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1204),
.A2(n_979),
.B1(n_1075),
.B2(n_1067),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1157),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1156),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1187),
.A2(n_1114),
.B1(n_1067),
.B2(n_1087),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1149),
.A2(n_1040),
.B1(n_968),
.B2(n_1080),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1154),
.A2(n_970),
.B1(n_1105),
.B2(n_1104),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1149),
.A2(n_1040),
.B1(n_1080),
.B2(n_983),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_1164),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1189),
.A2(n_983),
.B1(n_1078),
.B2(n_1066),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1205),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1193),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1178),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1179),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_SL g1253 ( 
.A(n_1207),
.Y(n_1253)
);

BUFx8_ASAP7_75t_L g1254 ( 
.A(n_1211),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1157),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_1105),
.B1(n_1061),
.B2(n_1087),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1198),
.A2(n_1122),
.B1(n_1078),
.B2(n_980),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1163),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1170),
.A2(n_1061),
.B1(n_1054),
.B2(n_1009),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1184),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1190),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1170),
.A2(n_1009),
.B1(n_1090),
.B2(n_1042),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1191),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1192),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1203),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1209),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1213),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1215),
.B(n_1128),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1161),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1213),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1214),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1208),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1195),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1195),
.A2(n_1189),
.B1(n_1042),
.B2(n_1030),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1151),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1159),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1196),
.A2(n_980),
.B1(n_1017),
.B2(n_1035),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1164),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1183),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1198),
.A2(n_980),
.B1(n_1017),
.B2(n_1037),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1188),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1198),
.A2(n_980),
.B1(n_1037),
.B2(n_1058),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1167),
.A2(n_980),
.B1(n_1058),
.B2(n_1037),
.Y(n_1283)
);

INVx6_ASAP7_75t_L g1284 ( 
.A(n_1159),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1209),
.A2(n_1024),
.B(n_1021),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1167),
.A2(n_980),
.B1(n_1005),
.B2(n_1018),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1167),
.B(n_1128),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1182),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1176),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1159),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1162),
.Y(n_1292)
);

BUFx2_ASAP7_75t_SL g1293 ( 
.A(n_1173),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1224),
.A2(n_1226),
.B1(n_1219),
.B2(n_1244),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1249),
.B(n_1036),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1267),
.B(n_1036),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1274),
.A2(n_980),
.B1(n_1167),
.B2(n_1051),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1227),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1220),
.Y(n_1299)
);

INVx5_ASAP7_75t_SL g1300 ( 
.A(n_1247),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1259),
.A2(n_990),
.B1(n_1110),
.B2(n_1109),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1274),
.A2(n_1167),
.B1(n_1051),
.B2(n_1018),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1259),
.A2(n_1018),
.B1(n_1020),
.B2(n_1011),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1246),
.A2(n_1018),
.B1(n_1020),
.B2(n_1011),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1278),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1270),
.B(n_986),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1249),
.B(n_986),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1230),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1262),
.A2(n_1020),
.B1(n_1029),
.B2(n_1011),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1222),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1262),
.A2(n_740),
.B(n_736),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1225),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1289),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1223),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1239),
.A2(n_1240),
.B1(n_1243),
.B2(n_1245),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1245),
.A2(n_1029),
.B1(n_1038),
.B2(n_1033),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1254),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1271),
.B(n_986),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1277),
.A2(n_1050),
.B1(n_1144),
.B2(n_1006),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1260),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1223),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_SL g1322 ( 
.A(n_1254),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1256),
.A2(n_1258),
.B1(n_1232),
.B2(n_1269),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1235),
.A2(n_1121),
.B1(n_754),
.B2(n_725),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1256),
.A2(n_1110),
.B1(n_716),
.B2(n_726),
.Y(n_1325)
);

BUFx4f_ASAP7_75t_SL g1326 ( 
.A(n_1242),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1248),
.A2(n_1029),
.B1(n_1038),
.B2(n_1033),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1290),
.A2(n_716),
.B1(n_726),
.B2(n_725),
.Y(n_1328)
);

OAI222xp33_ASAP7_75t_L g1329 ( 
.A1(n_1282),
.A2(n_1059),
.B1(n_1060),
.B2(n_1038),
.C1(n_1041),
.C2(n_1045),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1286),
.A2(n_1033),
.B1(n_1045),
.B2(n_1041),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1232),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1229),
.B(n_1173),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_SL g1333 ( 
.A1(n_1258),
.A2(n_1006),
.B1(n_1060),
.B2(n_1059),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1282),
.A2(n_1041),
.B1(n_1053),
.B2(n_1045),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1261),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1263),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1264),
.B(n_1146),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1228),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1257),
.A2(n_756),
.B(n_746),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1237),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1283),
.A2(n_1044),
.B1(n_993),
.B2(n_1053),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1280),
.A2(n_756),
.B1(n_762),
.B2(n_746),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1251),
.B(n_999),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1292),
.A2(n_762),
.B1(n_997),
.B2(n_1016),
.C(n_1013),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1238),
.A2(n_1044),
.B1(n_993),
.B2(n_1053),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1252),
.B(n_999),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1275),
.A2(n_1006),
.B(n_997),
.Y(n_1347)
);

OAI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1268),
.A2(n_984),
.B1(n_989),
.B2(n_993),
.C1(n_1010),
.C2(n_1111),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1250),
.B(n_1096),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1221),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1253),
.B(n_835),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1273),
.B(n_1019),
.C(n_1007),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1268),
.A2(n_999),
.B1(n_1019),
.B2(n_1010),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1293),
.A2(n_1144),
.B1(n_1181),
.B2(n_1180),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1272),
.A2(n_999),
.B1(n_1010),
.B2(n_989),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1253),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1265),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1281),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1231),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1287),
.A2(n_984),
.B1(n_1056),
.B2(n_761),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1233),
.A2(n_992),
.B(n_845),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1287),
.A2(n_1181),
.B1(n_1185),
.B2(n_1180),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1231),
.B(n_1209),
.Y(n_1363)
);

NOR2x1_ASAP7_75t_R g1364 ( 
.A(n_1266),
.B(n_1185),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1233),
.A2(n_1236),
.B1(n_1002),
.B2(n_1279),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1229),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1331),
.B(n_1229),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1295),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1298),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1325),
.A2(n_1002),
.B1(n_1236),
.B2(n_1183),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1294),
.A2(n_1153),
.B1(n_1168),
.B2(n_1158),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1294),
.A2(n_761),
.B1(n_759),
.B2(n_1056),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1318),
.B(n_1307),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1315),
.A2(n_1234),
.B1(n_1284),
.B2(n_1276),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1302),
.A2(n_761),
.B1(n_759),
.B2(n_1056),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1324),
.A2(n_1002),
.B1(n_1183),
.B2(n_992),
.Y(n_1376)
);

OAI222xp33_ASAP7_75t_L g1377 ( 
.A1(n_1323),
.A2(n_1063),
.B1(n_1096),
.B2(n_1102),
.C1(n_1109),
.C2(n_1013),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1297),
.A2(n_1302),
.B1(n_1304),
.B2(n_1301),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1310),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1297),
.A2(n_1039),
.B1(n_1102),
.B2(n_972),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1304),
.A2(n_1039),
.B1(n_972),
.B2(n_1115),
.Y(n_1381)
);

OAI221xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1311),
.A2(n_1016),
.B1(n_1063),
.B2(n_1021),
.C(n_1007),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1306),
.B(n_1241),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1319),
.A2(n_1276),
.B1(n_1284),
.B2(n_1234),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1301),
.A2(n_1039),
.B1(n_1136),
.B2(n_1125),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1340),
.A2(n_1039),
.B1(n_1148),
.B2(n_644),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1312),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1338),
.B(n_1241),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1366),
.B(n_1241),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1357),
.A2(n_1039),
.B1(n_644),
.B2(n_648),
.Y(n_1390)
);

AOI222xp33_ASAP7_75t_L g1391 ( 
.A1(n_1342),
.A2(n_672),
.B1(n_643),
.B2(n_644),
.C1(n_648),
.C2(n_654),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1308),
.A2(n_1039),
.B1(n_648),
.B2(n_654),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1303),
.A2(n_1288),
.B1(n_1079),
.B2(n_1108),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1352),
.A2(n_1183),
.B1(n_1288),
.B2(n_1158),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1320),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1337),
.A2(n_1344),
.B1(n_1333),
.B2(n_1336),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1328),
.A2(n_1183),
.B1(n_1168),
.B2(n_1169),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1361),
.A2(n_1169),
.B1(n_1291),
.B2(n_1255),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1335),
.B(n_1255),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1303),
.A2(n_1079),
.B1(n_1108),
.B2(n_1160),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1353),
.A2(n_643),
.B1(n_672),
.B2(n_654),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1353),
.A2(n_643),
.B1(n_672),
.B2(n_724),
.Y(n_1402)
);

AOI222xp33_ASAP7_75t_L g1403 ( 
.A1(n_1339),
.A2(n_724),
.B1(n_727),
.B2(n_730),
.C1(n_975),
.C2(n_976),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1358),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1327),
.A2(n_730),
.B1(n_727),
.B2(n_1008),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1296),
.B(n_1255),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1362),
.A2(n_1183),
.B1(n_1291),
.B2(n_730),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1327),
.A2(n_1062),
.B1(n_1065),
.B2(n_1103),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1330),
.A2(n_1062),
.B1(n_1065),
.B2(n_727),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1330),
.A2(n_1065),
.B1(n_1062),
.B2(n_1145),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1347),
.A2(n_1108),
.B1(n_1160),
.B2(n_1094),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1309),
.A2(n_1145),
.B1(n_1139),
.B2(n_1008),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1349),
.B(n_1317),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1351),
.A2(n_1291),
.B1(n_1188),
.B2(n_1216),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1354),
.A2(n_1057),
.B(n_1024),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1334),
.A2(n_1094),
.B1(n_1216),
.B2(n_1188),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1309),
.A2(n_1145),
.B1(n_1139),
.B2(n_1008),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1316),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1322),
.A2(n_1212),
.B1(n_1206),
.B2(n_1072),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1316),
.A2(n_639),
.B1(n_613),
.B2(n_678),
.C(n_652),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1322),
.A2(n_1212),
.B1(n_1206),
.B2(n_1266),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1326),
.A2(n_1216),
.B1(n_734),
.B2(n_737),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1326),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1334),
.A2(n_1355),
.B1(n_1360),
.B2(n_1345),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1355),
.A2(n_1003),
.B1(n_975),
.B2(n_976),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1341),
.A2(n_1210),
.B1(n_1057),
.B2(n_1285),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1356),
.A2(n_1210),
.B1(n_1285),
.B2(n_1218),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1365),
.A2(n_734),
.B1(n_713),
.B2(n_737),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1332),
.B(n_1177),
.Y(n_1430)
);

OAI222xp33_ASAP7_75t_L g1431 ( 
.A1(n_1360),
.A2(n_734),
.B1(n_713),
.B2(n_737),
.C1(n_1003),
.C2(n_613),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1300),
.A2(n_1210),
.B1(n_1218),
.B2(n_1201),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1329),
.A2(n_976),
.B1(n_975),
.B2(n_1210),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1314),
.A2(n_1003),
.B1(n_976),
.B2(n_401),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1332),
.B(n_1299),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1321),
.A2(n_1003),
.B1(n_401),
.B2(n_1026),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1350),
.B(n_1177),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1300),
.B(n_1177),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1305),
.A2(n_401),
.B1(n_1026),
.B2(n_1032),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1368),
.B(n_1300),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1372),
.A2(n_1026),
.B1(n_1032),
.B2(n_652),
.Y(n_1441)
);

OAI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1382),
.A2(n_678),
.B(n_639),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1398),
.A2(n_1348),
.B(n_1313),
.Y(n_1443)
);

NAND4xp25_ASAP7_75t_L g1444 ( 
.A(n_1376),
.B(n_62),
.C(n_63),
.D(n_64),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_1359),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1378),
.A2(n_636),
.B1(n_620),
.B2(n_618),
.C(n_631),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1416),
.B(n_1379),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1372),
.A2(n_1433),
.B1(n_1397),
.B2(n_1439),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1437),
.B(n_1359),
.C(n_1364),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1387),
.B(n_64),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1435),
.B(n_1363),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1395),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1388),
.A2(n_401),
.B(n_1363),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1371),
.A2(n_1032),
.B1(n_1120),
.B2(n_1200),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1373),
.B(n_1177),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1419),
.A2(n_1218),
.B1(n_1201),
.B2(n_1200),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1427),
.A2(n_1218),
.B1(n_1201),
.B2(n_1200),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1403),
.A2(n_67),
.B(n_68),
.Y(n_1458)
);

OAI21xp33_ASAP7_75t_L g1459 ( 
.A1(n_1406),
.A2(n_1396),
.B(n_1385),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1374),
.A2(n_1201),
.B1(n_1200),
.B2(n_1032),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_68),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1389),
.B(n_69),
.Y(n_1462)
);

NAND4xp25_ASAP7_75t_L g1463 ( 
.A(n_1439),
.B(n_1438),
.C(n_1367),
.D(n_1383),
.Y(n_1463)
);

OAI21xp33_ASAP7_75t_L g1464 ( 
.A1(n_1370),
.A2(n_1415),
.B(n_1394),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_70),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1404),
.B(n_71),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1425),
.A2(n_626),
.B1(n_615),
.B2(n_611),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1399),
.B(n_72),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1369),
.B(n_73),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_75),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1414),
.B(n_78),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1432),
.B(n_78),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1425),
.B(n_79),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1422),
.B(n_79),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1377),
.A2(n_1375),
.B1(n_1401),
.B2(n_1402),
.C(n_1384),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1411),
.B(n_80),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1375),
.B(n_81),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1393),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1391),
.B(n_615),
.C(n_611),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1407),
.B(n_618),
.Y(n_1480)
);

OAI21xp33_ASAP7_75t_L g1481 ( 
.A1(n_1423),
.A2(n_626),
.B(n_615),
.Y(n_1481)
);

NOR3xp33_ASAP7_75t_L g1482 ( 
.A(n_1417),
.B(n_636),
.C(n_620),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1400),
.A2(n_758),
.B1(n_752),
.B2(n_741),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1412),
.B(n_626),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1429),
.A2(n_631),
.B(n_83),
.Y(n_1485)
);

NOR3xp33_ASAP7_75t_L g1486 ( 
.A(n_1431),
.B(n_84),
.C(n_85),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1420),
.A2(n_631),
.B(n_95),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1386),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1380),
.B(n_96),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1418),
.B(n_97),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1401),
.B(n_98),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1436),
.B(n_752),
.C(n_741),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1410),
.B(n_102),
.Y(n_1493)
);

AND2x2_ASAP7_75t_SL g1494 ( 
.A(n_1402),
.B(n_103),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1436),
.A2(n_752),
.B1(n_741),
.B2(n_107),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1447),
.B(n_1434),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1445),
.B(n_1434),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1452),
.B(n_1405),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1405),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1451),
.B(n_1440),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1478),
.Y(n_1501)
);

NOR3xp33_ASAP7_75t_L g1502 ( 
.A(n_1444),
.B(n_1421),
.C(n_1390),
.Y(n_1502)
);

AND2x2_ASAP7_75t_SL g1503 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1392),
.C(n_1408),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1475),
.A2(n_1426),
.B1(n_1381),
.B2(n_121),
.Y(n_1505)
);

NOR3xp33_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1426),
.C(n_106),
.Y(n_1506)
);

AOI211xp5_ASAP7_75t_L g1507 ( 
.A1(n_1458),
.A2(n_104),
.B(n_122),
.C(n_128),
.Y(n_1507)
);

NOR3xp33_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_135),
.C(n_136),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1453),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1476),
.B(n_140),
.C(n_145),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1449),
.B(n_148),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1462),
.B(n_150),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1465),
.B(n_154),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1457),
.B(n_157),
.Y(n_1514)
);

NOR3xp33_ASAP7_75t_SL g1515 ( 
.A(n_1461),
.B(n_158),
.C(n_160),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1468),
.B(n_161),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1448),
.A2(n_162),
.B1(n_163),
.B2(n_167),
.Y(n_1517)
);

NAND4xp75_ASAP7_75t_L g1518 ( 
.A(n_1443),
.B(n_1494),
.C(n_1475),
.D(n_1472),
.Y(n_1518)
);

OAI31xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1459),
.A2(n_169),
.A3(n_170),
.B(n_172),
.Y(n_1519)
);

AO21x2_ASAP7_75t_L g1520 ( 
.A1(n_1469),
.A2(n_174),
.B(n_177),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1453),
.B(n_179),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1450),
.B(n_181),
.Y(n_1522)
);

OA211x2_ASAP7_75t_L g1523 ( 
.A1(n_1474),
.A2(n_185),
.B(n_186),
.C(n_187),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1463),
.B(n_188),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1471),
.A2(n_189),
.B(n_191),
.C(n_194),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1466),
.B(n_195),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

NAND4xp75_ASAP7_75t_L g1529 ( 
.A(n_1446),
.B(n_197),
.C(n_198),
.D(n_199),
.Y(n_1529)
);

NAND4xp25_ASAP7_75t_L g1530 ( 
.A(n_1477),
.B(n_200),
.C(n_206),
.D(n_207),
.Y(n_1530)
);

NOR4xp75_ASAP7_75t_L g1531 ( 
.A(n_1442),
.B(n_210),
.C(n_211),
.D(n_212),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_213),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1457),
.B(n_215),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1456),
.B(n_216),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1482),
.B(n_220),
.C(n_221),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1496),
.B(n_1456),
.Y(n_1537)
);

XNOR2x2_ASAP7_75t_L g1538 ( 
.A(n_1518),
.B(n_1446),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1527),
.Y(n_1539)
);

XNOR2xp5_ASAP7_75t_L g1540 ( 
.A(n_1512),
.B(n_1460),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1509),
.Y(n_1541)
);

XNOR2xp5_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1542)
);

XNOR2xp5_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1486),
.Y(n_1543)
);

XOR2x1_ASAP7_75t_L g1544 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1454),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1528),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1506),
.A2(n_1486),
.B1(n_1483),
.B2(n_1493),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1495),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1527),
.B(n_1482),
.Y(n_1550)
);

BUFx4f_ASAP7_75t_L g1551 ( 
.A(n_1534),
.Y(n_1551)
);

XOR2x2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.B(n_1491),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1481),
.C(n_1480),
.Y(n_1553)
);

NAND4xp75_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1483),
.C(n_1479),
.D(n_1467),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1516),
.B(n_1441),
.Y(n_1556)
);

NAND4xp75_ASAP7_75t_L g1557 ( 
.A(n_1503),
.B(n_1492),
.C(n_225),
.D(n_227),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1521),
.Y(n_1558)
);

NAND4xp75_ASAP7_75t_L g1559 ( 
.A(n_1503),
.B(n_222),
.C(n_228),
.D(n_230),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1516),
.B(n_231),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1524),
.B(n_233),
.C(n_234),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1528),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1522),
.B(n_238),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1496),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1547),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1562),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1539),
.B(n_1499),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1539),
.B(n_1521),
.Y(n_1568)
);

AO22x1_ASAP7_75t_L g1569 ( 
.A1(n_1537),
.A2(n_1534),
.B1(n_1532),
.B2(n_1533),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1539),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1541),
.Y(n_1571)
);

XNOR2x2_ASAP7_75t_L g1572 ( 
.A(n_1538),
.B(n_1514),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1551),
.A2(n_1505),
.B1(n_1514),
.B2(n_1510),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_R g1576 ( 
.A(n_1551),
.B(n_1526),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1555),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1558),
.Y(n_1579)
);

XOR2x2_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1580)
);

XOR2x2_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1549),
.Y(n_1582)
);

XNOR2xp5_ASAP7_75t_L g1583 ( 
.A(n_1540),
.B(n_1515),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

XOR2x2_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1531),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1581),
.A2(n_1545),
.B1(n_1549),
.B2(n_1552),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1567),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1582),
.A2(n_1551),
.B1(n_1545),
.B2(n_1548),
.Y(n_1588)
);

OA22x2_ASAP7_75t_L g1589 ( 
.A1(n_1572),
.A2(n_1546),
.B1(n_1560),
.B2(n_1550),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1584),
.Y(n_1590)
);

AO22x2_ASAP7_75t_L g1591 ( 
.A1(n_1572),
.A2(n_1544),
.B1(n_1559),
.B2(n_1557),
.Y(n_1591)
);

OA22x2_ASAP7_75t_L g1592 ( 
.A1(n_1583),
.A2(n_1581),
.B1(n_1573),
.B2(n_1564),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1575),
.Y(n_1593)
);

OA22x2_ASAP7_75t_L g1594 ( 
.A1(n_1564),
.A2(n_1544),
.B1(n_1556),
.B2(n_1517),
.Y(n_1594)
);

OAI22x1_ASAP7_75t_L g1595 ( 
.A1(n_1579),
.A2(n_1532),
.B1(n_1563),
.B2(n_1504),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1568),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1576),
.Y(n_1598)
);

OA22x2_ASAP7_75t_L g1599 ( 
.A1(n_1579),
.A2(n_1519),
.B1(n_1561),
.B2(n_1530),
.Y(n_1599)
);

OA22x2_ASAP7_75t_L g1600 ( 
.A1(n_1585),
.A2(n_1580),
.B1(n_1575),
.B2(n_1569),
.Y(n_1600)
);

OA22x2_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1553),
.B1(n_1563),
.B2(n_1554),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1566),
.B(n_1570),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1508),
.B1(n_1535),
.B2(n_1498),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1580),
.A2(n_1520),
.B1(n_1525),
.B2(n_1502),
.Y(n_1604)
);

AO22x2_ASAP7_75t_L g1605 ( 
.A1(n_1571),
.A2(n_1529),
.B1(n_1520),
.B2(n_242),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_SL g1607 ( 
.A(n_1588),
.B(n_1577),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1597),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1598),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1593),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1601),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1587),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1602),
.Y(n_1613)
);

XNOR2xp5_ASAP7_75t_L g1614 ( 
.A(n_1589),
.B(n_1578),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1595),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1604),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1608),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1609),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_SL g1620 ( 
.A(n_1616),
.Y(n_1620)
);

AOI22x1_ASAP7_75t_L g1621 ( 
.A1(n_1609),
.A2(n_1591),
.B1(n_1605),
.B2(n_1596),
.Y(n_1621)
);

AOI31xp33_ASAP7_75t_L g1622 ( 
.A1(n_1611),
.A2(n_1603),
.A3(n_1600),
.B(n_1592),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1606),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1610),
.Y(n_1624)
);

OA22x2_ASAP7_75t_L g1625 ( 
.A1(n_1611),
.A2(n_1594),
.B1(n_1591),
.B2(n_1599),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1617),
.A2(n_1605),
.B(n_1574),
.C(n_248),
.Y(n_1626)
);

NAND4xp25_ASAP7_75t_SL g1627 ( 
.A(n_1612),
.B(n_1574),
.C(n_241),
.D(n_251),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1619),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1625),
.A2(n_1614),
.B1(n_1615),
.B2(n_1613),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1623),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1622),
.A2(n_1607),
.B(n_252),
.C(n_255),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1625),
.A2(n_239),
.B1(n_259),
.B2(n_260),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1618),
.Y(n_1634)
);

AO22x2_ASAP7_75t_L g1635 ( 
.A1(n_1624),
.A2(n_366),
.B1(n_270),
.B2(n_274),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1621),
.A2(n_262),
.B1(n_275),
.B2(n_277),
.C(n_278),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1629),
.A2(n_1626),
.B1(n_1627),
.B2(n_283),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1628),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1632),
.A2(n_1636),
.B1(n_1635),
.B2(n_1633),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1630),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1634),
.Y(n_1641)
);

AO22x2_ASAP7_75t_L g1642 ( 
.A1(n_1631),
.A2(n_281),
.B1(n_282),
.B2(n_286),
.Y(n_1642)
);

AO22x1_ASAP7_75t_L g1643 ( 
.A1(n_1633),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1638),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1640),
.B(n_1641),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1637),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1643),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1642),
.A2(n_293),
.B1(n_297),
.B2(n_298),
.Y(n_1648)
);

AO22x2_ASAP7_75t_L g1649 ( 
.A1(n_1644),
.A2(n_1639),
.B1(n_303),
.B2(n_306),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1645),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1647),
.A2(n_302),
.B1(n_307),
.B2(n_309),
.Y(n_1651)
);

AND4x1_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_310),
.C(n_312),
.D(n_313),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1650),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1649),
.B(n_1648),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1651),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1652),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1654),
.Y(n_1658)
);

AO22x2_ASAP7_75t_L g1659 ( 
.A1(n_1656),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1655),
.A2(n_321),
.B1(n_322),
.B2(n_326),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1657),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1658),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1659),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1660),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1657),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1663),
.A2(n_327),
.B1(n_328),
.B2(n_330),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1662),
.A2(n_1665),
.B1(n_1661),
.B2(n_1663),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1664),
.A2(n_364),
.B1(n_337),
.B2(n_338),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1667),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1666),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1667),
.Y(n_1672)
);

AO22x2_ASAP7_75t_L g1673 ( 
.A1(n_1669),
.A2(n_1672),
.B1(n_1670),
.B2(n_1671),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1671),
.A2(n_336),
.B1(n_340),
.B2(n_341),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1671),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1673),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1674),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1675),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1676),
.A2(n_1678),
.B1(n_1677),
.B2(n_353),
.C(n_355),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_350),
.B(n_351),
.C(n_357),
.Y(n_1680)
);


endmodule