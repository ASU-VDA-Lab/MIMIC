module fake_ariane_41_n_2113 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2113);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2113;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_103),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_9),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_139),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_108),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_43),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_148),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_64),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_66),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_184),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_138),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_162),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_56),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_55),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_28),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_177),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_137),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_59),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_110),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_115),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_77),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_89),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_28),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_42),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_120),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_29),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_145),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_32),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_205),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_31),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_50),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_82),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_102),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_119),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_122),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_86),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_77),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_62),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_203),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_23),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_66),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_49),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_50),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_61),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_15),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_99),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_192),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_92),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_107),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_56),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_166),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_84),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_59),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_111),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_45),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_35),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_63),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_149),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_173),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_94),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_193),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_88),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_197),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_155),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_95),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_2),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_74),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_22),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_131),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_45),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_35),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_143),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_141),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_160),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_109),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_81),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_38),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_52),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_20),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_150),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_48),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_27),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_179),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_144),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_76),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_60),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_128),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_187),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_71),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_136),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_14),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_78),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_74),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_64),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_20),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_133),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_16),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_134),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_161),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_101),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_146),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_105),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_48),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_62),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_182),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_135),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_65),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_121),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_72),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_5),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_126),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_54),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_60),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_4),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_25),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_72),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_44),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_79),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_21),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_0),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_71),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_10),
.Y(n_364)
);

BUFx8_ASAP7_75t_SL g365 ( 
.A(n_152),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_151),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_21),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_70),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_90),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_51),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_183),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_33),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_19),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_53),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_6),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_31),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_18),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_17),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_96),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_65),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_116),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_69),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_3),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_1),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_33),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_93),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_13),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_114),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_68),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_7),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_178),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_38),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_204),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_26),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_186),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_46),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_185),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_168),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_12),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_164),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_37),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_165),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_100),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_210),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_210),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_217),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_217),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_218),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_276),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_218),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_365),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_229),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_229),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_380),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_306),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_238),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_382),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_215),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_244),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_223),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_244),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_242),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_266),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_224),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_249),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_306),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_242),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_249),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_252),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_283),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_221),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_344),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_344),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_252),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_296),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_323),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_221),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_253),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_253),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_259),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_211),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_301),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_259),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_260),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_322),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_260),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_261),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_261),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_211),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_322),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_265),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_265),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_336),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_285),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_324),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_285),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_332),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_289),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_333),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_231),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_241),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_289),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_298),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_221),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_298),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_305),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_208),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_305),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_336),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_312),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_312),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_315),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_364),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_400),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_364),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_207),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_209),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_315),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_219),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_232),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_328),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_328),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_330),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_248),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_222),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_233),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_392),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_227),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_330),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_337),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_236),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_337),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_221),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_227),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_354),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_359),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_243),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_245),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_341),
.Y(n_505)
);

INVxp33_ASAP7_75t_SL g506 ( 
.A(n_258),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_264),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_270),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_272),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_341),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_391),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_273),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_274),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_216),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_483),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_414),
.B(n_251),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_406),
.B(n_216),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_422),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

OR2x2_ASAP7_75t_SL g524 ( 
.A(n_465),
.B(n_319),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_421),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_428),
.A2(n_438),
.B1(n_432),
.B2(n_437),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_406),
.B(n_291),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_425),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_R g531 ( 
.A(n_413),
.B(n_360),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_407),
.B(n_291),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_469),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_499),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_429),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_481),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_491),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_435),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_446),
.B(n_404),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_447),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_408),
.B(n_308),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_441),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_408),
.B(n_308),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_437),
.A2(n_345),
.B1(n_334),
.B2(n_237),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_441),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_462),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_409),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_410),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_464),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_410),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_492),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_412),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_412),
.B(n_319),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_486),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_415),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_415),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_416),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_478),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_416),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_419),
.B(n_347),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_490),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_497),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_454),
.B(n_317),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_423),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_423),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_440),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_424),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_506),
.B(n_302),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_424),
.B(n_347),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_426),
.B(n_371),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_480),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_430),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_430),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_433),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_501),
.Y(n_590)
);

NAND2x1_ASAP7_75t_L g591 ( 
.A(n_433),
.B(n_220),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_434),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_502),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_439),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_507),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_511),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_439),
.B(n_371),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_525),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_529),
.A2(n_427),
.B1(n_494),
.B2(n_444),
.Y(n_601)
);

OA22x2_ASAP7_75t_L g602 ( 
.A1(n_529),
.A2(n_482),
.B1(n_431),
.B2(n_450),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_587),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_587),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_591),
.A2(n_444),
.B(n_443),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_527),
.B(n_466),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_575),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_527),
.B(n_418),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_539),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_516),
.B(n_513),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_529),
.A2(n_443),
.B1(n_448),
.B2(n_445),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_529),
.B(n_445),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_587),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_592),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_546),
.B(n_448),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_592),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_592),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_592),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_592),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_581),
.B(n_508),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_572),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_566),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_566),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_514),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_552),
.A2(n_279),
.B1(n_284),
.B2(n_278),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_520),
.A2(n_509),
.B1(n_500),
.B2(n_295),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_546),
.B(n_449),
.Y(n_637)
);

AO22x2_ASAP7_75t_L g638 ( 
.A1(n_552),
.A2(n_575),
.B1(n_521),
.B2(n_535),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_550),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_SL g640 ( 
.A1(n_521),
.A2(n_451),
.B(n_449),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_596),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_517),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_517),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_523),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_545),
.B(n_553),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_523),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_520),
.A2(n_304),
.B1(n_307),
.B2(n_290),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_550),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_549),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_576),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_598),
.B(n_417),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_534),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_545),
.B(n_451),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g657 ( 
.A1(n_572),
.A2(n_397),
.B(n_389),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_519),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_553),
.B(n_452),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_420),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_562),
.B(n_452),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_569),
.B(n_458),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_577),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_536),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_564),
.B(n_493),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_534),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_557),
.B(n_456),
.C(n_453),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

INVxp33_ASAP7_75t_SL g672 ( 
.A(n_530),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_577),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_580),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_537),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_580),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_549),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_549),
.A2(n_453),
.B1(n_457),
.B2(n_456),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_564),
.B(n_457),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_557),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_580),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_596),
.B(n_459),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_541),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_589),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_531),
.B(n_459),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_564),
.B(n_461),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_535),
.A2(n_311),
.B1(n_321),
.B2(n_310),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_411),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_589),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_559),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_536),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_591),
.A2(n_463),
.B(n_461),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_559),
.B(n_463),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_561),
.B(n_467),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_542),
.B(n_467),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_538),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_536),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_536),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_561),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_563),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_563),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_586),
.B(n_468),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_567),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_522),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_522),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_586),
.B(n_568),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_518),
.B(n_468),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

CKINVDCx8_ASAP7_75t_R g713 ( 
.A(n_579),
.Y(n_713)
);

OAI21xp33_ASAP7_75t_SL g714 ( 
.A1(n_582),
.A2(n_471),
.B(n_470),
.Y(n_714)
);

INVx5_ASAP7_75t_L g715 ( 
.A(n_522),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_526),
.B(n_540),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_564),
.B(n_549),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_528),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_548),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_571),
.B(n_470),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_528),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_574),
.A2(n_578),
.B1(n_585),
.B2(n_524),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_556),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_583),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_528),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_532),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_551),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_532),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_551),
.B(n_471),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_588),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_532),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_560),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_588),
.Y(n_736)
);

AND3x1_ASAP7_75t_L g737 ( 
.A(n_582),
.B(n_237),
.C(n_230),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_593),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_593),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_533),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_551),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_533),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_533),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_595),
.B(n_473),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_595),
.B(n_473),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_544),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_584),
.B(n_599),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_584),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_599),
.B(n_475),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_524),
.B(n_475),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_544),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_544),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_747),
.B(n_389),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_638),
.A2(n_477),
.B1(n_484),
.B2(n_476),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_614),
.A2(n_476),
.B1(n_484),
.B2(n_477),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_612),
.B(n_460),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_748),
.B(n_487),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_603),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_747),
.B(n_397),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_748),
.B(n_487),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_685),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_747),
.B(n_488),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_747),
.B(n_488),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_636),
.B(n_405),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_685),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_603),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_681),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_636),
.B(n_405),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_625),
.B(n_489),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_681),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_692),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_624),
.B(n_489),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_636),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_658),
.B(n_479),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_638),
.A2(n_496),
.B1(n_498),
.B2(n_495),
.Y(n_776)
);

BUFx5_ASAP7_75t_L g777 ( 
.A(n_692),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_609),
.B(n_565),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_652),
.B(n_495),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_652),
.B(n_677),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_642),
.B(n_246),
.C(n_230),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_691),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_691),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_677),
.B(n_496),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_730),
.B(n_498),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_692),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_725),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_628),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_636),
.B(n_505),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_741),
.B(n_505),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_730),
.B(n_510),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_725),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_741),
.B(n_510),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_725),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_603),
.B(n_221),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_741),
.B(n_220),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_628),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_733),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_710),
.B(n_313),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_614),
.A2(n_316),
.B1(n_234),
.B2(n_269),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_733),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_608),
.B(n_573),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_618),
.B(n_339),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_714),
.A2(n_329),
.B(n_318),
.C(n_246),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_642),
.B(n_455),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_741),
.B(n_234),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_638),
.A2(n_251),
.B1(n_381),
.B2(n_317),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_628),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_673),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_673),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_733),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_637),
.B(n_390),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_750),
.B(n_390),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_706),
.B(n_269),
.Y(n_815)
);

BUFx8_ASAP7_75t_L g816 ( 
.A(n_607),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_601),
.B(n_597),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_706),
.B(n_316),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_706),
.B(n_228),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_673),
.B(n_228),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_SL g821 ( 
.A1(n_632),
.A2(n_594),
.B1(n_590),
.B2(n_403),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_660),
.B(n_267),
.C(n_250),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_702),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_654),
.B(n_267),
.C(n_250),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_638),
.A2(n_251),
.B1(n_381),
.B2(n_326),
.Y(n_825)
);

AO221x1_ASAP7_75t_L g826 ( 
.A1(n_650),
.A2(n_254),
.B1(n_287),
.B2(n_385),
.C(n_292),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_614),
.A2(n_732),
.B1(n_640),
.B2(n_661),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_702),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_673),
.B(n_281),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_602),
.A2(n_251),
.B1(n_381),
.B2(n_326),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_749),
.B(n_268),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_673),
.B(n_281),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_732),
.B(n_268),
.Y(n_833)
);

NOR2x2_ASAP7_75t_L g834 ( 
.A(n_614),
.B(n_317),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_714),
.A2(n_554),
.B(n_547),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_735),
.B(n_275),
.C(n_271),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_600),
.B(n_206),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_603),
.B(n_366),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_626),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_602),
.A2(n_381),
.B1(n_317),
.B2(n_326),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_737),
.B(n_366),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_617),
.B(n_402),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_626),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_630),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_617),
.B(n_402),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_600),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_614),
.A2(n_256),
.B1(n_282),
.B2(n_399),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_617),
.B(n_323),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_602),
.A2(n_326),
.B1(n_254),
.B2(n_314),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_630),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_610),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_641),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_703),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_609),
.B(n_271),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_672),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_275),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_664),
.B(n_277),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_690),
.Y(n_858)
);

INVx8_ASAP7_75t_L g859 ( 
.A(n_679),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_698),
.B(n_212),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_641),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_657),
.A2(n_254),
.B1(n_314),
.B2(n_262),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_668),
.B(n_277),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_703),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_617),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_698),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_704),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_704),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_617),
.B(n_323),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_SL g870 ( 
.A(n_720),
.B(n_287),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_623),
.B(n_254),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_721),
.B(n_292),
.Y(n_872)
);

NOR2x1p5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_325),
.Y(n_873)
);

NAND2x1_ASAP7_75t_L g874 ( 
.A(n_627),
.B(n_547),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_607),
.B(n_293),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_613),
.B(n_293),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_708),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_632),
.B(n_335),
.C(n_331),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_679),
.B(n_294),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_690),
.B(n_294),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_717),
.B(n_318),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_688),
.B(n_329),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_688),
.B(n_350),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_683),
.B(n_338),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_657),
.A2(n_262),
.B1(n_361),
.B2(n_357),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_623),
.B(n_323),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_623),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_717),
.B(n_350),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_SL g890 ( 
.A(n_724),
.B(n_357),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_643),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_643),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_678),
.B(n_361),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_640),
.A2(n_213),
.B1(n_214),
.B2(n_225),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_351),
.C(n_348),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_668),
.B(n_368),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_727),
.B(n_353),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_712),
.B(n_368),
.Y(n_898)
);

O2A1O1Ixp5_ASAP7_75t_L g899 ( 
.A1(n_606),
.A2(n_383),
.B(n_387),
.C(n_385),
.Y(n_899)
);

OR2x2_ASAP7_75t_SL g900 ( 
.A(n_713),
.B(n_633),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_687),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_623),
.B(n_379),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_623),
.B(n_379),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_718),
.B(n_383),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_718),
.B(n_384),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_711),
.A2(n_226),
.B1(n_235),
.B2(n_239),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_723),
.A2(n_240),
.B1(n_247),
.B2(n_255),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_728),
.A2(n_387),
.B(n_384),
.C(n_388),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_728),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_716),
.B(n_388),
.C(n_355),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_646),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_646),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_697),
.B(n_358),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_736),
.B(n_362),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_738),
.B(n_739),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_738),
.B(n_363),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_705),
.B(n_367),
.C(n_370),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_653),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_648),
.A2(n_555),
.B(n_554),
.C(n_547),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_656),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_778),
.B(n_689),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_773),
.B(n_659),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_799),
.B(n_695),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_823),
.Y(n_924)
);

AND3x1_ASAP7_75t_L g925 ( 
.A(n_756),
.B(n_713),
.C(n_696),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_777),
.B(n_619),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_828),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_855),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_761),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_858),
.B(n_744),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_803),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_915),
.A2(n_745),
.B1(n_619),
.B2(n_670),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_846),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_920),
.B(n_653),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_882),
.B(n_670),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_864),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_895),
.B(n_373),
.C(n_372),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_775),
.A2(n_737),
.B1(n_619),
.B2(n_662),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_867),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_SL g941 ( 
.A(n_870),
.B(n_375),
.C(n_374),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_841),
.A2(n_662),
.B1(n_676),
.B2(n_663),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_757),
.B(n_663),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_868),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_806),
.B(n_657),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_758),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_854),
.B(n_665),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_866),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_760),
.B(n_665),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_816),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_606),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_762),
.B(n_763),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_865),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_899),
.A2(n_674),
.B(n_667),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_804),
.B(n_667),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_856),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_761),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_877),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_880),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_859),
.B(n_627),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_769),
.B(n_674),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_814),
.B(n_676),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_841),
.A2(n_682),
.B1(n_686),
.B2(n_629),
.Y(n_963)
);

AND2x6_ASAP7_75t_SL g964 ( 
.A(n_885),
.B(n_682),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_882),
.B(n_889),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_857),
.B(n_686),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_777),
.B(n_616),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_765),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_765),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_909),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_859),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_777),
.B(n_616),
.Y(n_972)
);

INVx6_ASAP7_75t_L g973 ( 
.A(n_816),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_758),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_839),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_839),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_873),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_859),
.A2(n_615),
.B1(n_604),
.B2(n_620),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_782),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_788),
.A2(n_605),
.B(n_604),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_843),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_863),
.B(n_629),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_843),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_774),
.B(n_631),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_889),
.B(n_694),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_SL g986 ( 
.A(n_870),
.B(n_377),
.C(n_376),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_844),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_851),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_859),
.B(n_900),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_779),
.B(n_631),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_784),
.B(n_785),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_821),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_782),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_758),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_817),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_791),
.B(n_634),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_753),
.B(n_634),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_826),
.A2(n_669),
.B1(n_635),
.B2(n_644),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_889),
.B(n_694),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_881),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_SL g1001 ( 
.A1(n_878),
.A2(n_378),
.B1(n_394),
.B2(n_396),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_808),
.A2(n_825),
.B1(n_759),
.B2(n_753),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_901),
.B(n_627),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_783),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_759),
.B(n_635),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_897),
.B(n_644),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_813),
.B(n_645),
.Y(n_1007)
);

INVx8_ASAP7_75t_L g1008 ( 
.A(n_758),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_844),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_837),
.B(n_666),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_886),
.A2(n_675),
.B1(n_684),
.B2(n_645),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_875),
.B(n_647),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_777),
.B(n_621),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_850),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_834),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_850),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_783),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_888),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_827),
.B(n_647),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_896),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_754),
.B(n_649),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_890),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_852),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_852),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_776),
.B(n_649),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_777),
.B(n_621),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_861),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_824),
.B(n_401),
.C(n_398),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_861),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_865),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_888),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_888),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_891),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_892),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_892),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_789),
.B(n_627),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_780),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_888),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_788),
.A2(n_605),
.B1(n_611),
.B2(n_615),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_777),
.B(n_611),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_777),
.B(n_620),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_755),
.B(n_622),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_911),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_879),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_911),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_912),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_912),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_822),
.B(n_781),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_918),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_883),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_865),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_833),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_789),
.B(n_655),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_797),
.B(n_622),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_797),
.B(n_651),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_913),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_810),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_918),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_872),
.B(n_655),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_831),
.B(n_669),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_800),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_790),
.A2(n_651),
.B(n_639),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_884),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_898),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_849),
.A2(n_671),
.B1(n_684),
.B2(n_680),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_904),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_SL g1068 ( 
.A(n_764),
.B(n_651),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_800),
.A2(n_809),
.B1(n_772),
.B2(n_786),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_862),
.A2(n_671),
.B1(n_675),
.B2(n_680),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_764),
.B(n_651),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_810),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_834),
.Y(n_1073)
);

INVx2_ASAP7_75t_SL g1074 ( 
.A(n_876),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_790),
.A2(n_639),
.B(n_701),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_809),
.B(n_693),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_893),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_840),
.A2(n_701),
.B1(n_699),
.B2(n_693),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_905),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_767),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_770),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_860),
.B(n_639),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_811),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_836),
.B(n_699),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_914),
.B(n_707),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_830),
.A2(n_729),
.B1(n_751),
.B2(n_746),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_907),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_894),
.A2(n_729),
.B1(n_751),
.B2(n_746),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_771),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_811),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_916),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_768),
.B(n_707),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_787),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_792),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_794),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_798),
.B(n_666),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_802),
.B(n_722),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_812),
.A2(n_666),
.B1(n_726),
.B2(n_742),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_793),
.A2(n_666),
.B1(n_752),
.B2(n_743),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_874),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_793),
.A2(n_666),
.B1(n_752),
.B2(n_743),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_835),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_819),
.A2(n_919),
.B(n_818),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_917),
.B(n_743),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_766),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_819),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_801),
.B(n_722),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_910),
.B(n_666),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_930),
.B(n_847),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_971),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_922),
.A2(n_796),
.B1(n_807),
.B2(n_805),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_952),
.A2(n_796),
.B1(n_807),
.B2(n_805),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_961),
.A2(n_818),
.B(n_815),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_991),
.A2(n_923),
.B(n_943),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_931),
.B(n_906),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1028),
.B(n_908),
.C(n_815),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_924),
.Y(n_1117)
);

OAI22x1_ASAP7_75t_L g1118 ( 
.A1(n_1087),
.A2(n_838),
.B1(n_842),
.B2(n_845),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_930),
.B(n_908),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1000),
.B(n_726),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1037),
.A2(n_829),
.B(n_820),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_949),
.A2(n_832),
.B(n_838),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_971),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_927),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1049),
.A2(n_842),
.B(n_845),
.C(n_887),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1091),
.A2(n_795),
.B(n_871),
.C(n_887),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_960),
.A2(n_731),
.B1(n_734),
.B2(n_740),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_936),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_967),
.A2(n_903),
.B(n_902),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1008),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_967),
.A2(n_903),
.B(n_902),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_960),
.A2(n_742),
.B1(n_734),
.B2(n_740),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1012),
.B(n_731),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1071),
.A2(n_869),
.B(n_848),
.C(n_752),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1053),
.A2(n_869),
.B(n_848),
.C(n_558),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1064),
.A2(n_554),
.B(n_555),
.C(n_558),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_965),
.A2(n_752),
.B1(n_343),
.B2(n_342),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_921),
.B(n_263),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1002),
.A2(n_346),
.B1(n_286),
.B2(n_288),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_956),
.B(n_0),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_1008),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1008),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_937),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_972),
.A2(n_719),
.B(n_715),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1002),
.A2(n_940),
.B1(n_958),
.B2(n_944),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_959),
.A2(n_349),
.B1(n_297),
.B2(n_299),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_973),
.B(n_379),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1071),
.A2(n_719),
.B(n_715),
.C(n_709),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_948),
.B(n_709),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1020),
.B(n_709),
.Y(n_1150)
);

AND2x6_ASAP7_75t_L g1151 ( 
.A(n_951),
.B(n_379),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1045),
.B(n_709),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_933),
.B(n_280),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_988),
.B(n_300),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1057),
.B(n_303),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_946),
.Y(n_1156)
);

OAI21xp33_ASAP7_75t_L g1157 ( 
.A1(n_941),
.A2(n_309),
.B(n_320),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1023),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_970),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1051),
.B(n_947),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_972),
.A2(n_719),
.B(n_715),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1037),
.A2(n_719),
.B(n_715),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1013),
.A2(n_719),
.B(n_715),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1013),
.A2(n_719),
.B(n_715),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_1042),
.B(n_1041),
.Y(n_1165)
);

AOI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1074),
.A2(n_709),
.B(n_327),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_928),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1022),
.A2(n_1103),
.B(n_1104),
.C(n_954),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_946),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1065),
.B(n_4),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_973),
.B(n_340),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_950),
.B(n_379),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1023),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_946),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_994),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1026),
.A2(n_386),
.B(n_356),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1102),
.A2(n_395),
.B1(n_393),
.B2(n_369),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1006),
.A2(n_352),
.B1(n_558),
.B2(n_555),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1027),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1057),
.B(n_6),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_953),
.B(n_80),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1052),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_995),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1067),
.B(n_7),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1079),
.A2(n_1003),
.B(n_939),
.C(n_989),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1041),
.A2(n_202),
.B(n_201),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1001),
.B(n_8),
.C(n_10),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_989),
.B(n_964),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_L g1189 ( 
.A(n_977),
.B(n_8),
.C(n_11),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_945),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_925),
.Y(n_1191)
);

OAI33xp33_ASAP7_75t_L g1192 ( 
.A1(n_934),
.A2(n_17),
.A3(n_18),
.B1(n_22),
.B2(n_23),
.B3(n_24),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_R g1193 ( 
.A(n_992),
.B(n_199),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1042),
.A2(n_195),
.B(n_194),
.Y(n_1194)
);

AO32x1_ASAP7_75t_L g1195 ( 
.A1(n_1069),
.A2(n_24),
.A3(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_935),
.B(n_30),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_935),
.A2(n_982),
.B1(n_963),
.B2(n_978),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_926),
.A2(n_191),
.B(n_181),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_926),
.A2(n_167),
.B(n_158),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1015),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_966),
.A2(n_1056),
.B(n_996),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1019),
.A2(n_1007),
.B(n_962),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_941),
.A2(n_30),
.B(n_34),
.C(n_36),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1073),
.B(n_37),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1038),
.B(n_39),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_994),
.B(n_41),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_994),
.B(n_83),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_955),
.A2(n_85),
.B(n_153),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1077),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_963),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1052),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1038),
.B(n_47),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1084),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_951),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1027),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_986),
.B(n_54),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1061),
.B(n_55),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1060),
.B(n_57),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1003),
.B(n_57),
.Y(n_1219)
);

O2A1O1Ixp5_ASAP7_75t_L g1220 ( 
.A1(n_1043),
.A2(n_58),
.B(n_61),
.C(n_63),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_986),
.B(n_58),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_975),
.B(n_67),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1104),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1080),
.B(n_70),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1052),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1056),
.A2(n_117),
.B(n_147),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_994),
.B(n_73),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_990),
.A2(n_113),
.B(n_142),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1075),
.A2(n_112),
.B(n_130),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1063),
.A2(n_106),
.B(n_129),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_976),
.B(n_73),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_942),
.A2(n_75),
.B(n_76),
.C(n_87),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_SL g1233 ( 
.A(n_938),
.B(n_75),
.C(n_91),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_938),
.Y(n_1234)
);

BUFx4f_ASAP7_75t_L g1235 ( 
.A(n_1082),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_980),
.A2(n_1054),
.B(n_932),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_985),
.A2(n_97),
.B1(n_98),
.B2(n_118),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1055),
.A2(n_1068),
.B(n_1043),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_981),
.B(n_123),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1052),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1039),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_983),
.B(n_987),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1055),
.A2(n_984),
.B(n_985),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_R g1244 ( 
.A(n_1039),
.B(n_124),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_999),
.A2(n_127),
.B(n_156),
.C(n_1085),
.Y(n_1245)
);

NOR2xp67_ASAP7_75t_L g1246 ( 
.A(n_1082),
.B(n_1039),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1009),
.B(n_1014),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_999),
.A2(n_1040),
.B(n_1100),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1016),
.B(n_1046),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1081),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1089),
.Y(n_1251)
);

AO22x1_ASAP7_75t_L g1252 ( 
.A1(n_1108),
.A2(n_1093),
.B1(n_1095),
.B2(n_1094),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1024),
.B(n_1036),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1106),
.A2(n_1048),
.B(n_1044),
.C(n_1059),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1021),
.A2(n_1025),
.B1(n_1034),
.B2(n_1050),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1039),
.B(n_974),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_946),
.Y(n_1257)
);

AO32x2_ASAP7_75t_L g1258 ( 
.A1(n_1098),
.A2(n_1105),
.A3(n_1032),
.B1(n_998),
.B2(n_1066),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1058),
.B(n_1072),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_974),
.B(n_1018),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1058),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1029),
.A2(n_1035),
.B1(n_1047),
.B2(n_1033),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1100),
.A2(n_1062),
.B(n_1092),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1029),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1033),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_997),
.A2(n_1005),
.B1(n_1047),
.B2(n_1035),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_929),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1268)
);

AOI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1111),
.A2(n_1107),
.B(n_1076),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1236),
.A2(n_998),
.B(n_1097),
.Y(n_1270)
);

OAI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_1109),
.A2(n_1078),
.B(n_1108),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1076),
.B1(n_1105),
.B2(n_1030),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1147),
.B(n_1031),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1158),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1118),
.A2(n_929),
.A3(n_1017),
.B(n_957),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1165),
.A2(n_979),
.B(n_957),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1168),
.A2(n_953),
.B(n_1030),
.C(n_1101),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1263),
.A2(n_968),
.B(n_969),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1129),
.A2(n_968),
.B(n_969),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1280)
);

AOI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1202),
.A2(n_1010),
.B(n_1076),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1238),
.A2(n_1088),
.B(n_1062),
.Y(n_1282)
);

AOI21xp33_ASAP7_75t_L g1283 ( 
.A1(n_1219),
.A2(n_1070),
.B(n_1011),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1167),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1201),
.A2(n_1248),
.B(n_1148),
.Y(n_1285)
);

AND2x6_ASAP7_75t_L g1286 ( 
.A(n_1206),
.B(n_974),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1113),
.A2(n_974),
.B(n_1018),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1185),
.B(n_1072),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1112),
.A2(n_1088),
.B(n_1070),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1235),
.Y(n_1290)
);

AOI221x1_ASAP7_75t_L g1291 ( 
.A1(n_1210),
.A2(n_1090),
.B1(n_1083),
.B2(n_1004),
.C(n_979),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1117),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1213),
.B(n_993),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1131),
.A2(n_993),
.B(n_1004),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1122),
.A2(n_1017),
.B(n_1096),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1187),
.A2(n_1099),
.B1(n_1083),
.B2(n_1090),
.Y(n_1296)
);

AOI211x1_ASAP7_75t_L g1297 ( 
.A1(n_1214),
.A2(n_1078),
.B(n_1066),
.C(n_1096),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1197),
.B(n_1255),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_L g1299 ( 
.A(n_1147),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1124),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1229),
.A2(n_1011),
.B(n_1086),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1128),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1134),
.A2(n_1083),
.A3(n_1090),
.B(n_1086),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1162),
.A2(n_1018),
.B(n_1083),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1230),
.A2(n_1018),
.B(n_1090),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1121),
.A2(n_1161),
.B(n_1144),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1160),
.B(n_1138),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1110),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1235),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1143),
.Y(n_1310)
);

NAND2xp33_ASAP7_75t_L g1311 ( 
.A(n_1116),
.B(n_1151),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1159),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1255),
.B(n_1242),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1243),
.A2(n_1245),
.B(n_1164),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1223),
.A2(n_1232),
.B1(n_1125),
.B2(n_1233),
.C(n_1237),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1175),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1217),
.A2(n_1218),
.B(n_1184),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1163),
.A2(n_1208),
.B(n_1239),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1253),
.B(n_1259),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1250),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1251),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1127),
.A2(n_1132),
.B(n_1228),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1147),
.A2(n_1206),
.B(n_1227),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1190),
.A2(n_1224),
.B1(n_1170),
.B2(n_1205),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1186),
.A2(n_1194),
.B(n_1181),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1264),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1191),
.B(n_1154),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1260),
.A2(n_1198),
.B(n_1199),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_1209),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1196),
.A2(n_1192),
.B1(n_1203),
.B2(n_1139),
.C(n_1234),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1226),
.A2(n_1178),
.B(n_1126),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1204),
.B(n_1140),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1254),
.A2(n_1267),
.A3(n_1179),
.B(n_1173),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1266),
.A2(n_1135),
.B(n_1136),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1200),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1175),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1212),
.A2(n_1227),
.B1(n_1180),
.B2(n_1222),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1266),
.A2(n_1262),
.B(n_1256),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1215),
.B(n_1265),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1157),
.A2(n_1189),
.B1(n_1231),
.B2(n_1216),
.C(n_1221),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1183),
.B(n_1120),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1141),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1149),
.A2(n_1133),
.B1(n_1150),
.B2(n_1152),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1261),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1156),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1220),
.A2(n_1157),
.B(n_1188),
.C(n_1155),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1182),
.A2(n_1225),
.B(n_1211),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1195),
.A2(n_1137),
.B(n_1166),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1176),
.A2(n_1151),
.B(n_1177),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1151),
.A2(n_1240),
.B(n_1182),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1172),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1171),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1151),
.B(n_1240),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_L g1355 ( 
.A(n_1141),
.B(n_1241),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1246),
.B(n_1110),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1172),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1211),
.A2(n_1225),
.B(n_1268),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1153),
.B(n_1110),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1146),
.A2(n_1123),
.B(n_1130),
.C(n_1142),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1172),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1156),
.B(n_1169),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1195),
.A2(n_1174),
.B(n_1257),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1156),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1258),
.A2(n_1195),
.A3(n_1244),
.B(n_1207),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1130),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1258),
.A2(n_1169),
.B(n_1174),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1123),
.A2(n_1142),
.B(n_1257),
.C(n_1258),
.Y(n_1368)
);

INVx3_ASAP7_75t_R g1369 ( 
.A(n_1193),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1235),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1109),
.A2(n_1119),
.B(n_1115),
.C(n_1219),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1109),
.B(n_636),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1117),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1138),
.B(n_1000),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1109),
.B(n_756),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1117),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1118),
.A2(n_1102),
.A3(n_1134),
.B(n_1125),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1109),
.A2(n_1119),
.B(n_1115),
.C(n_1219),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1109),
.B(n_756),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1110),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1109),
.B(n_756),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1117),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1109),
.B(n_756),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1160),
.B(n_778),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1236),
.A2(n_1125),
.B(n_1121),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1160),
.B(n_778),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1392)
);

NAND3x1_ASAP7_75t_L g1393 ( 
.A(n_1188),
.B(n_756),
.C(n_775),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1238),
.A2(n_1145),
.B(n_1114),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1246),
.B(n_971),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1236),
.A2(n_1114),
.B(n_1111),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1114),
.A2(n_1236),
.B(n_1201),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1109),
.A2(n_1119),
.B1(n_773),
.B2(n_1219),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1109),
.A2(n_756),
.B1(n_822),
.B2(n_824),
.C(n_870),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1109),
.B(n_756),
.Y(n_1403)
);

NAND2xp33_ASAP7_75t_L g1404 ( 
.A(n_1109),
.B(n_846),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_SL g1405 ( 
.A(n_1167),
.Y(n_1405)
);

INVx8_ASAP7_75t_L g1406 ( 
.A(n_1147),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1117),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1114),
.A2(n_1236),
.B(n_1201),
.Y(n_1411)
);

AOI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1111),
.A2(n_1219),
.B(n_1112),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1238),
.A2(n_1145),
.B(n_1114),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1115),
.A2(n_756),
.B1(n_775),
.B2(n_612),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1117),
.Y(n_1416)
);

OA22x2_ASAP7_75t_L g1417 ( 
.A1(n_1213),
.A2(n_821),
.B1(n_632),
.B2(n_1087),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1109),
.B(n_636),
.Y(n_1418)
);

AOI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1111),
.A2(n_1219),
.B(n_1112),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1114),
.A2(n_1236),
.B(n_1201),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1147),
.B(n_989),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1209),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1109),
.B(n_756),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1109),
.B(n_756),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1167),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1259),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1431)
);

AO31x2_ASAP7_75t_L g1432 ( 
.A1(n_1118),
.A2(n_1102),
.A3(n_1134),
.B(n_1125),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1165),
.A2(n_1263),
.B(n_1131),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1114),
.A2(n_1236),
.B(n_1201),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1209),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1158),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1202),
.A2(n_1252),
.B(n_1238),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1336),
.Y(n_1439)
);

CKINVDCx6p67_ASAP7_75t_R g1440 ( 
.A(n_1284),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1351),
.B(n_1286),
.Y(n_1441)
);

AO31x2_ASAP7_75t_L g1442 ( 
.A1(n_1291),
.A2(n_1368),
.A3(n_1285),
.B(n_1349),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1379),
.C(n_1371),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1292),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1405),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1382),
.A2(n_1384),
.B1(n_1403),
.B2(n_1425),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1300),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1426),
.B(n_1307),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1402),
.A2(n_1401),
.B1(n_1393),
.B2(n_1325),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1401),
.A2(n_1417),
.B1(n_1412),
.B2(n_1419),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1427),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1428),
.B(n_1320),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1391),
.A2(n_1408),
.B(n_1407),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1423),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1410),
.A2(n_1424),
.B(n_1420),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1398),
.A2(n_1434),
.B(n_1421),
.Y(n_1459)
);

NAND2x2_ASAP7_75t_L g1460 ( 
.A(n_1290),
.B(n_1309),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1429),
.A2(n_1433),
.B(n_1431),
.Y(n_1461)
);

INVx5_ASAP7_75t_L g1462 ( 
.A(n_1286),
.Y(n_1462)
);

OR2x6_ASAP7_75t_L g1463 ( 
.A(n_1324),
.B(n_1406),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1315),
.A2(n_1306),
.B(n_1326),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1437),
.A2(n_1279),
.B(n_1294),
.Y(n_1465)
);

AOI22x1_ASAP7_75t_L g1466 ( 
.A1(n_1318),
.A2(n_1394),
.B1(n_1413),
.B2(n_1329),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1351),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1286),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1302),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1325),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1308),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1406),
.B(n_1289),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1345),
.B(n_1386),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1289),
.A2(n_1415),
.B(n_1280),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1280),
.A2(n_1385),
.B(n_1415),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_L g1476 ( 
.A(n_1286),
.B(n_1350),
.Y(n_1476)
);

BUFx10_ASAP7_75t_L g1477 ( 
.A(n_1359),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1335),
.A2(n_1298),
.B(n_1363),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1295),
.A2(n_1287),
.B(n_1276),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1298),
.A2(n_1400),
.B(n_1396),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1308),
.Y(n_1482)
);

NAND2x1p5_ASAP7_75t_L g1483 ( 
.A(n_1299),
.B(n_1308),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1332),
.A2(n_1305),
.B(n_1278),
.Y(n_1484)
);

OR2x6_ASAP7_75t_SL g1485 ( 
.A(n_1390),
.B(n_1342),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1381),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1281),
.A2(n_1323),
.B(n_1282),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1353),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1282),
.A2(n_1301),
.B(n_1385),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1389),
.A2(n_1400),
.B(n_1392),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1347),
.B(n_1341),
.C(n_1331),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1389),
.A2(n_1396),
.B(n_1397),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1392),
.A2(n_1430),
.B(n_1397),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1320),
.B(n_1330),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1430),
.A2(n_1304),
.B(n_1339),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1288),
.A2(n_1270),
.B(n_1387),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1310),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1288),
.A2(n_1270),
.B(n_1387),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1348),
.A2(n_1354),
.B(n_1350),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1312),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1328),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1435),
.B(n_1404),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1354),
.A2(n_1313),
.B(n_1318),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1313),
.A2(n_1316),
.B(n_1362),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1297),
.B(n_1271),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1314),
.B(n_1409),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1314),
.B(n_1416),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1334),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1362),
.A2(n_1418),
.B(n_1372),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_SL g1510 ( 
.A(n_1343),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1338),
.B(n_1344),
.Y(n_1511)
);

CKINVDCx8_ASAP7_75t_R g1512 ( 
.A(n_1381),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1346),
.Y(n_1513)
);

NOR2xp67_ASAP7_75t_L g1514 ( 
.A(n_1370),
.B(n_1272),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1283),
.A2(n_1338),
.B(n_1311),
.Y(n_1515)
);

AO221x2_ASAP7_75t_L g1516 ( 
.A1(n_1417),
.A2(n_1296),
.B1(n_1365),
.B2(n_1321),
.C(n_1383),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1364),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1367),
.A2(n_1327),
.B(n_1317),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1334),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1274),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1322),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1373),
.B(n_1377),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1269),
.A2(n_1283),
.B(n_1340),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1317),
.A2(n_1337),
.B(n_1340),
.Y(n_1524)
);

INVxp67_ASAP7_75t_SL g1525 ( 
.A(n_1273),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1293),
.A2(n_1366),
.B(n_1361),
.Y(n_1526)
);

OAI21xp33_ASAP7_75t_L g1527 ( 
.A1(n_1360),
.A2(n_1269),
.B(n_1344),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1366),
.A2(n_1355),
.B1(n_1352),
.B2(n_1357),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1436),
.A2(n_1432),
.B(n_1378),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_SL g1530 ( 
.A1(n_1422),
.A2(n_1277),
.B(n_1273),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1378),
.A2(n_1432),
.B(n_1303),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1275),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1378),
.A2(n_1432),
.B(n_1303),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1395),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1275),
.Y(n_1535)
);

AO32x2_ASAP7_75t_L g1536 ( 
.A1(n_1275),
.A2(n_1303),
.A3(n_1365),
.B1(n_1422),
.B2(n_1369),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1395),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1324),
.B(n_1406),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1351),
.B(n_1286),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_SL g1541 ( 
.A(n_1338),
.B(n_1147),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1371),
.B2(n_1379),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1333),
.B(n_1380),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1369),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1292),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1428),
.B(n_1345),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_SL g1551 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1371),
.C(n_1379),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1299),
.B(n_713),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1371),
.B2(n_1379),
.Y(n_1556)
);

AO31x2_ASAP7_75t_L g1557 ( 
.A1(n_1291),
.A2(n_1368),
.A3(n_1285),
.B(n_1349),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1336),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1292),
.Y(n_1559)
);

A2O1A1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1371),
.C(n_1379),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1398),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1292),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1371),
.B2(n_1379),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1405),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1371),
.B2(n_1379),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1333),
.B(n_1380),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1405),
.Y(n_1568)
);

CKINVDCx11_ASAP7_75t_R g1569 ( 
.A(n_1336),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1286),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1414),
.B(n_1380),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1286),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1401),
.B(n_1109),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1289),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1414),
.A2(n_1380),
.B(n_1379),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1324),
.B(n_1406),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1292),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1428),
.B(n_1345),
.Y(n_1583)
);

CKINVDCx16_ASAP7_75t_R g1584 ( 
.A(n_1353),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1292),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1334),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1351),
.B(n_1286),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1333),
.B(n_1380),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1292),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1405),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1405),
.Y(n_1595)
);

CKINVDCx6p67_ASAP7_75t_R g1596 ( 
.A(n_1284),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1286),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1398),
.A2(n_1411),
.B(n_1399),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1401),
.B(n_1109),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1428),
.B(n_1345),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1319),
.A2(n_1388),
.B(n_1375),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1475),
.Y(n_1603)
);

CKINVDCx16_ASAP7_75t_R g1604 ( 
.A(n_1547),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1542),
.A2(n_1556),
.B(n_1564),
.C(n_1566),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1571),
.A2(n_1443),
.B1(n_1450),
.B2(n_1577),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1575),
.A2(n_1599),
.B(n_1551),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_SL g1608 ( 
.A1(n_1502),
.A2(n_1539),
.B(n_1438),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1547),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1439),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1571),
.A2(n_1560),
.B1(n_1501),
.B2(n_1470),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1455),
.B(n_1494),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1448),
.B(n_1446),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1550),
.B(n_1591),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1475),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1473),
.B(n_1506),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1507),
.B(n_1452),
.Y(n_1618)
);

AOI21x1_ASAP7_75t_SL g1619 ( 
.A1(n_1546),
.A2(n_1592),
.B(n_1567),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1560),
.A2(n_1501),
.B1(n_1452),
.B2(n_1561),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1441),
.B(n_1540),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1549),
.B(n_1583),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1522),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1457),
.B(n_1575),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1464),
.A2(n_1458),
.B(n_1456),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1558),
.B(n_1522),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1444),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1464),
.A2(n_1458),
.B(n_1456),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1447),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1493),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1493),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1461),
.A2(n_1543),
.B(n_1449),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1469),
.B(n_1497),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1515),
.A2(n_1491),
.B(n_1576),
.C(n_1511),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1517),
.B(n_1477),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1490),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1477),
.B(n_1485),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1500),
.B(n_1521),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1499),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1454),
.B(n_1513),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1548),
.B(n_1559),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1576),
.A2(n_1511),
.B(n_1527),
.C(n_1476),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1441),
.B(n_1540),
.Y(n_1643)
);

O2A1O1Ixp5_ASAP7_75t_L g1644 ( 
.A1(n_1528),
.A2(n_1540),
.B(n_1590),
.C(n_1441),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1562),
.B(n_1582),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1449),
.A2(n_1572),
.B(n_1600),
.Y(n_1646)
);

O2A1O1Ixp5_ASAP7_75t_L g1647 ( 
.A1(n_1590),
.A2(n_1525),
.B(n_1593),
.C(n_1585),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1511),
.A2(n_1460),
.B1(n_1510),
.B2(n_1596),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1440),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1520),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1499),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1478),
.B(n_1462),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1471),
.B(n_1486),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1482),
.B(n_1516),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1481),
.B(n_1474),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1496),
.A2(n_1498),
.B(n_1503),
.C(n_1504),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1516),
.B(n_1569),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1481),
.B(n_1474),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1490),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1584),
.Y(n_1661)
);

BUFx4f_ASAP7_75t_SL g1662 ( 
.A(n_1445),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1503),
.B(n_1492),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1496),
.A2(n_1498),
.B(n_1504),
.C(n_1514),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1541),
.A2(n_1581),
.B(n_1463),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1492),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1488),
.A2(n_1466),
.B1(n_1472),
.B2(n_1505),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1472),
.B(n_1534),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1463),
.A2(n_1581),
.B(n_1538),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1451),
.A2(n_1545),
.B(n_1598),
.Y(n_1670)
);

AOI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1554),
.A2(n_1565),
.B(n_1594),
.C(n_1526),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1505),
.A2(n_1568),
.B1(n_1445),
.B2(n_1595),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1505),
.A2(n_1568),
.B1(n_1595),
.B2(n_1459),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1530),
.A2(n_1552),
.B(n_1451),
.C(n_1459),
.Y(n_1674)
);

O2A1O1Ixp5_ASAP7_75t_L g1675 ( 
.A1(n_1532),
.A2(n_1519),
.B(n_1508),
.C(n_1587),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1512),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1463),
.A2(n_1538),
.B(n_1581),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1537),
.B(n_1589),
.Y(n_1678)
);

OA22x2_ASAP7_75t_L g1679 ( 
.A1(n_1538),
.A2(n_1467),
.B1(n_1529),
.B2(n_1533),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1537),
.B(n_1589),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1451),
.A2(n_1545),
.B1(n_1598),
.B2(n_1552),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1545),
.A2(n_1589),
.B1(n_1598),
.B2(n_1586),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1468),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1489),
.A2(n_1533),
.B(n_1531),
.C(n_1487),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1479),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1467),
.B(n_1518),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1552),
.B(n_1586),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1586),
.B(n_1483),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1570),
.A2(n_1597),
.B1(n_1573),
.B2(n_1479),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1479),
.A2(n_1487),
.B(n_1602),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1536),
.B(n_1509),
.Y(n_1691)
);

NOR2xp67_ASAP7_75t_L g1692 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1544),
.A2(n_1555),
.B(n_1580),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1524),
.B(n_1531),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1495),
.A2(n_1484),
.B(n_1465),
.C(n_1442),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1442),
.Y(n_1697)
);

CKINVDCx8_ASAP7_75t_R g1698 ( 
.A(n_1557),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1557),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1557),
.B(n_1484),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1553),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1553),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1563),
.A2(n_1578),
.B1(n_1572),
.B2(n_1574),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1579),
.B(n_1580),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1588),
.B(n_1480),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1571),
.A2(n_1414),
.B1(n_1443),
.B2(n_1450),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1455),
.B(n_1494),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1542),
.A2(n_1556),
.B(n_1566),
.C(n_1564),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1571),
.A2(n_1414),
.B1(n_1443),
.B2(n_1450),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1547),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1571),
.A2(n_1414),
.B1(n_1443),
.B2(n_1450),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_SL g1713 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1575),
.A2(n_1419),
.B(n_1412),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1444),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1455),
.B(n_1494),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1453),
.B(n_1546),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1443),
.A2(n_1419),
.B(n_1412),
.C(n_1371),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1453),
.B(n_1546),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1670),
.A2(n_1690),
.B(n_1696),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1656),
.B(n_1623),
.Y(n_1721)
);

NAND3xp33_ASAP7_75t_L g1722 ( 
.A(n_1707),
.B(n_1712),
.C(n_1710),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1629),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1613),
.B(n_1708),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1665),
.B(n_1669),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1620),
.A2(n_1612),
.B1(n_1606),
.B2(n_1654),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1678),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1695),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1693),
.A2(n_1659),
.B(n_1655),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1626),
.B(n_1691),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1715),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1716),
.B(n_1618),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1637),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1633),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1638),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1680),
.Y(n_1736)
);

AO21x2_ASAP7_75t_L g1737 ( 
.A1(n_1696),
.A2(n_1682),
.B(n_1681),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1677),
.B(n_1642),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1645),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1652),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1614),
.B(n_1627),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1624),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1641),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1639),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1630),
.Y(n_1745)
);

OAI222xp33_ASAP7_75t_L g1746 ( 
.A1(n_1605),
.A2(n_1709),
.B1(n_1634),
.B2(n_1607),
.C1(n_1714),
.C2(n_1658),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1611),
.Y(n_1747)
);

AO21x2_ASAP7_75t_L g1748 ( 
.A1(n_1687),
.A2(n_1684),
.B(n_1700),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1621),
.B(n_1643),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1630),
.Y(n_1750)
);

AO21x2_ASAP7_75t_L g1751 ( 
.A1(n_1699),
.A2(n_1697),
.B(n_1657),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_1604),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1631),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1631),
.B(n_1718),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1650),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1686),
.B(n_1688),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1640),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1685),
.B(n_1698),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1668),
.A2(n_1622),
.B1(n_1673),
.B2(n_1683),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1685),
.B(n_1698),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1635),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1603),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1717),
.B(n_1719),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1603),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1616),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1616),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1653),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1704),
.A2(n_1664),
.B(n_1663),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1718),
.B(n_1617),
.Y(n_1769)
);

AO21x2_ASAP7_75t_L g1770 ( 
.A1(n_1692),
.A2(n_1674),
.B(n_1703),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1636),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1636),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1660),
.B(n_1666),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1615),
.A2(n_1667),
.B1(n_1671),
.B2(n_1648),
.C(n_1672),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1666),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1675),
.Y(n_1776)
);

BUFx12f_ASAP7_75t_L g1777 ( 
.A(n_1649),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1701),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1644),
.Y(n_1779)
);

AO21x2_ASAP7_75t_L g1780 ( 
.A1(n_1702),
.A2(n_1706),
.B(n_1705),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1651),
.Y(n_1781)
);

NOR3xp33_ASAP7_75t_SL g1782 ( 
.A(n_1722),
.B(n_1609),
.C(n_1711),
.Y(n_1782)
);

NOR2x1p5_ASAP7_75t_L g1783 ( 
.A(n_1754),
.B(n_1610),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1754),
.B(n_1729),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1781),
.B(n_1651),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1727),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1778),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1722),
.B(n_1661),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1720),
.A2(n_1625),
.B(n_1628),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1744),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1777),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1780),
.B(n_1632),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1740),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1780),
.B(n_1632),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1780),
.B(n_1646),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1745),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1780),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1730),
.B(n_1646),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1730),
.B(n_1748),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1726),
.A2(n_1769),
.B1(n_1732),
.B2(n_1738),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1745),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1751),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1748),
.B(n_1646),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1748),
.B(n_1694),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1751),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1750),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1729),
.B(n_1689),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1772),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1753),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1748),
.B(n_1694),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1751),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1753),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1723),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1741),
.B(n_1625),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1723),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1776),
.B(n_1647),
.C(n_1661),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1729),
.B(n_1741),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1768),
.B(n_1679),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1744),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1731),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1808),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1784),
.B(n_1742),
.Y(n_1822)
);

NAND2x1_ASAP7_75t_L g1823 ( 
.A(n_1819),
.B(n_1757),
.Y(n_1823)
);

OAI321xp33_ASAP7_75t_L g1824 ( 
.A1(n_1800),
.A2(n_1738),
.A3(n_1779),
.B1(n_1774),
.B2(n_1769),
.C(n_1759),
.Y(n_1824)
);

OR2x6_ASAP7_75t_L g1825 ( 
.A(n_1816),
.B(n_1738),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1787),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1749),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1813),
.Y(n_1828)
);

NOR2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1791),
.B(n_1610),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1816),
.A2(n_1746),
.B(n_1725),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1818),
.A2(n_1779),
.B1(n_1738),
.B2(n_1774),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1813),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1800),
.A2(n_1732),
.B1(n_1733),
.B2(n_1738),
.C(n_1776),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_SL g1834 ( 
.A(n_1793),
.B(n_1725),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1808),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1817),
.B(n_1734),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1813),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1820),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1820),
.Y(n_1839)
);

AO21x2_ASAP7_75t_L g1840 ( 
.A1(n_1802),
.A2(n_1770),
.B(n_1765),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1793),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1784),
.B(n_1728),
.C(n_1773),
.Y(n_1842)
);

OAI21x1_ASAP7_75t_SL g1843 ( 
.A1(n_1790),
.A2(n_1757),
.B(n_1713),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1820),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1816),
.A2(n_1733),
.B1(n_1738),
.B2(n_1734),
.C(n_1735),
.Y(n_1845)
);

AOI33xp33_ASAP7_75t_L g1846 ( 
.A1(n_1792),
.A2(n_1763),
.A3(n_1743),
.B1(n_1728),
.B2(n_1735),
.B3(n_1739),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1784),
.A2(n_1746),
.B1(n_1739),
.B2(n_1743),
.C(n_1770),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1788),
.A2(n_1752),
.B1(n_1777),
.B2(n_1662),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1815),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1791),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1782),
.A2(n_1788),
.B1(n_1783),
.B2(n_1799),
.Y(n_1851)
);

AOI331xp33_ASAP7_75t_L g1852 ( 
.A1(n_1796),
.A2(n_1747),
.A3(n_1771),
.B1(n_1775),
.B2(n_1619),
.B3(n_1662),
.C1(n_1608),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1815),
.Y(n_1853)
);

INVx5_ASAP7_75t_SL g1854 ( 
.A(n_1785),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1818),
.A2(n_1770),
.B1(n_1760),
.B2(n_1758),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1786),
.B(n_1740),
.Y(n_1856)
);

AO21x2_ASAP7_75t_L g1857 ( 
.A1(n_1802),
.A2(n_1770),
.B(n_1764),
.Y(n_1857)
);

NOR4xp25_ASAP7_75t_SL g1858 ( 
.A(n_1819),
.B(n_1796),
.C(n_1812),
.D(n_1809),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1799),
.B(n_1767),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_SL g1860 ( 
.A1(n_1799),
.A2(n_1758),
.B(n_1760),
.Y(n_1860)
);

AOI33xp33_ASAP7_75t_L g1861 ( 
.A1(n_1792),
.A2(n_1763),
.A3(n_1728),
.B1(n_1761),
.B2(n_1775),
.B3(n_1771),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1818),
.A2(n_1724),
.B1(n_1736),
.B2(n_1727),
.C(n_1721),
.Y(n_1862)
);

NAND4xp25_ASAP7_75t_SL g1863 ( 
.A(n_1799),
.B(n_1676),
.C(n_1761),
.D(n_1777),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1818),
.A2(n_1764),
.B1(n_1762),
.B2(n_1765),
.C(n_1766),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1817),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1782),
.Y(n_1866)
);

AOI221xp5_ASAP7_75t_L g1867 ( 
.A1(n_1817),
.A2(n_1766),
.B1(n_1762),
.B2(n_1736),
.C(n_1756),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1793),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1783),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1803),
.A2(n_1737),
.B1(n_1721),
.B2(n_1773),
.C(n_1755),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1814),
.B(n_1786),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1828),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1832),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1847),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1859),
.B(n_1798),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1826),
.A2(n_1789),
.B(n_1802),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1840),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1837),
.Y(n_1878)
);

OA21x2_ASAP7_75t_L g1879 ( 
.A1(n_1870),
.A2(n_1789),
.B(n_1802),
.Y(n_1879)
);

INVx4_ASAP7_75t_L g1880 ( 
.A(n_1850),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1838),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1859),
.B(n_1798),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1839),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1840),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1822),
.B(n_1814),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1840),
.Y(n_1886)
);

INVx4_ASAP7_75t_SL g1887 ( 
.A(n_1825),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1844),
.Y(n_1888)
);

INVx3_ASAP7_75t_SL g1889 ( 
.A(n_1825),
.Y(n_1889)
);

OA21x2_ASAP7_75t_L g1890 ( 
.A1(n_1830),
.A2(n_1805),
.B(n_1811),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1850),
.B(n_1609),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1857),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1849),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1846),
.B(n_1814),
.Y(n_1894)
);

INVx4_ASAP7_75t_L g1895 ( 
.A(n_1825),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1821),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1835),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1853),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1868),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1848),
.B(n_1711),
.Y(n_1900)
);

AND4x1_ASAP7_75t_L g1901 ( 
.A(n_1831),
.B(n_1803),
.C(n_1804),
.D(n_1810),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1836),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1857),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1846),
.B(n_1814),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1824),
.A2(n_1855),
.B(n_1845),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1861),
.B(n_1796),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1871),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1871),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1861),
.B(n_1801),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1869),
.B(n_1649),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1834),
.B(n_1790),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1827),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1822),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1896),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1876),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1874),
.B(n_1867),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.B(n_1899),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1911),
.B(n_1827),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1911),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1911),
.B(n_1827),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1874),
.A2(n_1866),
.B1(n_1851),
.B2(n_1833),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1872),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1899),
.B(n_1875),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1894),
.B(n_1864),
.Y(n_1924)
);

AND2x4_ASAP7_75t_SL g1925 ( 
.A(n_1880),
.B(n_1895),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1906),
.B(n_1842),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1905),
.A2(n_1860),
.B(n_1866),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1872),
.Y(n_1928)
);

NAND2x1_ASAP7_75t_L g1929 ( 
.A(n_1897),
.B(n_1843),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1873),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1882),
.B(n_1854),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1882),
.B(n_1854),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1894),
.B(n_1798),
.Y(n_1933)
);

NAND4xp25_ASAP7_75t_SL g1934 ( 
.A(n_1904),
.B(n_1795),
.C(n_1794),
.D(n_1792),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1882),
.B(n_1880),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1873),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1878),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1880),
.B(n_1854),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1897),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1887),
.B(n_1803),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1896),
.Y(n_1941)
);

NAND4xp25_ASAP7_75t_L g1942 ( 
.A(n_1904),
.B(n_1792),
.C(n_1794),
.D(n_1795),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1878),
.Y(n_1943)
);

NOR3xp33_ASAP7_75t_L g1944 ( 
.A(n_1905),
.B(n_1863),
.C(n_1797),
.Y(n_1944)
);

OAI33xp33_ASAP7_75t_L g1945 ( 
.A1(n_1909),
.A2(n_1865),
.A3(n_1797),
.B1(n_1807),
.B2(n_1856),
.B3(n_1806),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1881),
.Y(n_1946)
);

CKINVDCx16_ASAP7_75t_R g1947 ( 
.A(n_1880),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1876),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1909),
.A2(n_1852),
.B(n_1856),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1907),
.B(n_1854),
.Y(n_1950)
);

NAND2x1_ASAP7_75t_L g1951 ( 
.A(n_1895),
.B(n_1841),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1900),
.B(n_1869),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1881),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1907),
.B(n_1868),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1924),
.B(n_1908),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1939),
.B(n_1908),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1922),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1922),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1928),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1923),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1914),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1928),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1923),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1926),
.B(n_1902),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1930),
.Y(n_1965)
);

OAI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1927),
.A2(n_1916),
.B(n_1949),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1939),
.B(n_1902),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1930),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1941),
.B(n_1901),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1926),
.B(n_1901),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1954),
.B(n_1883),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1915),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1936),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1915),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1936),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1954),
.B(n_1883),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1913),
.B(n_1885),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1915),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1937),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1947),
.B(n_1888),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1947),
.B(n_1888),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1937),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1948),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1927),
.B(n_1893),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1942),
.A2(n_1885),
.B(n_1804),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1913),
.B(n_1893),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1942),
.B(n_1898),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1944),
.B(n_1898),
.Y(n_1988)
);

NOR2xp67_ASAP7_75t_L g1989 ( 
.A(n_1919),
.B(n_1895),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1943),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1948),
.Y(n_1991)
);

NAND2xp33_ASAP7_75t_L g1992 ( 
.A(n_1921),
.B(n_1829),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1935),
.B(n_1858),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1966),
.B(n_1943),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1970),
.A2(n_1921),
.B1(n_1895),
.B2(n_1889),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1960),
.B(n_1935),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1963),
.B(n_1917),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1963),
.B(n_1917),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1961),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1993),
.B(n_1912),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1955),
.B(n_1946),
.Y(n_2002)
);

CKINVDCx16_ASAP7_75t_R g2003 ( 
.A(n_1955),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1957),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1957),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1993),
.B(n_1912),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1992),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1977),
.B(n_1933),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1959),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1989),
.B(n_1940),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1959),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1988),
.B(n_1918),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1992),
.A2(n_1945),
.B(n_1934),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1964),
.B(n_1946),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1962),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_1956),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1962),
.Y(n_2017)
);

INVx4_ASAP7_75t_L g2018 ( 
.A(n_1965),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1969),
.A2(n_1879),
.B1(n_1940),
.B2(n_1889),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1987),
.B(n_1918),
.Y(n_2020)
);

NOR2x1_ASAP7_75t_L g2021 ( 
.A(n_1984),
.B(n_1951),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2005),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1994),
.A2(n_1929),
.B(n_1967),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2003),
.A2(n_1987),
.B1(n_1985),
.B2(n_1925),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_2003),
.A2(n_1879),
.B1(n_1940),
.B2(n_1991),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2005),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2017),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2000),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1998),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_2007),
.B(n_2000),
.Y(n_2030)
);

NOR3xp33_ASAP7_75t_L g2031 ( 
.A(n_1994),
.B(n_1964),
.C(n_1965),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1995),
.A2(n_1879),
.B1(n_1940),
.B2(n_1972),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2017),
.Y(n_2033)
);

OAI221xp5_ASAP7_75t_SL g2034 ( 
.A1(n_2007),
.A2(n_2013),
.B1(n_2019),
.B2(n_2016),
.C(n_2012),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1996),
.Y(n_2035)
);

AOI222xp33_ASAP7_75t_L g2036 ( 
.A1(n_2016),
.A2(n_1986),
.B1(n_1974),
.B2(n_1991),
.C1(n_1983),
.C2(n_1972),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1998),
.B(n_1971),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_2008),
.B(n_1977),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1998),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_2008),
.B(n_1976),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_SL g2041 ( 
.A(n_1995),
.B(n_1910),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_2000),
.B(n_1952),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1999),
.B(n_1925),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_R g2045 ( 
.A1(n_2034),
.A2(n_1996),
.B1(n_2013),
.B2(n_2011),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2029),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_2039),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2038),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2022),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2030),
.B(n_1999),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2030),
.B(n_2009),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2028),
.Y(n_2052)
);

OAI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_2025),
.A2(n_1889),
.B1(n_1879),
.B2(n_2021),
.Y(n_2053)
);

INVx1_ASAP7_75t_SL g2054 ( 
.A(n_2044),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2042),
.B(n_1999),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_SL g2056 ( 
.A(n_2042),
.B(n_1997),
.Y(n_2056)
);

AND2x4_ASAP7_75t_L g2057 ( 
.A(n_2028),
.B(n_1997),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2031),
.A2(n_1879),
.B1(n_1983),
.B2(n_1974),
.Y(n_2058)
);

NOR4xp25_ASAP7_75t_L g2059 ( 
.A(n_2052),
.B(n_2034),
.C(n_2026),
.D(n_2033),
.Y(n_2059)
);

AOI211xp5_ASAP7_75t_L g2060 ( 
.A1(n_2053),
.A2(n_2031),
.B(n_2023),
.C(n_2032),
.Y(n_2060)
);

AOI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2058),
.A2(n_2043),
.B1(n_2035),
.B2(n_2024),
.C(n_2002),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2055),
.B(n_2012),
.Y(n_2062)
);

NAND3xp33_ASAP7_75t_SL g2063 ( 
.A(n_2056),
.B(n_2036),
.C(n_2041),
.Y(n_2063)
);

NAND4xp75_ASAP7_75t_L g2064 ( 
.A(n_2051),
.B(n_2021),
.C(n_2027),
.D(n_2006),
.Y(n_2064)
);

NAND4xp75_ASAP7_75t_L g2065 ( 
.A(n_2050),
.B(n_2001),
.C(n_2006),
.D(n_2020),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2048),
.A2(n_2001),
.B1(n_2006),
.B2(n_2012),
.Y(n_2066)
);

AOI221xp5_ASAP7_75t_L g2067 ( 
.A1(n_2045),
.A2(n_2002),
.B1(n_2014),
.B2(n_2037),
.C(n_2015),
.Y(n_2067)
);

AO22x1_ASAP7_75t_L g2068 ( 
.A1(n_2050),
.A2(n_2018),
.B1(n_2009),
.B2(n_2010),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2055),
.B(n_2057),
.Y(n_2069)
);

AOI311xp33_ASAP7_75t_L g2070 ( 
.A1(n_2049),
.A2(n_2011),
.A3(n_2004),
.B(n_2015),
.C(n_2014),
.Y(n_2070)
);

OAI21xp33_ASAP7_75t_L g2071 ( 
.A1(n_2054),
.A2(n_2001),
.B(n_2020),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2069),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2059),
.A2(n_2048),
.B1(n_2049),
.B2(n_2047),
.C(n_2046),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2063),
.A2(n_2057),
.B1(n_2047),
.B2(n_2020),
.Y(n_2074)
);

AOI221x1_ASAP7_75t_L g2075 ( 
.A1(n_2071),
.A2(n_2046),
.B1(n_2057),
.B2(n_2009),
.C(n_2018),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2062),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2066),
.B(n_2040),
.Y(n_2077)
);

O2A1O1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_2060),
.A2(n_2004),
.B(n_1973),
.C(n_1975),
.Y(n_2078)
);

OAI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2067),
.A2(n_2018),
.B1(n_2009),
.B2(n_1951),
.C(n_1978),
.Y(n_2079)
);

OAI31xp33_ASAP7_75t_L g2080 ( 
.A1(n_2079),
.A2(n_1925),
.A3(n_2010),
.B(n_2064),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2073),
.B(n_2065),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2074),
.B(n_2068),
.Y(n_2082)
);

XOR2x2_ASAP7_75t_L g2083 ( 
.A(n_2077),
.B(n_2061),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2072),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2076),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2078),
.B(n_1997),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2075),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2084),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2086),
.B(n_2018),
.Y(n_2089)
);

CKINVDCx16_ASAP7_75t_R g2090 ( 
.A(n_2085),
.Y(n_2090)
);

AOI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2081),
.A2(n_2010),
.B(n_2070),
.C(n_1990),
.Y(n_2091)
);

AND3x4_ASAP7_75t_L g2092 ( 
.A(n_2083),
.B(n_2010),
.C(n_1978),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2087),
.B(n_1980),
.Y(n_2093)
);

NOR3x2_ASAP7_75t_L g2094 ( 
.A(n_2090),
.B(n_2081),
.C(n_2080),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2092),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2088),
.Y(n_2096)
);

NOR4xp25_ASAP7_75t_L g2097 ( 
.A(n_2093),
.B(n_2082),
.C(n_1973),
.D(n_1990),
.Y(n_2097)
);

OA22x2_ASAP7_75t_L g2098 ( 
.A1(n_2095),
.A2(n_2089),
.B1(n_2091),
.B2(n_2010),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2096),
.Y(n_2099)
);

AOI322xp5_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_2094),
.A3(n_2097),
.B1(n_1948),
.B2(n_1982),
.C1(n_1968),
.C2(n_1975),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2098),
.A2(n_1982),
.B1(n_1968),
.B2(n_1979),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2100),
.B(n_1958),
.Y(n_2102)
);

AO22x2_ASAP7_75t_L g2103 ( 
.A1(n_2101),
.A2(n_1981),
.B1(n_1919),
.B2(n_1929),
.Y(n_2103)
);

AO22x2_ASAP7_75t_L g2104 ( 
.A1(n_2102),
.A2(n_1919),
.B1(n_1953),
.B2(n_1950),
.Y(n_2104)
);

AO22x2_ASAP7_75t_L g2105 ( 
.A1(n_2103),
.A2(n_1919),
.B1(n_1953),
.B2(n_1950),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_SL g2106 ( 
.A1(n_2104),
.A2(n_1891),
.B1(n_1676),
.B2(n_1862),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_SL g2107 ( 
.A1(n_2105),
.A2(n_1890),
.B1(n_1823),
.B2(n_1841),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_2106),
.A2(n_1920),
.B(n_1938),
.Y(n_2108)
);

AOI22x1_ASAP7_75t_L g2109 ( 
.A1(n_2108),
.A2(n_2107),
.B1(n_1938),
.B2(n_1920),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_1884),
.B(n_1877),
.Y(n_2110)
);

AOI222xp33_ASAP7_75t_L g2111 ( 
.A1(n_2110),
.A2(n_1892),
.B1(n_1877),
.B2(n_1884),
.C1(n_1886),
.C2(n_1903),
.Y(n_2111)
);

AOI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_2111),
.A2(n_1903),
.B1(n_1877),
.B2(n_1884),
.C(n_1886),
.Y(n_2112)
);

AOI211xp5_ASAP7_75t_L g2113 ( 
.A1(n_2112),
.A2(n_1932),
.B(n_1931),
.C(n_1886),
.Y(n_2113)
);


endmodule