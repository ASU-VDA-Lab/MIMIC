module fake_ariane_76_n_1765 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1765);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1765;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_64),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_22),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_132),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_77),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_17),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_28),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_47),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_59),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_73),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_93),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_75),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_81),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_30),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_110),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_104),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_49),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_92),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_156),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_84),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_139),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_58),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_45),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_37),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_19),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_36),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_98),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_24),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_47),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_46),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_1),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_69),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_39),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_34),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_49),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_86),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_130),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_62),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_143),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_63),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_90),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_54),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_46),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_31),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_102),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_40),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_53),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_99),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_78),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_159),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_108),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_116),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_134),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_105),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_88),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_15),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_45),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_37),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_22),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_74),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_33),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_67),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_94),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_125),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_19),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_55),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_96),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_66),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_31),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_121),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_106),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_76),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_10),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_54),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_17),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_117),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_4),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_51),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_51),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_41),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_48),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_42),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_27),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_112),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_23),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_23),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_20),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_3),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_151),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_123),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_163),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_231),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_232),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_166),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_172),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_172),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_173),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_161),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_173),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_175),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_223),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_161),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_182),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_182),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_168),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_189),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_168),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_189),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_221),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_188),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_188),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_217),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_274),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_235),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_235),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_232),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_274),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_279),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_220),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_221),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_235),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_195),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_200),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_235),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_202),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_202),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_229),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_200),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_178),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_291),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_260),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_260),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_230),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_262),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_281),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_180),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_205),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_281),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_205),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_232),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_232),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_291),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_291),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_273),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_292),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_214),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_291),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_292),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_293),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_165),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_293),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_214),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_345),
.B(n_209),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_224),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_331),
.A2(n_246),
.B1(n_317),
.B2(n_216),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_353),
.B(n_224),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_396),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_227),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_325),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_349),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_241),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_321),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_321),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_364),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_334),
.B(n_365),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_227),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_329),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_249),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_360),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_362),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_332),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_332),
.B(n_241),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_345),
.B(n_282),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_333),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_336),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_336),
.B(n_282),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_315),
.Y(n_444)
);

NOR2x1_ASAP7_75t_L g445 ( 
.A(n_337),
.B(n_338),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_335),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_337),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_372),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_335),
.A2(n_316),
.B1(n_318),
.B2(n_222),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_322),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_341),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_343),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_315),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_369),
.B(n_249),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_326),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_346),
.B(n_253),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_378),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_390),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_375),
.B(n_183),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_348),
.B(n_295),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_355),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_348),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_370),
.B(n_295),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_371),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_375),
.B(n_263),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_427),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_327),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_424),
.B(n_388),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_405),
.B(n_253),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_427),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_427),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_407),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_458),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_448),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_448),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

OAI22xp33_ASAP7_75t_L g497 ( 
.A1(n_450),
.A2(n_388),
.B1(n_393),
.B2(n_389),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_452),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_452),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_401),
.B(n_386),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_367),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_452),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_452),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_452),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_415),
.B(n_389),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_469),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_419),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_446),
.B(n_387),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_469),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_401),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_393),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_457),
.B(n_382),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_471),
.B(n_461),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_402),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_425),
.B(n_383),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_429),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_421),
.B(n_383),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_421),
.B(n_385),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_421),
.A2(n_240),
.B1(n_196),
.B2(n_193),
.Y(n_533)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_445),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_458),
.Y(n_535)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_464),
.B(n_342),
.C(n_339),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_421),
.A2(n_309),
.B1(n_211),
.B2(n_228),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_447),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_465),
.A2(n_303),
.B1(n_233),
.B2(n_234),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_451),
.B(n_351),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_438),
.B(n_385),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_438),
.B(n_377),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_324),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_406),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_408),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_408),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_408),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_462),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_451),
.B(n_352),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_472),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_418),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_472),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_409),
.A2(n_347),
.B1(n_376),
.B2(n_384),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_440),
.B(n_391),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_451),
.B(n_356),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_423),
.B(n_392),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_423),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_418),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_428),
.B(n_357),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_436),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_445),
.B(n_263),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_428),
.B(n_392),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_410),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_433),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_438),
.B(n_185),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_403),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_438),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_400),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_409),
.A2(n_296),
.B1(n_237),
.B2(n_239),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_410),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_437),
.B(n_358),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_439),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_439),
.Y(n_594)
);

AOI21x1_ASAP7_75t_L g595 ( 
.A1(n_400),
.A2(n_361),
.B(n_359),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_441),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_454),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_467),
.B(n_160),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_440),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_459),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_404),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_404),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_411),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_465),
.B(n_368),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_411),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_465),
.B(n_373),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_410),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_412),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_467),
.A2(n_290),
.B1(n_244),
.B2(n_250),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_412),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_410),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_468),
.B(n_251),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_422),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_422),
.Y(n_622)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_599),
.B(n_442),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_474),
.B(n_463),
.C(n_460),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_573),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_586),
.B(n_468),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_468),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_519),
.B(n_468),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_477),
.A2(n_442),
.B1(n_459),
.B2(n_443),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_477),
.B(n_443),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_573),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_508),
.B(n_416),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_477),
.B(n_443),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_503),
.B(n_418),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_515),
.A2(n_276),
.B1(n_275),
.B2(n_272),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_573),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_526),
.B(n_416),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_534),
.B(n_443),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_528),
.B(n_417),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_482),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_502),
.B(n_417),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_536),
.B(n_255),
.C(n_254),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_503),
.B(n_418),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_502),
.B(n_418),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_582),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_503),
.B(n_444),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_497),
.B(n_306),
.C(n_299),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_579),
.A2(n_459),
.B1(n_456),
.B2(n_444),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_502),
.A2(n_459),
.B1(n_208),
.B2(n_320),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_535),
.B(n_456),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_495),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_503),
.B(n_269),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_520),
.A2(n_410),
.B(n_287),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_578),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_535),
.B(n_379),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_546),
.B(n_257),
.C(n_256),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_579),
.A2(n_459),
.B1(n_306),
.B2(n_310),
.Y(n_659)
);

AND2x6_ASAP7_75t_SL g660 ( 
.A(n_510),
.B(n_299),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_502),
.B(n_459),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_513),
.B(n_414),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_551),
.B(n_459),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_242),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_501),
.B(n_420),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_578),
.B(n_261),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_482),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_605),
.B(n_380),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_610),
.B(n_265),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_476),
.B(n_268),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_552),
.B(n_434),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_610),
.B(n_294),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_549),
.B(n_269),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_482),
.B(n_287),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_583),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_482),
.B(n_302),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_579),
.A2(n_302),
.B1(n_320),
.B2(n_313),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_605),
.B(n_278),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_546),
.A2(n_310),
.B1(n_311),
.B2(n_314),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_565),
.B(n_313),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_489),
.B(n_381),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_571),
.B(n_311),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_394),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_583),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_591),
.B(n_314),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_545),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_483),
.B(n_520),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_593),
.B(n_395),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_483),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_579),
.A2(n_184),
.B1(n_319),
.B2(n_198),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_593),
.B(n_397),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_594),
.B(n_286),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_596),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_483),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_578),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_594),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_483),
.B(n_258),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_483),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_570),
.B(n_297),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_483),
.B(n_258),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_578),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_612),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_612),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_488),
.B(n_300),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_301),
.Y(n_709)
);

NAND2x1_ASAP7_75t_L g710 ( 
.A(n_490),
.B(n_277),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_533),
.B(n_162),
.Y(n_711)
);

BUFx6f_ASAP7_75t_SL g712 ( 
.A(n_579),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_569),
.B(n_305),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_597),
.B(n_307),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_545),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_598),
.B(n_312),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_522),
.B(n_277),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_598),
.B(n_167),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_533),
.A2(n_174),
.B1(n_298),
.B2(n_289),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_600),
.B(n_169),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_563),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_579),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_563),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_540),
.B(n_170),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_R g725 ( 
.A(n_511),
.B(n_171),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_540),
.B(n_176),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_537),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_620),
.B(n_584),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_530),
.B(n_0),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_600),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_601),
.B(n_177),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_601),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_602),
.B(n_179),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_531),
.B(n_2),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_550),
.B(n_2),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_615),
.B(n_4),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_579),
.A2(n_277),
.B1(n_308),
.B2(n_186),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_537),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_602),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_603),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_522),
.B(n_277),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_5),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_603),
.B(n_181),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_190),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_523),
.B(n_277),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_616),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_566),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_523),
.B(n_277),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_524),
.B(n_5),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_604),
.A2(n_288),
.B1(n_285),
.B2(n_284),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_524),
.B(n_277),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_616),
.B(n_7),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_490),
.B(n_277),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_619),
.B(n_7),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_478),
.B(n_277),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_621),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_566),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_478),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_490),
.B(n_191),
.Y(n_760)
);

INVxp33_ASAP7_75t_L g761 ( 
.A(n_592),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_580),
.B(n_192),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_621),
.B(n_8),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_490),
.B(n_194),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_507),
.B(n_8),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_622),
.B(n_525),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_525),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_589),
.B(n_197),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_529),
.B(n_538),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_537),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_529),
.Y(n_771)
);

OR2x6_ASAP7_75t_SL g772 ( 
.A(n_538),
.B(n_283),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_542),
.A2(n_280),
.B(n_271),
.C(n_270),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_542),
.A2(n_267),
.B1(n_266),
.B2(n_264),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_507),
.B(n_9),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_543),
.B(n_259),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_543),
.B(n_252),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_547),
.B(n_248),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_548),
.B(n_247),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_585),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_521),
.Y(n_781)
);

NOR2x1p5_ASAP7_75t_L g782 ( 
.A(n_478),
.B(n_245),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_507),
.B(n_9),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_507),
.B(n_243),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_646),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_655),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_652),
.B(n_478),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_647),
.B(n_498),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_647),
.A2(n_498),
.B1(n_504),
.B2(n_558),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_629),
.A2(n_498),
.B1(n_504),
.B2(n_558),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_548),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_662),
.Y(n_792)
);

INVx5_ASAP7_75t_L g793 ( 
.A(n_627),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_655),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_768),
.A2(n_504),
.B1(n_498),
.B2(n_564),
.Y(n_795)
);

NAND2x1p5_ASAP7_75t_L g796 ( 
.A(n_722),
.B(n_606),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_656),
.B(n_699),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_678),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_688),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_627),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_633),
.B(n_555),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_700),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_631),
.A2(n_634),
.B1(n_672),
.B2(n_719),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_672),
.B(n_703),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_730),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_719),
.A2(n_564),
.B1(n_568),
.B2(n_614),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_761),
.B(n_568),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_673),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_683),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_690),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_735),
.B(n_486),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_638),
.B(n_504),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_697),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_653),
.A2(n_671),
.B1(n_648),
.B2(n_706),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_665),
.B(n_473),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_653),
.A2(n_480),
.B1(n_475),
.B2(n_481),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_685),
.B(n_588),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_732),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_735),
.B(n_486),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_641),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_739),
.B(n_486),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_740),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_656),
.B(n_505),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_746),
.B(n_754),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_682),
.A2(n_713),
.B1(n_736),
.B2(n_658),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_767),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_707),
.B(n_505),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_705),
.B(n_505),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_715),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_638),
.B(n_588),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_771),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_473),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_640),
.B(n_642),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_757),
.B(n_506),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_721),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_682),
.A2(n_607),
.B1(n_617),
.B2(n_614),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_657),
.B(n_506),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_641),
.B(n_475),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_668),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_641),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_668),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_639),
.B(n_506),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_769),
.B(n_480),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_671),
.B(n_481),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_692),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_641),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_651),
.B(n_606),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_669),
.B(n_607),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_675),
.B(n_608),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_651),
.B(n_608),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_695),
.Y(n_853)
);

AO22x1_ASAP7_75t_L g854 ( 
.A1(n_624),
.A2(n_606),
.B1(n_213),
.B2(n_212),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_670),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_689),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_623),
.B(n_606),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_711),
.A2(n_609),
.B1(n_617),
.B2(n_611),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_766),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_742),
.B(n_609),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_723),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_747),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_782),
.B(n_606),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_670),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_725),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_674),
.B(n_479),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_758),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_670),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_626),
.B(n_611),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_728),
.B(n_479),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_763),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_625),
.B(n_606),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_708),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_670),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_484),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_628),
.B(n_499),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_725),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_632),
.B(n_637),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_752),
.B(n_755),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_664),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_693),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_693),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_693),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_R g884 ( 
.A(n_712),
.B(n_595),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_780),
.Y(n_885)
);

CKINVDCx16_ASAP7_75t_R g886 ( 
.A(n_772),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_752),
.B(n_499),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_781),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_660),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_755),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_693),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_724),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_643),
.B(n_484),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_759),
.B(n_514),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_663),
.B(n_485),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_759),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_744),
.B(n_485),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_681),
.B(n_487),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_726),
.B(n_514),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_661),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_702),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_729),
.B(n_487),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_749),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_649),
.B(n_517),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_636),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_702),
.Y(n_906)
);

NOR2x1_ASAP7_75t_R g907 ( 
.A(n_666),
.B(n_199),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_681),
.B(n_517),
.Y(n_908)
);

AND3x1_ASAP7_75t_L g909 ( 
.A(n_729),
.B(n_518),
.C(n_613),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_712),
.B(n_491),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_649),
.B(n_491),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_630),
.B(n_492),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_702),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_734),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_749),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_676),
.B(n_492),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_696),
.B(n_709),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_714),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_716),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_734),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_686),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_737),
.A2(n_493),
.B1(n_494),
.B2(n_496),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_717),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_765),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_718),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_691),
.A2(n_493),
.B(n_516),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_684),
.B(n_494),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_762),
.B(n_496),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_717),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_694),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_774),
.B(n_500),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_750),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_702),
.B(n_650),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_720),
.B(n_500),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_691),
.A2(n_509),
.B(n_516),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_765),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_774),
.B(n_509),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_727),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_775),
.B(n_512),
.Y(n_939)
);

INVxp67_ASAP7_75t_SL g940 ( 
.A(n_727),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_512),
.Y(n_941)
);

NOR2x1p5_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_518),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_727),
.B(n_518),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_727),
.B(n_518),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_737),
.A2(n_553),
.B1(n_556),
.B2(n_521),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_783),
.B(n_532),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_680),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_659),
.A2(n_553),
.B1(n_532),
.B2(n_554),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_738),
.B(n_527),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_733),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_783),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_743),
.B(n_738),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_645),
.A2(n_618),
.B1(n_613),
.B2(n_527),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_644),
.B(n_554),
.Y(n_954)
);

AND2x6_ASAP7_75t_L g955 ( 
.A(n_738),
.B(n_556),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_741),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_741),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_745),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_738),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_770),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_644),
.B(n_557),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_745),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_748),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_770),
.B(n_537),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_770),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_794),
.B(n_595),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_813),
.B(n_770),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_791),
.A2(n_667),
.B(n_698),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_791),
.A2(n_635),
.B(n_764),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_804),
.Y(n_970)
);

CKINVDCx6p67_ASAP7_75t_R g971 ( 
.A(n_786),
.Y(n_971)
);

CKINVDCx6p67_ASAP7_75t_R g972 ( 
.A(n_815),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_843),
.B(n_951),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_849),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_785),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_809),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_805),
.A2(n_659),
.B1(n_679),
.B2(n_677),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_843),
.B(n_677),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_834),
.B(n_776),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_879),
.A2(n_779),
.B1(n_778),
.B2(n_777),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_921),
.B(n_679),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_925),
.B(n_760),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_793),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_792),
.B(n_557),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_798),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_811),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_914),
.B(n_773),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_792),
.B(n_760),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_SL g990 ( 
.A(n_905),
.B(n_784),
.C(n_764),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_932),
.B(n_784),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_873),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_804),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_804),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_801),
.A2(n_635),
.B(n_751),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_879),
.A2(n_751),
.B(n_748),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_801),
.A2(n_753),
.B(n_756),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_816),
.B(n_753),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_930),
.B(n_710),
.Y(n_999)
);

BUFx8_ASAP7_75t_L g1000 ( 
.A(n_889),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_924),
.B(n_537),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_946),
.A2(n_654),
.B(n_704),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_847),
.B(n_559),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_946),
.A2(n_704),
.B(n_701),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_853),
.B(n_561),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_799),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_955),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_886),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_827),
.A2(n_701),
.B1(n_559),
.B2(n_561),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_793),
.B(n_527),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_918),
.B(n_527),
.Y(n_1011)
);

AO21x2_ASAP7_75t_L g1012 ( 
.A1(n_939),
.A2(n_562),
.B(n_618),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_939),
.A2(n_613),
.B(n_590),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_856),
.B(n_562),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_813),
.B(n_567),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_865),
.B(n_613),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_955),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_952),
.A2(n_590),
.B(n_541),
.C(n_560),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_936),
.B(n_537),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_837),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_920),
.B(n_590),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_890),
.A2(n_590),
.B(n_574),
.C(n_560),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_SL g1024 ( 
.A(n_817),
.B(n_919),
.C(n_915),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_903),
.A2(n_574),
.B(n_560),
.C(n_541),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_941),
.A2(n_541),
.B(n_574),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_802),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_820),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_947),
.A2(n_544),
.B1(n_581),
.B2(n_203),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_810),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_941),
.A2(n_581),
.B(n_544),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_835),
.B(n_544),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_877),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_813),
.B(n_587),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_871),
.A2(n_226),
.B1(n_206),
.B2(n_207),
.C(n_210),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_859),
.B(n_544),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_810),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_835),
.A2(n_581),
.B(n_544),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_826),
.A2(n_581),
.B1(n_544),
.B2(n_219),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_950),
.B(n_581),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_841),
.B(n_14),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_917),
.B(n_581),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_908),
.A2(n_887),
.B(n_845),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_887),
.A2(n_587),
.B(n_575),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_824),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_826),
.A2(n_204),
.B(n_215),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_845),
.A2(n_587),
.B(n_575),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_803),
.A2(n_238),
.B1(n_236),
.B2(n_225),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_885),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_808),
.B(n_892),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_821),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_819),
.B(n_14),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_793),
.B(n_587),
.Y(n_1054)
);

AND2x6_ASAP7_75t_L g1055 ( 
.A(n_933),
.B(n_60),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_846),
.A2(n_575),
.B1(n_567),
.B2(n_18),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_860),
.A2(n_575),
.B(n_567),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_866),
.B(n_15),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_849),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_928),
.A2(n_567),
.B(n_56),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_810),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_954),
.A2(n_149),
.B(n_148),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_880),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_899),
.A2(n_16),
.B(n_21),
.C(n_25),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_861),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_934),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_828),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_829),
.B(n_32),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_926),
.A2(n_935),
.B(n_961),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_833),
.B(n_34),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_938),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_787),
.B(n_795),
.C(n_807),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_814),
.A2(n_38),
.B(n_42),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_909),
.A2(n_854),
.B1(n_850),
.B2(n_851),
.C(n_898),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_823),
.A2(n_43),
.B(n_44),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_862),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_867),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_900),
.B(n_43),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_888),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_900),
.B(n_875),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_875),
.B(n_44),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_933),
.A2(n_50),
.B1(n_52),
.B2(n_61),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_SL g1083 ( 
.A1(n_893),
.A2(n_52),
.B1(n_65),
.B2(n_68),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_832),
.B(n_852),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_821),
.B(n_85),
.Y(n_1085)
);

OAI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_904),
.A2(n_100),
.B1(n_113),
.B2(n_124),
.Y(n_1086)
);

AND2x2_ASAP7_75t_SL g1087 ( 
.A(n_910),
.B(n_127),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_876),
.A2(n_138),
.B1(n_147),
.B2(n_869),
.C(n_893),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_923),
.A2(n_958),
.B(n_956),
.C(n_963),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_855),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_896),
.B(n_907),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_844),
.B(n_876),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_961),
.A2(n_916),
.B(n_964),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_878),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_844),
.B(n_838),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_929),
.A2(n_962),
.B(n_957),
.C(n_789),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_878),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_943),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_836),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_916),
.B(n_904),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_836),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_870),
.B(n_788),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_823),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_790),
.A2(n_912),
.B1(n_911),
.B2(n_818),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_793),
.B(n_960),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_901),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_855),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_902),
.A2(n_894),
.B(n_830),
.C(n_927),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_987),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1044),
.A2(n_998),
.B(n_1104),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1051),
.B(n_944),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1073),
.A2(n_894),
.B1(n_937),
.B2(n_931),
.C(n_912),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1092),
.B(n_911),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1093),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_991),
.B(n_842),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1024),
.B(n_842),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_989),
.B(n_949),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_974),
.B(n_842),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_1004),
.B(n_1002),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_1104),
.A2(n_913),
.A3(n_938),
.B(n_965),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_992),
.B(n_858),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1039),
.A2(n_897),
.B(n_895),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1056),
.A2(n_942),
.B1(n_960),
.B2(n_800),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_971),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1084),
.B(n_881),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1103),
.B(n_881),
.Y(n_1126)
);

AO31x2_ASAP7_75t_L g1127 ( 
.A1(n_1100),
.A2(n_981),
.A3(n_1089),
.B(n_995),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_980),
.A2(n_840),
.B(n_940),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1099),
.B(n_864),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_968),
.A2(n_922),
.B(n_953),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_1080),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1073),
.A2(n_839),
.B1(n_797),
.B2(n_825),
.C(n_945),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_986),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_997),
.A2(n_1060),
.B(n_1026),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1096),
.A2(n_1040),
.A3(n_1025),
.B(n_1101),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_983),
.B(n_974),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_985),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1013),
.A2(n_948),
.B(n_949),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1095),
.A2(n_1045),
.B(n_1037),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1040),
.A2(n_965),
.A3(n_884),
.B(n_910),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1007),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1006),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1094),
.A2(n_955),
.A3(n_872),
.B(n_863),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1056),
.A2(n_863),
.B(n_857),
.C(n_959),
.Y(n_1144)
);

AO31x2_ASAP7_75t_L g1145 ( 
.A1(n_1097),
.A2(n_955),
.A3(n_872),
.B(n_864),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1059),
.B(n_960),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_SL g1147 ( 
.A1(n_1070),
.A2(n_944),
.B(n_857),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1075),
.A2(n_848),
.B1(n_906),
.B2(n_891),
.C(n_883),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1027),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1034),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1098),
.B(n_967),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1000),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1019),
.A2(n_796),
.B(n_800),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1048),
.A2(n_800),
.B(n_822),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1108),
.A2(n_822),
.B(n_842),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1062),
.A2(n_822),
.B(n_874),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_996),
.A2(n_822),
.B(n_874),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_855),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_996),
.A2(n_874),
.B(n_868),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1088),
.A2(n_868),
.B(n_882),
.C(n_883),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1075),
.A2(n_882),
.B1(n_883),
.B2(n_891),
.Y(n_1161)
);

NOR4xp25_ASAP7_75t_L g1162 ( 
.A(n_1064),
.B(n_882),
.C(n_891),
.D(n_906),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1043),
.B(n_906),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1057),
.A2(n_1022),
.B(n_1001),
.Y(n_1164)
);

AOI31xp67_ASAP7_75t_L g1165 ( 
.A1(n_1020),
.A2(n_1009),
.A3(n_1082),
.B(n_978),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1087),
.B(n_1074),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_SL g1167 ( 
.A(n_1082),
.B(n_1066),
.C(n_1063),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1072),
.A2(n_1023),
.B(n_990),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1050),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1015),
.A2(n_1105),
.B(n_1005),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1058),
.A2(n_978),
.B1(n_999),
.B2(n_1067),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1009),
.A2(n_1102),
.B(n_1003),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1106),
.A2(n_1065),
.A3(n_977),
.B(n_1014),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1086),
.A2(n_1007),
.B(n_1018),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1083),
.A2(n_1047),
.B(n_1011),
.C(n_988),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1053),
.A2(n_1047),
.B(n_1078),
.Y(n_1176)
);

AO22x2_ASAP7_75t_L g1177 ( 
.A1(n_1076),
.A2(n_1079),
.B1(n_1077),
.B2(n_1029),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1105),
.A2(n_1054),
.B(n_1010),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1007),
.B(n_1018),
.Y(n_1180)
);

AOI22x1_ASAP7_75t_L g1181 ( 
.A1(n_1083),
.A2(n_1010),
.B1(n_1071),
.B2(n_984),
.Y(n_1181)
);

INVx3_ASAP7_75t_SL g1182 ( 
.A(n_1008),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1054),
.A2(n_1071),
.B(n_1081),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1021),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1018),
.A2(n_1012),
.B(n_1041),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1012),
.A2(n_966),
.B(n_982),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1000),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1091),
.A2(n_979),
.B(n_1068),
.C(n_1042),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1049),
.A2(n_1036),
.B1(n_1030),
.B2(n_973),
.C(n_1017),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1085),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_976),
.A2(n_984),
.A3(n_1055),
.B(n_1085),
.Y(n_1191)
);

AND3x2_ASAP7_75t_L g1192 ( 
.A(n_1090),
.B(n_1085),
.C(n_1055),
.Y(n_1192)
);

AOI21xp33_ASAP7_75t_L g1193 ( 
.A1(n_967),
.A2(n_1035),
.B(n_1016),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1055),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1055),
.A2(n_1035),
.B(n_1016),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_970),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1016),
.A2(n_1035),
.B(n_993),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_970),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_993),
.A2(n_994),
.B(n_1031),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_993),
.B(n_994),
.Y(n_1200)
);

AO32x2_ASAP7_75t_L g1201 ( 
.A1(n_1107),
.A2(n_994),
.A3(n_1031),
.B1(n_1038),
.B2(n_1061),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1031),
.B(n_1038),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1107),
.Y(n_1203)
);

AOI221x1_ASAP7_75t_L g1204 ( 
.A1(n_1038),
.A2(n_1075),
.B1(n_1073),
.B2(n_1064),
.C(n_879),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1061),
.B(n_1107),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1061),
.A2(n_1104),
.A3(n_1100),
.B(n_1044),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1051),
.B(n_805),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_991),
.B(n_510),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1024),
.B(n_510),
.C(n_951),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_992),
.B(n_805),
.Y(n_1210)
);

AO21x2_ASAP7_75t_L g1211 ( 
.A1(n_1012),
.A2(n_1044),
.B(n_969),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_975),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1007),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_992),
.B(n_805),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_SL g1215 ( 
.A(n_1007),
.B(n_815),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1073),
.A2(n_1092),
.B(n_879),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1051),
.B(n_805),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_998),
.A2(n_879),
.B(n_477),
.C(n_920),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1104),
.A2(n_1100),
.A3(n_1044),
.B(n_1093),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1093),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1051),
.B(n_805),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1051),
.B(n_805),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_975),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_972),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_975),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_992),
.B(n_805),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_992),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1093),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1007),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1093),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1069),
.A2(n_1044),
.B(n_969),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_975),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_992),
.B(n_805),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1093),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1044),
.A2(n_879),
.B(n_477),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1044),
.A2(n_879),
.B(n_1092),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_972),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1044),
.A2(n_879),
.B(n_1092),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1051),
.B(n_805),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_967),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1044),
.A2(n_879),
.B(n_1092),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1051),
.B(n_805),
.Y(n_1242)
);

O2A1O1Ixp5_ASAP7_75t_SL g1243 ( 
.A1(n_1033),
.A2(n_1020),
.B(n_1001),
.C(n_1073),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1024),
.B(n_510),
.C(n_951),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1007),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_972),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_990),
.A2(n_920),
.B1(n_890),
.B2(n_879),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1044),
.A2(n_879),
.B(n_1092),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1104),
.A2(n_1100),
.A3(n_1044),
.B(n_1093),
.Y(n_1249)
);

CKINVDCx8_ASAP7_75t_R g1250 ( 
.A(n_1008),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1085),
.B(n_967),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1206),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1171),
.B(n_1175),
.C(n_1110),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1230),
.A2(n_1234),
.B(n_1134),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1109),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1171),
.A2(n_1218),
.B1(n_1208),
.B2(n_1110),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1235),
.A2(n_1238),
.B(n_1236),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1177),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_L g1260 ( 
.A(n_1141),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1235),
.A2(n_1248),
.B(n_1241),
.Y(n_1261)
);

AOI221xp5_ASAP7_75t_L g1262 ( 
.A1(n_1167),
.A2(n_1247),
.B1(n_1166),
.B2(n_1176),
.C(n_1216),
.Y(n_1262)
);

NAND2x1_ASAP7_75t_L g1263 ( 
.A(n_1229),
.B(n_1215),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1112),
.A2(n_1139),
.B(n_1164),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1122),
.A2(n_1170),
.B(n_1185),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1117),
.B(n_1221),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1183),
.A2(n_1174),
.B(n_1231),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1222),
.B(n_1239),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1204),
.A2(n_1123),
.A3(n_1160),
.B(n_1113),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1242),
.A2(n_1247),
.B1(n_1227),
.B2(n_1189),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1161),
.A2(n_1130),
.B(n_1186),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1112),
.A2(n_1130),
.B(n_1132),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1152),
.A2(n_1187),
.B1(n_1190),
.B2(n_1124),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1136),
.B(n_1111),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1206),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1210),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1150),
.Y(n_1277)
);

CKINVDCx8_ASAP7_75t_R g1278 ( 
.A(n_1151),
.Y(n_1278)
);

NOR2xp67_ASAP7_75t_SL g1279 ( 
.A(n_1250),
.B(n_1224),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1161),
.A2(n_1188),
.B1(n_1233),
.B2(n_1226),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1214),
.B(n_1131),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1125),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1176),
.A2(n_1121),
.B1(n_1123),
.B2(n_1251),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1251),
.A2(n_1137),
.B1(n_1181),
.B2(n_1169),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1132),
.A2(n_1157),
.B(n_1159),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1201),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1186),
.A2(n_1162),
.B(n_1168),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1162),
.A2(n_1211),
.B(n_1159),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1195),
.B(n_1251),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1144),
.A2(n_1116),
.B1(n_1148),
.B2(n_1113),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1195),
.A2(n_1128),
.B(n_1125),
.C(n_1180),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1231),
.A2(n_1119),
.B(n_1243),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1201),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1133),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1209),
.A2(n_1244),
.B(n_1155),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1119),
.A2(n_1156),
.B(n_1154),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1142),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1115),
.B(n_1158),
.C(n_1199),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1182),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1237),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1206),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1151),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1246),
.B(n_1196),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1178),
.Y(n_1304)
);

AOI222xp33_ASAP7_75t_L g1305 ( 
.A1(n_1149),
.A2(n_1223),
.B1(n_1225),
.B2(n_1232),
.C1(n_1212),
.C2(n_1184),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1147),
.A2(n_1153),
.B(n_1179),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1194),
.B(n_1197),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1173),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1173),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1126),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1126),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1163),
.A2(n_1202),
.B(n_1200),
.C(n_1129),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1201),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1129),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1163),
.A2(n_1193),
.B(n_1199),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1172),
.A2(n_1192),
.B1(n_1138),
.B2(n_1193),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1138),
.A2(n_1229),
.B(n_1172),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1198),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1203),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1246),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1200),
.B(n_1202),
.C(n_1205),
.Y(n_1321)
);

NAND2xp33_ASAP7_75t_SL g1322 ( 
.A(n_1141),
.B(n_1245),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1165),
.A2(n_1240),
.B1(n_1146),
.B2(n_1118),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1140),
.A2(n_1120),
.B(n_1191),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1120),
.A2(n_1127),
.A3(n_1249),
.B(n_1219),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1219),
.A2(n_1249),
.B(n_1120),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1140),
.A2(n_1191),
.B(n_1135),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1240),
.B(n_1191),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1127),
.A2(n_1249),
.A3(n_1219),
.B(n_1135),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1141),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1135),
.A2(n_1145),
.B(n_1140),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1143),
.B(n_1213),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1145),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1145),
.A2(n_1220),
.B(n_1114),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1143),
.B(n_1024),
.C(n_951),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1143),
.B(n_1195),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1218),
.A2(n_879),
.B(n_477),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1190),
.A2(n_1123),
.A3(n_1104),
.B1(n_1067),
.B2(n_981),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1240),
.B(n_1007),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1251),
.B(n_1195),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1185),
.A2(n_1139),
.B(n_1134),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_1152),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1114),
.A2(n_1228),
.B(n_1220),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1109),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1177),
.Y(n_1346)
);

OAI221xp5_ASAP7_75t_L g1347 ( 
.A1(n_1218),
.A2(n_827),
.B1(n_1171),
.B2(n_624),
.C(n_1024),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1195),
.B(n_1251),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1218),
.A2(n_879),
.B(n_477),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1114),
.A2(n_1228),
.B(n_1220),
.Y(n_1350)
);

OAI21xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1110),
.A2(n_879),
.B(n_477),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_SL g1352 ( 
.A1(n_1218),
.A2(n_879),
.B(n_1235),
.C(n_1110),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1109),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_1208),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1218),
.A2(n_879),
.B(n_477),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1195),
.B(n_1251),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1206),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1206),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1166),
.B(n_951),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1109),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1167),
.A2(n_477),
.B1(n_1166),
.B2(n_827),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1171),
.A2(n_951),
.B1(n_879),
.B2(n_477),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1114),
.A2(n_1228),
.B(n_1220),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1207),
.B(n_1217),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1204),
.A2(n_1185),
.A3(n_1139),
.B(n_1218),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1117),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1171),
.A2(n_951),
.B1(n_879),
.B2(n_477),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_SL g1369 ( 
.A(n_1152),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1250),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1218),
.A2(n_879),
.B(n_477),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1209),
.B(n_865),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1177),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1224),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1171),
.A2(n_1082),
.B1(n_951),
.B2(n_879),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1167),
.A2(n_477),
.B1(n_1166),
.B2(n_827),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1292),
.A2(n_1255),
.B(n_1258),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1359),
.A2(n_1347),
.B1(n_1343),
.B2(n_1257),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1370),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1277),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1375),
.B(n_1276),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1351),
.A2(n_1376),
.B(n_1349),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1274),
.Y(n_1384)
);

BUFx4f_ASAP7_75t_L g1385 ( 
.A(n_1320),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1292),
.A2(n_1255),
.B(n_1350),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1337),
.A2(n_1371),
.B(n_1355),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1363),
.A2(n_1368),
.B(n_1376),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1352),
.A2(n_1253),
.B(n_1261),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1270),
.A2(n_1359),
.B(n_1352),
.C(n_1377),
.Y(n_1391)
);

O2A1O1Ixp5_ASAP7_75t_L g1392 ( 
.A1(n_1291),
.A2(n_1295),
.B(n_1290),
.C(n_1335),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1362),
.A2(n_1377),
.B(n_1262),
.C(n_1280),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1291),
.A2(n_1342),
.B(n_1272),
.Y(n_1394)
);

AOI221x1_ASAP7_75t_SL g1395 ( 
.A1(n_1254),
.A2(n_1361),
.B1(n_1341),
.B2(n_1268),
.C(n_1365),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1256),
.B(n_1345),
.Y(n_1396)
);

OA22x2_ASAP7_75t_L g1397 ( 
.A1(n_1340),
.A2(n_1304),
.B1(n_1281),
.B2(n_1289),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1370),
.Y(n_1398)
);

CKINVDCx6p67_ASAP7_75t_R g1399 ( 
.A(n_1369),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1343),
.Y(n_1400)
);

AND2x2_ASAP7_75t_SL g1401 ( 
.A(n_1286),
.B(n_1293),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1362),
.A2(n_1283),
.B1(n_1353),
.B2(n_1360),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1326),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1252),
.A2(n_1358),
.B(n_1275),
.C(n_1301),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1289),
.B(n_1348),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1283),
.A2(n_1372),
.B1(n_1272),
.B2(n_1284),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1275),
.A2(n_1357),
.B(n_1282),
.C(n_1263),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1354),
.B(n_1367),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1302),
.B(n_1354),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1342),
.A2(n_1272),
.B(n_1264),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1294),
.B(n_1297),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1305),
.B(n_1318),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1284),
.A2(n_1299),
.B1(n_1300),
.B2(n_1374),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1319),
.B(n_1313),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1287),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1320),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1299),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1300),
.A2(n_1303),
.B1(n_1298),
.B2(n_1323),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1312),
.A2(n_1310),
.B(n_1311),
.C(n_1314),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1259),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_1369),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1346),
.B(n_1373),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1323),
.A2(n_1278),
.B1(n_1340),
.B2(n_1273),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1321),
.B(n_1269),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1330),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1338),
.A2(n_1316),
.B(n_1348),
.C(n_1356),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1269),
.B(n_1330),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1269),
.B(n_1312),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1269),
.B(n_1315),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1315),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1338),
.A2(n_1287),
.B(n_1271),
.C(n_1285),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1315),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1338),
.A2(n_1271),
.B(n_1285),
.C(n_1288),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1260),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1307),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1338),
.B(n_1288),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1329),
.B(n_1325),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1260),
.A2(n_1316),
.B1(n_1339),
.B2(n_1307),
.Y(n_1438)
);

AND2x2_ASAP7_75t_SL g1439 ( 
.A(n_1336),
.B(n_1328),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1307),
.B(n_1332),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1264),
.A2(n_1296),
.B(n_1267),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_SL g1442 ( 
.A1(n_1328),
.A2(n_1264),
.B(n_1336),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1339),
.A2(n_1333),
.B(n_1327),
.C(n_1309),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1329),
.B(n_1325),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1265),
.A2(n_1344),
.B(n_1334),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1333),
.A2(n_1344),
.B1(n_1279),
.B2(n_1308),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1366),
.B(n_1327),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1366),
.B(n_1322),
.Y(n_1448)
);

BUFx8_ASAP7_75t_L g1449 ( 
.A(n_1306),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1324),
.A2(n_1331),
.B1(n_1317),
.B2(n_1334),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1364),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1266),
.B(n_1274),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1292),
.A2(n_1255),
.B(n_1258),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1289),
.B(n_1348),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1292),
.A2(n_1255),
.B(n_1350),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1276),
.B(n_1281),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1363),
.A2(n_1368),
.B(n_1347),
.C(n_1257),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1276),
.B(n_1281),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1313),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1320),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1375),
.B(n_1276),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1410),
.A2(n_1429),
.B(n_1394),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1441),
.A2(n_1424),
.B(n_1445),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1420),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1449),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1401),
.B(n_1436),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1417),
.B(n_1400),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1452),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1388),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1457),
.B(n_1459),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1460),
.B(n_1414),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1395),
.B(n_1384),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_1408),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1460),
.B(n_1422),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1408),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1449),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1458),
.A2(n_1391),
.B1(n_1393),
.B2(n_1383),
.C(n_1379),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1411),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1427),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1396),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_SL g1482 ( 
.A(n_1380),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1403),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1402),
.A2(n_1423),
.B1(n_1406),
.B2(n_1453),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1382),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1398),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1381),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1430),
.A2(n_1432),
.B(n_1451),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1448),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1426),
.B(n_1428),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1435),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1437),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1444),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1426),
.B(n_1439),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1419),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1415),
.A2(n_1390),
.B(n_1392),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1409),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1407),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1407),
.Y(n_1500)
);

INVxp67_ASAP7_75t_R g1501 ( 
.A(n_1418),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1446),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1431),
.A2(n_1433),
.B(n_1387),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1440),
.B(n_1439),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1433),
.A2(n_1443),
.B(n_1447),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1450),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1425),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1404),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1463),
.B(n_1378),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1378),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1378),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1467),
.B(n_1454),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1489),
.B(n_1412),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1467),
.B(n_1454),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1458),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1478),
.A2(n_1389),
.B1(n_1393),
.B2(n_1413),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1484),
.A2(n_1397),
.B1(n_1391),
.B2(n_1399),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1483),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1466),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1506),
.B(n_1456),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1506),
.B(n_1464),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1466),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1475),
.B(n_1386),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1477),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1497),
.B(n_1386),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1461),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1488),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1397),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1469),
.B(n_1405),
.Y(n_1530)
);

AND2x2_ASAP7_75t_SL g1531 ( 
.A(n_1494),
.B(n_1455),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1392),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1484),
.A2(n_1438),
.B1(n_1421),
.B2(n_1434),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1508),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1485),
.B(n_1442),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1519),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1518),
.A2(n_1494),
.B1(n_1503),
.B2(n_1490),
.Y(n_1537)
);

OAI33xp33_ASAP7_75t_L g1538 ( 
.A1(n_1513),
.A2(n_1510),
.A3(n_1529),
.B1(n_1524),
.B2(n_1479),
.B3(n_1471),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1519),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1535),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1520),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1516),
.A2(n_1501),
.B1(n_1495),
.B2(n_1496),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1471),
.Y(n_1543)
);

AOI31xp33_ASAP7_75t_L g1544 ( 
.A1(n_1532),
.A2(n_1507),
.A3(n_1476),
.B(n_1468),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1519),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1521),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1516),
.A2(n_1501),
.B1(n_1495),
.B2(n_1496),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1532),
.B(n_1522),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1512),
.B(n_1481),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1510),
.B(n_1475),
.Y(n_1550)
);

AOI221xp5_ASAP7_75t_L g1551 ( 
.A1(n_1532),
.A2(n_1502),
.B1(n_1503),
.B2(n_1508),
.C(n_1500),
.Y(n_1551)
);

AOI211xp5_ASAP7_75t_L g1552 ( 
.A1(n_1515),
.A2(n_1522),
.B(n_1509),
.C(n_1511),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1470),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_SL g1554 ( 
.A(n_1520),
.B(n_1486),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1518),
.A2(n_1477),
.B1(n_1480),
.B2(n_1491),
.C(n_1500),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_SL g1556 ( 
.A(n_1533),
.B(n_1499),
.C(n_1487),
.Y(n_1556)
);

OAI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1533),
.A2(n_1480),
.B1(n_1491),
.B2(n_1499),
.C(n_1465),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1533),
.A2(n_1465),
.B1(n_1492),
.B2(n_1493),
.C(n_1479),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1515),
.A2(n_1503),
.B1(n_1505),
.B2(n_1504),
.Y(n_1559)
);

AND2x4_ASAP7_75t_SL g1560 ( 
.A(n_1530),
.B(n_1498),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1512),
.B(n_1514),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1551),
.A2(n_1526),
.B(n_1528),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1559),
.A2(n_1526),
.B(n_1528),
.Y(n_1563)
);

INVx4_ASAP7_75t_SL g1564 ( 
.A(n_1541),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1552),
.B(n_1522),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1559),
.A2(n_1517),
.B(n_1528),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_SL g1568 ( 
.A(n_1537),
.B(n_1547),
.C(n_1542),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1536),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

INVxp33_ASAP7_75t_L g1573 ( 
.A(n_1554),
.Y(n_1573)
);

BUFx8_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1548),
.B(n_1522),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1550),
.B(n_1524),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1578)
);

AO21x1_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1534),
.B(n_1511),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1557),
.B(n_1509),
.C(n_1511),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1540),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1546),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1564),
.B(n_1560),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1573),
.B(n_1482),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1573),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_SL g1587 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1564),
.B(n_1560),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1564),
.B(n_1509),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1569),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1567),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1564),
.B(n_1549),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1569),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1574),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1564),
.B(n_1509),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1564),
.B(n_1511),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1549),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1581),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1520),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1568),
.B(n_1523),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1543),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1570),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1570),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1565),
.C(n_1562),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1567),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1570),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

AND2x2_ASAP7_75t_SL g1617 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1571),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1579),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1579),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1568),
.Y(n_1623)
);

NAND4xp25_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1525),
.C(n_1527),
.D(n_1555),
.Y(n_1624)
);

NOR2xp67_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1556),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1582),
.A2(n_1534),
.B(n_1527),
.C(n_1558),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1623),
.B(n_1579),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1575),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1597),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1577),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1582),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1619),
.B(n_1612),
.Y(n_1632)
);

NAND2x2_ASAP7_75t_L g1633 ( 
.A(n_1587),
.B(n_1525),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1619),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1585),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1592),
.B(n_1575),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1595),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1599),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1625),
.B(n_1579),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

AO22x1_ASAP7_75t_L g1642 ( 
.A1(n_1621),
.A2(n_1574),
.B1(n_1525),
.B2(n_1568),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1576),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1595),
.B(n_1578),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1609),
.B(n_1576),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1595),
.B(n_1385),
.Y(n_1646)
);

NOR3xp33_ASAP7_75t_L g1647 ( 
.A(n_1612),
.B(n_1538),
.C(n_1583),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1626),
.B(n_1525),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1625),
.A2(n_1617),
.B(n_1624),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1602),
.B(n_1574),
.Y(n_1650)
);

NAND4xp25_ASAP7_75t_L g1651 ( 
.A(n_1590),
.B(n_1596),
.C(n_1605),
.D(n_1589),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1606),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1606),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1608),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1584),
.B(n_1578),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1584),
.B(n_1578),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1608),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1590),
.B(n_1571),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1588),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1610),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1661)
);

NAND2x1_ASAP7_75t_L g1662 ( 
.A(n_1588),
.B(n_1583),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1636),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1635),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1647),
.A2(n_1617),
.B1(n_1591),
.B2(n_1614),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1629),
.B(n_1605),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1662),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1634),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1646),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1659),
.Y(n_1671)
);

INVx3_ASAP7_75t_SL g1672 ( 
.A(n_1631),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1627),
.B(n_1609),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1639),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1628),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1646),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_1589),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1653),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1631),
.B(n_1655),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1641),
.B(n_1603),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1640),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1640),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1656),
.B(n_1601),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1664),
.A2(n_1627),
.B1(n_1649),
.B2(n_1633),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1665),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1665),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1671),
.B(n_1647),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1669),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1666),
.A2(n_1649),
.B1(n_1642),
.B2(n_1591),
.C(n_1614),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1674),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1664),
.A2(n_1617),
.B1(n_1648),
.B2(n_1600),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1682),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1684),
.A2(n_1562),
.B1(n_1563),
.B2(n_1650),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1674),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1672),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1673),
.A2(n_1651),
.B(n_1562),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1675),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1672),
.A2(n_1600),
.B1(n_1598),
.B2(n_1589),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1672),
.A2(n_1600),
.B1(n_1598),
.B2(n_1589),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1668),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1692),
.B(n_1682),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1693),
.A2(n_1686),
.B1(n_1562),
.B2(n_1673),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1699),
.B(n_1677),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1699),
.B(n_1677),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1702),
.B(n_1668),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1704),
.B(n_1670),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1690),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1708),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1708),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1694),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1710),
.A2(n_1703),
.B(n_1696),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1715),
.A2(n_1700),
.B1(n_1689),
.B2(n_1698),
.C(n_1691),
.Y(n_1721)
);

NAND4xp25_ASAP7_75t_L g1722 ( 
.A(n_1709),
.B(n_1670),
.C(n_1668),
.D(n_1707),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1645),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1713),
.A2(n_1670),
.B(n_1695),
.C(n_1697),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1713),
.A2(n_1676),
.B(n_1701),
.Y(n_1725)
);

AOI221x1_ASAP7_75t_L g1726 ( 
.A1(n_1714),
.A2(n_1670),
.B1(n_1687),
.B2(n_1678),
.C(n_1685),
.Y(n_1726)
);

INVxp33_ASAP7_75t_L g1727 ( 
.A(n_1709),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1717),
.A2(n_1687),
.B1(n_1681),
.B2(n_1685),
.C(n_1706),
.Y(n_1728)
);

OAI21xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1711),
.A2(n_1680),
.B(n_1688),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1727),
.B(n_1711),
.Y(n_1730)
);

OAI32xp33_ASAP7_75t_L g1731 ( 
.A1(n_1729),
.A2(n_1718),
.A3(n_1719),
.B1(n_1712),
.B2(n_1681),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1723),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1726),
.Y(n_1733)
);

AOI211xp5_ASAP7_75t_L g1734 ( 
.A1(n_1720),
.A2(n_1718),
.B(n_1705),
.C(n_1679),
.Y(n_1734)
);

OAI21xp33_ASAP7_75t_L g1735 ( 
.A1(n_1721),
.A2(n_1667),
.B(n_1680),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1733),
.B(n_1724),
.C(n_1722),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1730),
.B(n_1732),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1734),
.B(n_1688),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1731),
.B(n_1725),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1735),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1732),
.B(n_1728),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1730),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1737),
.Y(n_1743)
);

AND3x4_ASAP7_75t_L g1744 ( 
.A(n_1740),
.B(n_1679),
.C(n_1416),
.Y(n_1744)
);

XNOR2xp5_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1679),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_L g1746 ( 
.A(n_1741),
.B(n_1679),
.C(n_1658),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1739),
.B(n_1598),
.C(n_1600),
.D(n_1661),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1745),
.A2(n_1736),
.B(n_1742),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1743),
.B(n_1421),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1746),
.A2(n_1385),
.B(n_1660),
.C(n_1598),
.Y(n_1750)
);

NAND4xp25_ASAP7_75t_L g1751 ( 
.A(n_1748),
.B(n_1747),
.C(n_1744),
.D(n_1661),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1751),
.B(n_1750),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1752),
.Y(n_1753)
);

XNOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1752),
.B(n_1749),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1658),
.B1(n_1643),
.B2(n_1637),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1755),
.A2(n_1611),
.B1(n_1618),
.B2(n_1616),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1756),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1758),
.Y(n_1759)
);

XNOR2xp5_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1601),
.Y(n_1760)
);

AO21x1_ASAP7_75t_L g1761 ( 
.A1(n_1759),
.A2(n_1611),
.B(n_1618),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1761),
.B(n_1760),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1616),
.B1(n_1615),
.B2(n_1610),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1615),
.B1(n_1604),
.B2(n_1603),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1622),
.B(n_1620),
.C(n_1613),
.Y(n_1765)
);


endmodule