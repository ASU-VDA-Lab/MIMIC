module fake_netlist_6_4227_n_96 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_96);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_96;

wire n_52;
wire n_91;
wire n_46;
wire n_88;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_92;
wire n_42;
wire n_90;
wire n_54;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_78;
wire n_84;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_55;
wire n_94;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI21x1_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_16),
.B(n_14),
.Y(n_33)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_7),
.B(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx8_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

XNOR2x1_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_1),
.Y(n_43)
);

NOR2x1_ASAP7_75t_L g44 ( 
.A(n_6),
.B(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_6),
.Y(n_46)
);

NOR2xp67_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

AOI221xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.C(n_7),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_2),
.C(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_22),
.C(n_46),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_31),
.C(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_36),
.C(n_34),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_31),
.B(n_41),
.C(n_40),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_33),
.B(n_28),
.C(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_38),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_45),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_47),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AND2x4_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_68),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_78),
.B(n_77),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_35),
.Y(n_86)
);

OAI211xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_44),
.B(n_61),
.C(n_74),
.Y(n_87)
);

OAI221xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_72),
.B1(n_70),
.B2(n_67),
.C(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_85),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_73),
.B1(n_75),
.B2(n_37),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_71),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_94),
.Y(n_96)
);


endmodule