module fake_jpeg_18922_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_58),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_28),
.Y(n_66)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_24),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_26),
.B(n_22),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_40),
.C(n_37),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_76),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_39),
.B1(n_41),
.B2(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_87),
.B1(n_47),
.B2(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_20),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_50),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_86),
.B1(n_57),
.B2(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_82),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_41),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_46),
.C(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_43),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_41),
.B1(n_38),
.B2(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_102),
.B1(n_70),
.B2(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_46),
.Y(n_128)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_27),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_64),
.B1(n_63),
.B2(n_73),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_127),
.B1(n_138),
.B2(n_75),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_65),
.B1(n_69),
.B2(n_72),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_80),
.B(n_69),
.C(n_76),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_100),
.B1(n_28),
.B2(n_21),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_80),
.B1(n_83),
.B2(n_49),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_45),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_84),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_75),
.B1(n_56),
.B2(n_45),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_46),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_97),
.B1(n_103),
.B2(n_107),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_17),
.B(n_30),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_16),
.B(n_22),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_136),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_137),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_111),
.B1(n_109),
.B2(n_75),
.Y(n_138)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_152),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_135),
.B1(n_115),
.B2(n_131),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_90),
.B1(n_84),
.B2(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_124),
.B1(n_132),
.B2(n_121),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_108),
.C(n_45),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_27),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_108),
.C(n_56),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_108),
.C(n_56),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_114),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_133),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_20),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_21),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_100),
.C(n_91),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_29),
.C(n_24),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_122),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_30),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_176),
.B1(n_180),
.B2(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_131),
.B1(n_137),
.B2(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_149),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_124),
.B1(n_121),
.B2(n_126),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_26),
.B1(n_22),
.B2(n_17),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_147),
.C(n_164),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_28),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_197),
.B1(n_198),
.B2(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_200),
.B(n_201),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_142),
.B(n_145),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_208),
.C(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_206),
.B1(n_210),
.B2(n_212),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_209),
.B1(n_211),
.B2(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_163),
.C(n_142),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_154),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_173),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_161),
.B(n_143),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_189),
.B1(n_179),
.B2(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_226),
.B1(n_227),
.B2(n_230),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_183),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_203),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_229),
.C(n_231),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_189),
.B1(n_191),
.B2(n_174),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_174),
.B1(n_190),
.B2(n_184),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_171),
.C(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_172),
.B1(n_157),
.B2(n_167),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_167),
.C(n_140),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_195),
.B1(n_209),
.B2(n_194),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_239),
.B1(n_234),
.B2(n_237),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_202),
.CI(n_201),
.CON(n_237),
.SN(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_212),
.B1(n_214),
.B2(n_196),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_157),
.B1(n_153),
.B2(n_29),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_29),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_245),
.Y(n_251)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_221),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_29),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_255),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_245),
.C(n_243),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_218),
.C(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_229),
.B1(n_219),
.B2(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_256),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_8),
.B1(n_1),
.B2(n_3),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_235),
.C(n_240),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_261),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_10),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_235),
.C(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_264),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_10),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_10),
.B(n_4),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_15),
.B(n_5),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_251),
.C(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_9),
.C(n_4),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_11),
.C(n_5),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_6),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_258),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_278)
);

XOR2x1_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_6),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_7),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_7),
.B(n_12),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_15),
.C(n_7),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_278),
.C(n_277),
.Y(n_282)
);

O2A1O1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_13),
.B(n_14),
.C(n_0),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_13),
.Y(n_284)
);


endmodule