module fake_jpeg_30885_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_1),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_2),
.B(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_2),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_22),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_27),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_39),
.B1(n_38),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_15),
.B1(n_25),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_38),
.B1(n_36),
.B2(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_30),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_24),
.B1(n_19),
.B2(n_23),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_70),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_11),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_67),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_10),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_72),
.B1(n_52),
.B2(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_40),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_72),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_45),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_54),
.B1(n_44),
.B2(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_82),
.B1(n_70),
.B2(n_30),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_66),
.B1(n_71),
.B2(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_94),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_79),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_75),
.B1(n_83),
.B2(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_50),
.B(n_44),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_7),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_103),
.C(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_95),
.B1(n_91),
.B2(n_90),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_84),
.B(n_73),
.C(n_74),
.D(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_4),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_99),
.C(n_98),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_109),
.C(n_108),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_43),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_119),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_114),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_112),
.B(n_121),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_124),
.B(n_120),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_113),
.B(n_41),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_41),
.Y(n_126)
);


endmodule