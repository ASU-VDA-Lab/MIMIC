module fake_jpeg_1291_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_42),
.B(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_16),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_16),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_8),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_21),
.C(n_23),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_53),
.C(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_51),
.B1(n_26),
.B2(n_43),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_25),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_19),
.B1(n_32),
.B2(n_33),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_17),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_12),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_94),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_102),
.B(n_40),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_17),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_106),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_9),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_100),
.Y(n_129)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_48),
.B(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_109),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_24),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_108),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_58),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_5),
.B(n_6),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_87),
.B(n_103),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_111),
.Y(n_146)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_55),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_106),
.C(n_95),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_119),
.C(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_85),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_91),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_139),
.C(n_142),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_84),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_99),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_99),
.C(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_112),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_110),
.C(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_157),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_160),
.C(n_161),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_123),
.B1(n_98),
.B2(n_127),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_143),
.B1(n_145),
.B2(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_112),
.B1(n_127),
.B2(n_114),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_145),
.B1(n_118),
.B2(n_113),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_117),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_113),
.C(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_117),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_137),
.C(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_149),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_169),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_105),
.B(n_138),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_121),
.B(n_138),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_163),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_152),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_149),
.C(n_150),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_168),
.B(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_180),
.B1(n_166),
.B2(n_172),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_115),
.B1(n_76),
.B2(n_96),
.Y(n_180)
);

OAI31xp33_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_184),
.A3(n_187),
.B(n_115),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_168),
.B(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_165),
.B(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_189),
.B(n_191),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_171),
.B(n_63),
.Y(n_189)
);

OR2x6_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_8),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_96),
.A3(n_80),
.B1(n_76),
.B2(n_41),
.C1(n_115),
.C2(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_80),
.A3(n_12),
.B1(n_14),
.B2(n_7),
.C1(n_74),
.C2(n_66),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_190),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_196),
.B1(n_193),
.B2(n_74),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_69),
.Y(n_199)
);


endmodule