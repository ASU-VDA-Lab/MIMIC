module fake_jpeg_29820_n_55 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_29),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_23),
.B1(n_21),
.B2(n_5),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_24),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_6),
.C(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_36),
.C(n_7),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_8),
.C(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_47),
.B1(n_39),
.B2(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_43),
.C(n_8),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_31),
.CI(n_34),
.CON(n_55),
.SN(n_55)
);


endmodule