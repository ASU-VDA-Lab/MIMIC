module fake_netlist_1_9155_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
BUFx6f_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_5), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
AOI21xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_0), .B(n_1), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_9), .B(n_0), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_3), .B(n_4), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
XNOR2x2_ASAP7_75t_SL g18 ( .A(n_16), .B(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx4_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
NAND2x1p5_ASAP7_75t_L g21 ( .A(n_19), .B(n_9), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_10), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
XNOR2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_18), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_20), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_21), .B1(n_9), .B2(n_8), .Y(n_27) );
endmodule