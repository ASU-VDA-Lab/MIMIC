module fake_jpeg_2079_n_191 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_191);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_47),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_0),
.Y(n_87)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_67),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_61),
.B1(n_50),
.B2(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_65),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.C(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_86),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_54),
.Y(n_98)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_61),
.B(n_49),
.C(n_56),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_80),
.B1(n_77),
.B2(n_84),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_123),
.B1(n_4),
.B2(n_5),
.Y(n_139)
);

OA22x2_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_61),
.B1(n_60),
.B2(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_60),
.B(n_71),
.C(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_50),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_64),
.C(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_58),
.B1(n_55),
.B2(n_52),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_48),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_102),
.B1(n_103),
.B2(n_60),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_21),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_142),
.B(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_46),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_34),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_116),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_116),
.C(n_32),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_153),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_24),
.C(n_23),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_12),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_4),
.B(n_6),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_9),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_161),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_133),
.CI(n_127),
.CON(n_158),
.SN(n_158)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_140),
.A3(n_134),
.B1(n_143),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_7),
.B(n_8),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_166),
.Y(n_173)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_167),
.B1(n_161),
.B2(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_10),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_171),
.B(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_154),
.C(n_168),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_151),
.B1(n_145),
.B2(n_158),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_146),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_152),
.Y(n_178)
);

XOR2x1_ASAP7_75t_SL g180 ( 
.A(n_178),
.B(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_180),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_178),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_177),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_179),
.B(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_15),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_16),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_17),
.C(n_18),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_18),
.Y(n_191)
);


endmodule