module fake_jpeg_23020_n_63 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx2_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_0),
.B(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_15),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_15),
.B(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_34),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_14),
.B(n_13),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.C(n_12),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_21),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_22),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_48),
.B1(n_37),
.B2(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_22),
.B1(n_24),
.B2(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_47),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_51),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_46),
.B(n_49),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_38),
.C(n_24),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_50),
.A3(n_38),
.B1(n_24),
.B2(n_18),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_16),
.B(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_61),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_6),
.Y(n_63)
);


endmodule