module real_jpeg_23874_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_2),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_104),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_2),
.B(n_50),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_5),
.B(n_47),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_5),
.B(n_85),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_6),
.B(n_47),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_6),
.B(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_6),
.B(n_50),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_6),
.B(n_85),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_29),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_6),
.B(n_25),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_6),
.B(n_34),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_8),
.B(n_25),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_8),
.B(n_85),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_8),
.B(n_50),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_8),
.Y(n_263)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_9),
.B(n_10),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_10),
.B(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_10),
.B(n_47),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_10),
.B(n_85),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_10),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_10),
.B(n_38),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_10),
.B(n_29),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_10),
.B(n_25),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_85),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_11),
.B(n_50),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_11),
.B(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_11),
.B(n_47),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_11),
.B(n_38),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_11),
.B(n_29),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_11),
.B(n_34),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_47),
.Y(n_177)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_12),
.B(n_85),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_12),
.B(n_25),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_13),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_13),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_13),
.B(n_50),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_47),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_13),
.B(n_38),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_13),
.B(n_29),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_15),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_15),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_157),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_15),
.B(n_85),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_15),
.B(n_50),
.Y(n_272)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_29),
.Y(n_72)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_17),
.Y(n_148)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_17),
.Y(n_194)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_17),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.C(n_52),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_119),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_64),
.Y(n_63)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.CI(n_32),
.CON(n_23),
.SN(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_26),
.B(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.C(n_39),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_33),
.B(n_97),
.Y(n_96)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_34),
.Y(n_249)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_41),
.B(n_52),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.C(n_49),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_43),
.B(n_46),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_59),
.C(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_44),
.A2(n_49),
.B1(n_60),
.B2(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_45),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_46),
.B(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_82),
.B1(n_83),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_49),
.B(n_80),
.C(n_83),
.Y(n_117)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_50),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_112),
.C(n_118),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_76),
.A2(n_77),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_96),
.C(n_98),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_78),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_88),
.C(n_92),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_79),
.B(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_101),
.C(n_106),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_83),
.A2(n_87),
.B1(n_101),
.B2(n_102),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_84),
.B(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_88),
.B(n_92),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_88)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_331),
.SN(n_331)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_92),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.CI(n_95),
.CON(n_92),
.SN(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.C(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_368),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_96),
.Y(n_368)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.C(n_111),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_100),
.B(n_355),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_101),
.A2(n_102),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_101),
.B(n_309),
.C(n_310),
.Y(n_330)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_106),
.B(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_341),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_111),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_111),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_111),
.B(n_337),
.C(n_340),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_112),
.B(n_118),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_117),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_113),
.A2(n_114),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_116),
.B(n_117),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_369),
.C(n_370),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_357),
.C(n_358),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_345),
.C(n_346),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_321),
.C(n_322),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_290),
.C(n_291),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_255),
.C(n_256),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_224),
.C(n_225),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_199),
.C(n_200),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_159),
.C(n_170),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_143),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_131),
.B(n_138),
.C(n_143),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_139),
.B(n_141),
.C(n_142),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_144),
.B(n_152),
.C(n_153),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_158),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_158),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_169),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_195),
.C(n_196),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.C(n_185),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.C(n_190),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_213),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_214),
.C(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_207),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_209),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.CI(n_212),
.CON(n_209),
.SN(n_209)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_221),
.B2(n_222),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_240),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.C(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_236),
.C(n_239),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_231),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.CI(n_234),
.CON(n_231),
.SN(n_231)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_247),
.C(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_247),
.B1(n_253),
.B2(n_254),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_280),
.C(n_281),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_251),
.C(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_276),
.B2(n_289),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_277),
.C(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_261),
.C(n_269),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_269),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_265),
.C(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_275),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_317),
.C(n_318),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.CI(n_288),
.CON(n_282),
.SN(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_319),
.B2(n_320),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_292),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_311),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_311),
.C(n_319),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_302),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_303),
.C(n_304),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_298),
.C(n_300),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_310),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_325),
.C(n_344),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_332),
.B2(n_344),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_335),
.C(n_336),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_343),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_340),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_356),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_350),
.C(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_353),
.C(n_354),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_361),
.C(n_366),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_365),
.B2(n_366),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_371),
.Y(n_372)
);


endmodule