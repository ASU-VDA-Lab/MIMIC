module fake_jpeg_6291_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_51;
wire n_245;
wire n_47;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_247;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_212;
wire n_240;
wire n_56;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_273;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_22),
.B1(n_19),
.B2(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_51),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_29),
.B(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_65),
.B1(n_68),
.B2(n_16),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_25),
.C(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_16),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_22),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_29),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_43),
.B1(n_29),
.B2(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_74),
.B1(n_77),
.B2(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_21),
.B1(n_26),
.B2(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_82),
.B1(n_31),
.B2(n_24),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_30),
.B1(n_24),
.B2(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_87),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_32),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_32),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_101),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_58),
.C(n_46),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_98),
.B(n_99),
.CI(n_115),
.CON(n_144),
.SN(n_144)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_31),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_84),
.B1(n_91),
.B2(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_76),
.B1(n_93),
.B2(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_109),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_106),
.B(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_117),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_53),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_63),
.B1(n_59),
.B2(n_50),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_116),
.B1(n_74),
.B2(n_94),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_53),
.C(n_64),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_50),
.B1(n_34),
.B2(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_127),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_149),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_117),
.B(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_142),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_105),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_73),
.B1(n_76),
.B2(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_96),
.B(n_93),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_76),
.B1(n_85),
.B2(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_108),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_157),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_134),
.B(n_113),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_98),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_166),
.C(n_167),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_104),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_110),
.B1(n_130),
.B2(n_128),
.Y(n_182)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_170),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_125),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_119),
.C(n_115),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_119),
.C(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_78),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_174),
.Y(n_196)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_124),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_125),
.B(n_113),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_132),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_138),
.B(n_103),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_181),
.A2(n_186),
.B(n_199),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_156),
.B1(n_174),
.B2(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_124),
.B1(n_149),
.B2(n_136),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_191),
.B1(n_203),
.B2(n_175),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_144),
.C(n_134),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_192),
.C(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_147),
.B1(n_144),
.B2(n_101),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_144),
.C(n_147),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_101),
.B1(n_92),
.B2(n_120),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_198),
.B1(n_163),
.B2(n_161),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_122),
.C(n_78),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_92),
.B1(n_122),
.B2(n_80),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_135),
.B(n_92),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_180),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_32),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_164),
.C(n_176),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_140),
.B1(n_35),
.B2(n_37),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_206),
.B1(n_223),
.B2(n_226),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_177),
.B1(n_173),
.B2(n_155),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_150),
.B(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_214),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_173),
.B(n_150),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_168),
.C(n_165),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_227),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_151),
.B1(n_165),
.B2(n_140),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_172),
.B(n_160),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_189),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_197),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_197),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_201),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_245),
.C(n_246),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_20),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_20),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_226),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_64),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_254),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_263),
.B1(n_256),
.B2(n_262),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_224),
.B(n_214),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_262),
.B(n_263),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_217),
.B1(n_222),
.B2(n_209),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_244),
.A2(n_205),
.B1(n_206),
.B2(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_223),
.B(n_241),
.C(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_233),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_259),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_219),
.B(n_223),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_233),
.A2(n_221),
.B(n_1),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_235),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_11),
.B(n_15),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_237),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_133),
.C(n_140),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_256),
.B(n_251),
.C(n_2),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_56),
.C(n_47),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_12),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_279),
.B(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_71),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_268),
.B(n_271),
.Y(n_283)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_278),
.A3(n_270),
.B1(n_275),
.B2(n_269),
.C1(n_280),
.C2(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_270),
.A3(n_40),
.B1(n_56),
.B2(n_47),
.C1(n_10),
.C2(n_15),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_279),
.A2(n_14),
.A3(n_13),
.B1(n_10),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_3),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_286),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_292),
.B(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_5),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_284),
.C(n_285),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_5),
.B(n_6),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_5),
.B1(n_6),
.B2(n_247),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_5),
.B(n_6),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_298),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_294),
.Y(n_302)
);


endmodule