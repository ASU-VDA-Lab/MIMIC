module fake_netlist_1_6264_n_10 (n_3, n_1, n_2, n_0, n_10);
input n_3;
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_8;
wire n_7;
AND2x2_ASAP7_75t_L g4 ( .A(n_3), .B(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_2), .B(n_1), .Y(n_5) );
AND2x2_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
NOR2x1_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
AOI22xp5_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_4), .B1(n_0), .B2(n_2), .Y(n_8) );
NAND4xp25_ASAP7_75t_L g9 ( .A(n_8), .B(n_7), .C(n_0), .D(n_3), .Y(n_9) );
OAI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_1), .B1(n_3), .B2(n_8), .Y(n_10) );
endmodule