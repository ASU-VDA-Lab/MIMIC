module fake_netlist_5_1822_n_2829 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2829);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2829;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1547;
wire n_1070;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_1276;
wire n_702;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_1644;
wire n_762;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_703;
wire n_698;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

BUFx10_ASAP7_75t_L g615 ( 
.A(n_142),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_167),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_453),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_457),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_117),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_259),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_195),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_226),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_55),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_48),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_81),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_218),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_115),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_484),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_570),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_5),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_34),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_117),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_122),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_519),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_465),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_591),
.B(n_396),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_407),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_196),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_524),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_207),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_483),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_269),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_438),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_276),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_383),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_316),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_595),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_464),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_274),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_360),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_173),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_43),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_590),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_270),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_541),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_97),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_126),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_2),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_476),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_372),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_511),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_391),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_339),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_463),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_357),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_280),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_61),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_314),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_212),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_413),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_512),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_36),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_157),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_257),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_364),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_533),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_507),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_397),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_532),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_459),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_293),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_504),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_509),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_382),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_458),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_306),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_614),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_74),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_549),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_94),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_304),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_441),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_130),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_280),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_110),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_170),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_361),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_592),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_52),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_83),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_471),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_352),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_501),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_76),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_279),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_472),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_212),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_284),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_156),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_345),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_89),
.Y(n_714)
);

BUFx5_ASAP7_75t_L g715 ( 
.A(n_121),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_410),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_26),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_85),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_293),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_163),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_98),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_189),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_252),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_114),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_350),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_115),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_587),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_432),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_4),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_276),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_84),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_69),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_385),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_77),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_33),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_247),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_107),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_489),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_560),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_309),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_564),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_356),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_466),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_302),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_266),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_409),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_285),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_424),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_300),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_184),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_450),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_73),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_410),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_294),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_439),
.Y(n_755)
);

BUFx5_ASAP7_75t_L g756 ( 
.A(n_554),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_465),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_387),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_443),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_334),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_586),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_343),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_239),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_361),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_254),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_365),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_597),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_583),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_378),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_19),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_80),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_613),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_299),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_102),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_55),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_581),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_388),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_561),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_126),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_99),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_451),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_147),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_239),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_420),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_454),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_400),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_250),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_456),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_259),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_209),
.Y(n_791)
);

CKINVDCx14_ASAP7_75t_R g792 ( 
.A(n_338),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_226),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_467),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_334),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_73),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_389),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_295),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_461),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_345),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_153),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_285),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_357),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_397),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_573),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_468),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_304),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_70),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_379),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_325),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_455),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_26),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_215),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_469),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_405),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_107),
.Y(n_816)
);

CKINVDCx14_ASAP7_75t_R g817 ( 
.A(n_365),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_91),
.Y(n_818)
);

CKINVDCx16_ASAP7_75t_R g819 ( 
.A(n_490),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_23),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_264),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_326),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_419),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_542),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_548),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_168),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_545),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_563),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_525),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_85),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_64),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_399),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_388),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_544),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_481),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_260),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_531),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_64),
.Y(n_838)
);

CKINVDCx14_ASAP7_75t_R g839 ( 
.A(n_406),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_445),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_192),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_96),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_153),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_282),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_347),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_48),
.Y(n_846)
);

BUFx10_ASAP7_75t_L g847 ( 
.A(n_309),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_231),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_552),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_462),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_487),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_232),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_495),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_198),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_450),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_452),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_555),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_498),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_218),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_121),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_247),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_538),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_270),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_460),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_715),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_624),
.B(n_0),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_715),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_715),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_715),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_622),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_715),
.Y(n_871)
);

INVxp33_ASAP7_75t_L g872 ( 
.A(n_650),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_715),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_715),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_746),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_746),
.Y(n_876)
);

INVxp33_ASAP7_75t_SL g877 ( 
.A(n_626),
.Y(n_877)
);

INVxp33_ASAP7_75t_L g878 ( 
.A(n_713),
.Y(n_878)
);

INVxp33_ASAP7_75t_L g879 ( 
.A(n_760),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_842),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_842),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_696),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_619),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_842),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_619),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_622),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_792),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_619),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_838),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_619),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_792),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_668),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_714),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_718),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_668),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_668),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_850),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_850),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_850),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_615),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_852),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_817),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_615),
.Y(n_906)
);

INVxp33_ASAP7_75t_SL g907 ( 
.A(n_626),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_817),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_852),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_729),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_729),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_839),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_839),
.B(n_1),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_759),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_759),
.Y(n_915)
);

INVxp33_ASAP7_75t_SL g916 ( 
.A(n_627),
.Y(n_916)
);

INVxp33_ASAP7_75t_SL g917 ( 
.A(n_627),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_806),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_816),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_806),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_692),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_816),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_816),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_816),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_647),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_629),
.Y(n_926)
);

INVxp33_ASAP7_75t_L g927 ( 
.A(n_631),
.Y(n_927)
);

INVxp33_ASAP7_75t_L g928 ( 
.A(n_636),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_638),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_692),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_639),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_617),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_652),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_756),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_618),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_653),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_756),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_756),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_654),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_658),
.B(n_0),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_620),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_621),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_649),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_615),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_625),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_679),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_659),
.Y(n_947)
);

INVxp33_ASAP7_75t_SL g948 ( 
.A(n_861),
.Y(n_948)
);

INVxp33_ASAP7_75t_SL g949 ( 
.A(n_861),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_660),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_756),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_679),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_623),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_756),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_623),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_655),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_756),
.Y(n_957)
);

BUFx2_ASAP7_75t_SL g958 ( 
.A(n_827),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_665),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_669),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_827),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_670),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_858),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_616),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_634),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_946),
.B(n_679),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_884),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_867),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_867),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_921),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_819),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_871),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_871),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_934),
.Y(n_975)
);

AND2x6_ASAP7_75t_L g976 ( 
.A(n_934),
.B(n_773),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_937),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_885),
.B(n_635),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_870),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_923),
.B(n_628),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_938),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_884),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_924),
.B(n_628),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_910),
.B(n_798),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_938),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_911),
.B(n_798),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_865),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_868),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_869),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_886),
.Y(n_991)
);

INVx5_ASAP7_75t_L g992 ( 
.A(n_951),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_914),
.B(n_846),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_870),
.B(n_640),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_886),
.B(n_630),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_873),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_958),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_874),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_889),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_915),
.B(n_918),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_951),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_920),
.B(n_846),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_887),
.B(n_709),
.Y(n_1003)
);

INVxp33_ASAP7_75t_SL g1004 ( 
.A(n_894),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_925),
.B(n_856),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_889),
.Y(n_1006)
);

BUFx12f_ASAP7_75t_L g1007 ( 
.A(n_887),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_954),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_954),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_891),
.B(n_893),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_891),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_875),
.B(n_635),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_925),
.B(n_856),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_876),
.B(n_704),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_880),
.B(n_704),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_957),
.B(n_773),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_893),
.B(n_630),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_896),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_957),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_888),
.B(n_824),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_896),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_888),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_964),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_895),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_897),
.B(n_824),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_964),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_897),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_892),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_898),
.B(n_825),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_892),
.B(n_858),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_881),
.B(n_767),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1001),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_974),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_974),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_994),
.B(n_877),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_1001),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_974),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1008),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_978),
.B(n_900),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_967),
.B(n_978),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_988),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1003),
.A2(n_913),
.B1(n_826),
.B2(n_859),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_988),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_988),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1008),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_989),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_1001),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_967),
.B(n_767),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_972),
.A2(n_826),
.B1(n_859),
.B2(n_747),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1008),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_989),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_1024),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_1000),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_989),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_978),
.B(n_904),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

BUFx8_ASAP7_75t_L g1058 ( 
.A(n_1007),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_998),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_998),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_R g1061 ( 
.A(n_1004),
.B(n_932),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_967),
.B(n_905),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_990),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_972),
.B(n_905),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_1001),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_967),
.B(n_882),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1019),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_978),
.B(n_908),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1018),
.B(n_908),
.Y(n_1069)
);

CKINVDCx16_ASAP7_75t_R g1070 ( 
.A(n_1007),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_1005),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_998),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1018),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1018),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1019),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1019),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1023),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_990),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_990),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1020),
.B(n_877),
.Y(n_1080)
);

NOR2x1_ASAP7_75t_L g1081 ( 
.A(n_995),
.B(n_673),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1023),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1005),
.B(n_899),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1012),
.B(n_901),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1023),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_969),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_977),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_969),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_977),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_969),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_977),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1012),
.B(n_902),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_1007),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1012),
.B(n_909),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_976),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_973),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_990),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_973),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_973),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_973),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1013),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1013),
.B(n_943),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_995),
.B(n_912),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_977),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1022),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_982),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1031),
.A2(n_747),
.B1(n_916),
.B2(n_907),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_982),
.Y(n_1109)
);

CKINVDCx8_ASAP7_75t_R g1110 ( 
.A(n_997),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1000),
.B(n_943),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_982),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_980),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_982),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_980),
.B(n_912),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1017),
.A2(n_837),
.B(n_828),
.Y(n_1116)
);

AND3x2_ASAP7_75t_L g1117 ( 
.A(n_1028),
.B(n_637),
.C(n_644),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_968),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_999),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_SL g1120 ( 
.A(n_1028),
.B(n_965),
.C(n_935),
.Y(n_1120)
);

AND2x6_ASAP7_75t_L g1121 ( 
.A(n_1012),
.B(n_828),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_985),
.B(n_956),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1113),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1041),
.B(n_990),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1041),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1034),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1041),
.B(n_990),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1034),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1041),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1073),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1065),
.B(n_996),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1103),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1035),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1053),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1073),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1035),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1103),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1074),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1049),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1074),
.Y(n_1140)
);

AND3x2_ASAP7_75t_L g1141 ( 
.A(n_1036),
.B(n_823),
.C(n_903),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_1080),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1122),
.B(n_958),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1065),
.B(n_996),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_1043),
.B(n_837),
.Y(n_1145)
);

NOR2x1p5_ASAP7_75t_L g1146 ( 
.A(n_1120),
.B(n_1022),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1113),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1033),
.B(n_996),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1062),
.A2(n_1022),
.B1(n_1017),
.B2(n_1025),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1071),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1066),
.Y(n_1151)
);

CKINVDCx14_ASAP7_75t_R g1152 ( 
.A(n_1106),
.Y(n_1152)
);

NOR2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1106),
.B(n_932),
.Y(n_1153)
);

NOR2x1p5_ASAP7_75t_L g1154 ( 
.A(n_1104),
.B(n_935),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1111),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1064),
.B(n_907),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_1033),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1066),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1065),
.B(n_996),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1122),
.B(n_878),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1111),
.B(n_879),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1033),
.B(n_996),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1038),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1038),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1039),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1039),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1033),
.B(n_996),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_1116),
.A2(n_738),
.B(n_706),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1102),
.B(n_941),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1046),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1054),
.B(n_941),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1066),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1043),
.B(n_1068),
.C(n_945),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1115),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1054),
.B(n_1083),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1046),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1037),
.B(n_1025),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1051),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1118),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1051),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1067),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1037),
.B(n_1030),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_L g1184 ( 
.A(n_1049),
.B(n_773),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_SL g1185 ( 
.A(n_1084),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1049),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1037),
.B(n_981),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1067),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_1081),
.B(n_945),
.C(n_942),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1118),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1066),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1083),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1040),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1040),
.Y(n_1194)
);

INVx8_ASAP7_75t_L g1195 ( 
.A(n_1049),
.Y(n_1195)
);

INVxp33_ASAP7_75t_SL g1196 ( 
.A(n_1108),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1048),
.B(n_981),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1049),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1048),
.B(n_773),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1075),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1048),
.B(n_829),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1075),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1048),
.B(n_829),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1056),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1056),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1076),
.Y(n_1206)
);

INVx8_ASAP7_75t_L g1207 ( 
.A(n_1049),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1049),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1084),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1084),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1114),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_L g1212 ( 
.A(n_1121),
.B(n_1081),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1084),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1092),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1114),
.B(n_829),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1114),
.B(n_829),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1076),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1092),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1077),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1092),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1077),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1092),
.B(n_1095),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1095),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1063),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1095),
.Y(n_1225)
);

CKINVDCx6p67_ASAP7_75t_R g1226 ( 
.A(n_1070),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1069),
.B(n_916),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1110),
.B(n_942),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1095),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1114),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1087),
.B(n_984),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1082),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1082),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1096),
.B(n_1119),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1121),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1087),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1096),
.B(n_1119),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1117),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1050),
.B(n_966),
.C(n_984),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1085),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1085),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1058),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1089),
.B(n_966),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1042),
.Y(n_1244)
);

INVx8_ASAP7_75t_L g1245 ( 
.A(n_1121),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1089),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1091),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1121),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1091),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1042),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1105),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1044),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1105),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1044),
.Y(n_1254)
);

BUFx4f_ASAP7_75t_L g1255 ( 
.A(n_1121),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1110),
.B(n_883),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1096),
.B(n_777),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1045),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1045),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1109),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1108),
.A2(n_849),
.B1(n_862),
.B2(n_930),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1125),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1161),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1227),
.B(n_961),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1129),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_1189),
.B(n_890),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1236),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1160),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1246),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1143),
.B(n_1175),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1247),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1249),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1244),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1157),
.B(n_1047),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1251),
.Y(n_1275)
);

XNOR2x2_ASAP7_75t_L g1276 ( 
.A(n_1261),
.B(n_1050),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1253),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1244),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1260),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1250),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1157),
.B(n_1047),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1157),
.B(n_1070),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1177),
.A2(n_1101),
.B(n_1100),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1226),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1235),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1130),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1226),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1173),
.B(n_906),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1132),
.B(n_985),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1227),
.B(n_963),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1169),
.B(n_1093),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1138),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1179),
.B(n_1052),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1140),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1171),
.B(n_1093),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1147),
.Y(n_1297)
);

INVxp33_ASAP7_75t_L g1298 ( 
.A(n_1134),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1151),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1183),
.A2(n_1116),
.B(n_1055),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1150),
.B(n_944),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_R g1302 ( 
.A(n_1196),
.B(n_917),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1158),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1196),
.B(n_917),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1158),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1152),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1250),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1158),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1172),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1195),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1172),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1155),
.B(n_872),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1172),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1191),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1191),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1191),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1252),
.Y(n_1317)
);

NOR2xp67_ASAP7_75t_L g1318 ( 
.A(n_1239),
.B(n_987),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1252),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1254),
.Y(n_1320)
);

XOR2xp5_ASAP7_75t_L g1321 ( 
.A(n_1152),
.B(n_971),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1254),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1155),
.B(n_987),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1137),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1258),
.Y(n_1325)
);

OR2x2_ASAP7_75t_SL g1326 ( 
.A(n_1145),
.B(n_866),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1258),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1259),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1259),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1180),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1137),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1142),
.B(n_948),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1190),
.Y(n_1333)
);

INVx4_ASAP7_75t_SL g1334 ( 
.A(n_1185),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1230),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1242),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1194),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1194),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1142),
.B(n_948),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1204),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1204),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1240),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1142),
.B(n_949),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1240),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1241),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1241),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_1112),
.B(n_1109),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1187),
.B(n_1052),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1209),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1210),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1126),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1213),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1197),
.A2(n_1059),
.B(n_1055),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1214),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1146),
.B(n_1061),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1218),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1156),
.B(n_949),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_1058),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1228),
.B(n_993),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1223),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1192),
.B(n_993),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1225),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1229),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1174),
.B(n_633),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1222),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1211),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1211),
.Y(n_1367)
);

XOR2xp5_ASAP7_75t_L g1368 ( 
.A(n_1123),
.B(n_1058),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1145),
.B(n_662),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1231),
.A2(n_1060),
.B(n_1059),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1193),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1205),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

XOR2xp5_ASAP7_75t_L g1374 ( 
.A(n_1123),
.B(n_1058),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1126),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1128),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1242),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1128),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1256),
.B(n_1002),
.Y(n_1379)
);

BUFx5_ASAP7_75t_L g1380 ( 
.A(n_1248),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1238),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1154),
.B(n_1243),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1133),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1149),
.B(n_1002),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1133),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1136),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1136),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1141),
.B(n_707),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1153),
.B(n_927),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1186),
.B(n_1096),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_1185),
.Y(n_1391)
);

INVxp67_ASAP7_75t_SL g1392 ( 
.A(n_1124),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1163),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1124),
.B(n_711),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1139),
.B(n_928),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1245),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1139),
.B(n_931),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1163),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1164),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1164),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1165),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1165),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1166),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1166),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1215),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1170),
.B(n_1060),
.Y(n_1406)
);

XOR2xp5_ASAP7_75t_L g1407 ( 
.A(n_1139),
.B(n_642),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1170),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1176),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1176),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1178),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1178),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1224),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1181),
.B(n_1072),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1139),
.B(n_956),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1181),
.B(n_1072),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1182),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1185),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1182),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1188),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1127),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1188),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1200),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1200),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1202),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1198),
.B(n_1014),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1215),
.Y(n_1427)
);

XOR2xp5_ASAP7_75t_L g1428 ( 
.A(n_1198),
.B(n_657),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1216),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1199),
.B(n_804),
.Y(n_1430)
);

XOR2xp5_ASAP7_75t_L g1431 ( 
.A(n_1198),
.B(n_661),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1199),
.B(n_864),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1202),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1206),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1206),
.Y(n_1435)
);

INVxp33_ASAP7_75t_L g1436 ( 
.A(n_1216),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1217),
.B(n_1112),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1217),
.Y(n_1438)
);

OR2x2_ASAP7_75t_SL g1439 ( 
.A(n_1198),
.B(n_866),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1195),
.B(n_940),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1219),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1208),
.B(n_1014),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1208),
.B(n_1014),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1219),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1201),
.B(n_825),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1221),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1221),
.Y(n_1447)
);

AND2x6_ASAP7_75t_L g1448 ( 
.A(n_1208),
.B(n_1063),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1232),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1232),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1233),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1168),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1245),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1186),
.B(n_1096),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1245),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1235),
.B(n_926),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1233),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1168),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1208),
.B(n_1014),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1357),
.B(n_1201),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1357),
.B(n_1203),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_1413),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1312),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_SL g1464 ( 
.A(n_1296),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1319),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1264),
.B(n_1291),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1297),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1270),
.B(n_1186),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1395),
.B(n_1186),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1439),
.A2(n_1255),
.B1(n_1195),
.B2(n_1207),
.Y(n_1470)
);

NAND2xp33_ASAP7_75t_L g1471 ( 
.A(n_1310),
.B(n_1195),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1273),
.Y(n_1472)
);

NAND2xp33_ASAP7_75t_SL g1473 ( 
.A(n_1396),
.B(n_1235),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1278),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1304),
.B(n_1203),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1397),
.B(n_1255),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1263),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1284),
.Y(n_1478)
);

CKINVDCx14_ASAP7_75t_R g1479 ( 
.A(n_1321),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1322),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1304),
.B(n_1148),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1310),
.B(n_1207),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1276),
.A2(n_1121),
.B1(n_1212),
.B2(n_1235),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1394),
.B(n_1131),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1382),
.A2(n_1212),
.B1(n_1121),
.B2(n_1207),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1359),
.B(n_1248),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1325),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1327),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1263),
.A2(n_1207),
.B1(n_1184),
.B2(n_1245),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1280),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1365),
.B(n_1144),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1332),
.B(n_1343),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1334),
.B(n_1234),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1421),
.B(n_1159),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1268),
.A2(n_1184),
.B1(n_1237),
.B2(n_1234),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1268),
.B(n_1248),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1301),
.B(n_940),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1389),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1292),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1364),
.B(n_1015),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1285),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1364),
.B(n_1015),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1339),
.B(n_1162),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1328),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1421),
.B(n_1167),
.Y(n_1505)
);

NAND2xp33_ASAP7_75t_SL g1506 ( 
.A(n_1453),
.B(n_1224),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1323),
.B(n_1224),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1379),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1339),
.B(n_1237),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1324),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1369),
.B(n_1015),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1329),
.Y(n_1512)
);

NOR2xp67_ASAP7_75t_SL g1513 ( 
.A(n_1310),
.B(n_1096),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1369),
.B(n_1015),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1348),
.B(n_1086),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1344),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1298),
.B(n_641),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1345),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1307),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1324),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1317),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1346),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1430),
.A2(n_1257),
.B(n_1032),
.C(n_689),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1330),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1331),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1358),
.A2(n_703),
.B1(n_705),
.B2(n_693),
.C(n_684),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1320),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1287),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1333),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1342),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1334),
.B(n_1257),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1351),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1348),
.B(n_1086),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1331),
.B(n_643),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1294),
.B(n_1088),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1376),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1294),
.B(n_1088),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1430),
.A2(n_1032),
.B1(n_1094),
.B2(n_1090),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1326),
.B(n_929),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1302),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1392),
.B(n_1090),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1392),
.B(n_1094),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1432),
.B(n_936),
.C(n_933),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1337),
.B(n_645),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1334),
.B(n_939),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1455),
.A2(n_676),
.B1(n_680),
.B2(n_663),
.Y(n_1546)
);

BUFx4f_ASAP7_75t_L g1547 ( 
.A(n_1440),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1285),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1384),
.A2(n_1032),
.B1(n_1099),
.B2(n_1097),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1361),
.B(n_1032),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1338),
.B(n_1097),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1371),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1290),
.B(n_616),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1340),
.B(n_1099),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1341),
.B(n_646),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1306),
.B(n_682),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1286),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1289),
.B(n_1100),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1285),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1293),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1372),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1295),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1456),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1419),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1290),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1407),
.B(n_648),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1413),
.A2(n_1078),
.B(n_1063),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1447),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1267),
.B(n_1101),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1418),
.B(n_947),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1269),
.B(n_1107),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1456),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1428),
.B(n_651),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1271),
.B(n_1272),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1391),
.B(n_950),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1275),
.B(n_1107),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1336),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1377),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1277),
.B(n_968),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1318),
.A2(n_632),
.B1(n_672),
.B2(n_671),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1279),
.A2(n_671),
.B1(n_672),
.B2(n_632),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1288),
.B(n_1266),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1375),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1418),
.B(n_959),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1448),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1378),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1388),
.B(n_616),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1274),
.A2(n_1079),
.B(n_1078),
.Y(n_1588)
);

BUFx5_ASAP7_75t_L g1589 ( 
.A(n_1448),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1262),
.B(n_983),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1370),
.B(n_1078),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1383),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1415),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1370),
.B(n_1078),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1385),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1355),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1265),
.B(n_983),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1386),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1282),
.B(n_685),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1349),
.B(n_667),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1431),
.A2(n_1445),
.B1(n_1426),
.B2(n_1443),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1387),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1436),
.B(n_1373),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1368),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1350),
.A2(n_690),
.B1(n_701),
.B2(n_686),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1381),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1440),
.A2(n_677),
.B1(n_688),
.B2(n_675),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1352),
.B(n_656),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1354),
.B(n_1356),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1393),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1360),
.B(n_664),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1448),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1440),
.A2(n_1310),
.B1(n_1363),
.B2(n_1362),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1335),
.B(n_991),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1398),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1442),
.B(n_675),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1299),
.A2(n_1305),
.B1(n_1308),
.B2(n_1303),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1399),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1309),
.B(n_666),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1400),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_L g1621 ( 
.A(n_1380),
.B(n_1079),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1311),
.B(n_1079),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1459),
.B(n_677),
.Y(n_1623)
);

AND2x2_ASAP7_75t_SL g1624 ( 
.A(n_1458),
.B(n_688),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1405),
.A2(n_716),
.B(n_723),
.C(n_721),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1313),
.A2(n_739),
.B1(n_741),
.B2(n_727),
.Y(n_1626)
);

AND2x2_ASAP7_75t_SL g1627 ( 
.A(n_1314),
.B(n_698),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1401),
.Y(n_1628)
);

NOR2xp67_ASAP7_75t_SL g1629 ( 
.A(n_1315),
.B(n_761),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1402),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1316),
.B(n_962),
.C(n_960),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1366),
.B(n_1098),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1367),
.B(n_1098),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1403),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1374),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1353),
.B(n_1098),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1404),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1427),
.A2(n_772),
.B1(n_779),
.B2(n_768),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1353),
.B(n_1098),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1429),
.A2(n_678),
.B1(n_687),
.B2(n_683),
.C(n_674),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1274),
.A2(n_1098),
.B(n_1057),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1408),
.B(n_991),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1409),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_L g1644 ( 
.A(n_1380),
.B(n_805),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1410),
.A2(n_744),
.B1(n_757),
.B2(n_730),
.C(n_724),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1417),
.B(n_691),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1420),
.B(n_1006),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1422),
.B(n_1006),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1423),
.A2(n_835),
.B1(n_851),
.B2(n_834),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1424),
.B(n_1010),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1425),
.B(n_1010),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1433),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1380),
.B(n_853),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1434),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1435),
.B(n_953),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1452),
.B(n_695),
.C(n_694),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1438),
.B(n_857),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_SL g1659 ( 
.A(n_1281),
.B(n_698),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1448),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1441),
.A2(n_774),
.B(n_775),
.C(n_766),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1444),
.B(n_1029),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1446),
.B(n_1029),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1621),
.A2(n_1281),
.B(n_1300),
.Y(n_1664)
);

CKINVDCx11_ASAP7_75t_R g1665 ( 
.A(n_1528),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1586),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1460),
.A2(n_1283),
.B(n_1300),
.C(n_1449),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1461),
.A2(n_1475),
.B(n_1481),
.C(n_1466),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1471),
.A2(n_1283),
.B(n_1390),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1492),
.B(n_1450),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1592),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1601),
.A2(n_1457),
.B1(n_1451),
.B2(n_1406),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1482),
.A2(n_1390),
.B(n_1406),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1503),
.B(n_1414),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1510),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1624),
.B(n_1380),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1595),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1501),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1467),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1501),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1500),
.B(n_1414),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1509),
.A2(n_1416),
.B1(n_1437),
.B2(n_1347),
.Y(n_1682)
);

BUFx4f_ASAP7_75t_L g1683 ( 
.A(n_1577),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1563),
.B(n_1416),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1602),
.Y(n_1685)
);

A2O1A1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1596),
.A2(n_1437),
.B(n_784),
.C(n_789),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1484),
.A2(n_1454),
.B(n_1380),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1644),
.A2(n_1470),
.B(n_1476),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1499),
.B(n_1380),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1582),
.A2(n_794),
.B(n_797),
.C(n_783),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1470),
.A2(n_1448),
.B(n_975),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1612),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1491),
.A2(n_975),
.B(n_979),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1502),
.B(n_801),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1615),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1511),
.B(n_802),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1578),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1515),
.A2(n_979),
.B(n_975),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1514),
.B(n_813),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1507),
.A2(n_1016),
.B(n_976),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1612),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1515),
.A2(n_979),
.B(n_975),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1533),
.A2(n_979),
.B(n_975),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1603),
.A2(n_1657),
.B(n_1608),
.C(n_1611),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1477),
.B(n_667),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1647),
.A2(n_822),
.B(n_830),
.C(n_821),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1498),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1593),
.B(n_841),
.Y(n_1708)
);

BUFx12f_ASAP7_75t_L g1709 ( 
.A(n_1606),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1570),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1533),
.A2(n_986),
.B(n_979),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_R g1712 ( 
.A(n_1479),
.B(n_1464),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1508),
.B(n_845),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1627),
.B(n_667),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1524),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1550),
.B(n_854),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1494),
.B(n_697),
.Y(n_1717)
);

O2A1O1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1640),
.A2(n_740),
.B(n_765),
.C(n_734),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1505),
.B(n_1565),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1535),
.A2(n_986),
.B(n_979),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1618),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1612),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1620),
.Y(n_1723)
);

AO21x1_ASAP7_75t_L g1724 ( 
.A1(n_1613),
.A2(n_740),
.B(n_734),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1628),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1552),
.B(n_953),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1535),
.A2(n_992),
.B(n_986),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1575),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1574),
.B(n_699),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1501),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1539),
.A2(n_778),
.B(n_815),
.C(n_765),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1540),
.B(n_700),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1463),
.B(n_681),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1495),
.A2(n_1016),
.B(n_976),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1609),
.B(n_702),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1566),
.B(n_710),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1529),
.B(n_712),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1557),
.B(n_1560),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1483),
.A2(n_1016),
.B(n_976),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1537),
.A2(n_992),
.B(n_986),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1573),
.A2(n_719),
.B1(n_720),
.B2(n_717),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1537),
.A2(n_992),
.B(n_986),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1562),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1630),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1660),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1654),
.A2(n_992),
.B(n_986),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1625),
.A2(n_815),
.B(n_778),
.C(n_955),
.Y(n_1747)
);

AOI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1659),
.A2(n_1594),
.B(n_1591),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1553),
.A2(n_725),
.B1(n_726),
.B2(n_722),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1587),
.A2(n_955),
.B(n_922),
.C(n_919),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1660),
.Y(n_1751)
);

INVx11_ASAP7_75t_L g1752 ( 
.A(n_1520),
.Y(n_1752)
);

NAND2xp33_ASAP7_75t_L g1753 ( 
.A(n_1589),
.B(n_728),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1591),
.A2(n_1026),
.B(n_1009),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1661),
.A2(n_708),
.B(n_771),
.C(n_681),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1525),
.B(n_731),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_R g1757 ( 
.A(n_1506),
.B(n_470),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1619),
.A2(n_733),
.B(n_736),
.C(n_735),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1583),
.Y(n_1759)
);

AO21x1_ASAP7_75t_L g1760 ( 
.A1(n_1613),
.A2(n_3),
.B(n_2),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1616),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1634),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1547),
.A2(n_737),
.B1(n_742),
.B2(n_732),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1600),
.B(n_681),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1636),
.A2(n_1016),
.B(n_976),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1561),
.B(n_743),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1636),
.A2(n_1016),
.B(n_976),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1637),
.Y(n_1768)
);

CKINVDCx10_ASAP7_75t_R g1769 ( 
.A(n_1616),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1544),
.A2(n_745),
.B1(n_749),
.B2(n_748),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1555),
.A2(n_1534),
.B1(n_1623),
.B2(n_1616),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1485),
.A2(n_750),
.B(n_753),
.C(n_751),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1598),
.Y(n_1773)
);

AO22x1_ASAP7_75t_L g1774 ( 
.A1(n_1545),
.A2(n_752),
.B1(n_755),
.B2(n_754),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1651),
.B(n_758),
.Y(n_1775)
);

OAI321xp33_ASAP7_75t_L g1776 ( 
.A1(n_1526),
.A2(n_812),
.A3(n_771),
.B1(n_847),
.B2(n_781),
.C(n_708),
.Y(n_1776)
);

AO21x1_ASAP7_75t_L g1777 ( 
.A1(n_1496),
.A2(n_4),
.B(n_3),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1623),
.A2(n_762),
.B1(n_764),
.B2(n_763),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1623),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1563),
.B(n_708),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1610),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1643),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1548),
.B(n_999),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1465),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1652),
.B(n_1497),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1563),
.B(n_771),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1559),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1548),
.Y(n_1788)
);

INVxp33_ASAP7_75t_SL g1789 ( 
.A(n_1556),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1639),
.A2(n_1588),
.B(n_1462),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1641),
.A2(n_1009),
.B(n_992),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1559),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1570),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1486),
.A2(n_1009),
.B(n_992),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1584),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1480),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1653),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1572),
.B(n_769),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1517),
.B(n_770),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1487),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1559),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1572),
.B(n_776),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1655),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1541),
.A2(n_1026),
.B(n_1009),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1572),
.B(n_780),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1532),
.Y(n_1806)
);

AO21x1_ASAP7_75t_L g1807 ( 
.A1(n_1607),
.A2(n_6),
.B(n_5),
.Y(n_1807)
);

AO21x1_ASAP7_75t_L g1808 ( 
.A1(n_1607),
.A2(n_1580),
.B(n_1468),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1646),
.B(n_1579),
.Y(n_1809)
);

NOR2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1478),
.B(n_1545),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1656),
.B(n_782),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1488),
.B(n_785),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1584),
.B(n_781),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1546),
.B(n_781),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1541),
.A2(n_1009),
.B(n_1026),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1469),
.A2(n_1016),
.B(n_976),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1542),
.A2(n_1009),
.B(n_1026),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1547),
.B(n_812),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1542),
.A2(n_1016),
.B(n_976),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1567),
.A2(n_1473),
.B(n_1489),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1504),
.B(n_786),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1512),
.B(n_787),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1516),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1518),
.B(n_788),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1493),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1522),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1536),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1631),
.B(n_812),
.Y(n_1828)
);

NOR2xp67_ASAP7_75t_L g1829 ( 
.A(n_1604),
.B(n_1635),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1543),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1564),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1568),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_R g1833 ( 
.A(n_1599),
.B(n_473),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1530),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1590),
.B(n_790),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1617),
.A2(n_793),
.B1(n_795),
.B2(n_791),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1597),
.B(n_796),
.Y(n_1837)
);

AO21x1_ASAP7_75t_L g1838 ( 
.A1(n_1632),
.A2(n_7),
.B(n_6),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1472),
.B(n_799),
.Y(n_1839)
);

BUFx4f_ASAP7_75t_L g1840 ( 
.A(n_1493),
.Y(n_1840)
);

OAI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1543),
.A2(n_807),
.B(n_803),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1474),
.A2(n_1519),
.B1(n_1521),
.B2(n_1490),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1658),
.B(n_847),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1638),
.B(n_800),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1549),
.A2(n_1016),
.B(n_809),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1527),
.B(n_808),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1614),
.B(n_810),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1642),
.B(n_811),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1585),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1642),
.B(n_1648),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1585),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1558),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1569),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1626),
.B(n_847),
.Y(n_1854)
);

AO21x1_ASAP7_75t_L g1855 ( 
.A1(n_1633),
.A2(n_8),
.B(n_7),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1648),
.B(n_814),
.Y(n_1856)
);

NOR3xp33_ASAP7_75t_L g1857 ( 
.A(n_1668),
.B(n_1645),
.C(n_1581),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1793),
.Y(n_1858)
);

NAND2x1_ASAP7_75t_L g1859 ( 
.A(n_1684),
.B(n_1629),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1704),
.A2(n_1581),
.B(n_1523),
.C(n_1649),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1664),
.A2(n_1662),
.B(n_1649),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1799),
.A2(n_1605),
.B1(n_1650),
.B2(n_1531),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1670),
.A2(n_1809),
.B1(n_1771),
.B2(n_1674),
.Y(n_1863)
);

AND2x2_ASAP7_75t_SL g1864 ( 
.A(n_1840),
.B(n_1531),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1785),
.B(n_1551),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1844),
.A2(n_1662),
.B(n_1663),
.C(n_1571),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_R g1867 ( 
.A(n_1697),
.B(n_1589),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1679),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1736),
.B(n_1554),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1738),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1810),
.B(n_1576),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1728),
.B(n_818),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1673),
.A2(n_1669),
.B(n_1850),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1789),
.B(n_820),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1715),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1688),
.A2(n_1622),
.B(n_1538),
.Y(n_1876)
);

AND3x2_ASAP7_75t_L g1877 ( 
.A(n_1814),
.B(n_1622),
.C(n_1589),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1665),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1696),
.B(n_831),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1719),
.B(n_832),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1717),
.B(n_833),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1714),
.A2(n_840),
.B(n_843),
.C(n_836),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1840),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1852),
.B(n_844),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1753),
.A2(n_1513),
.B(n_1589),
.Y(n_1885)
);

O2A1O1Ixp5_ASAP7_75t_L g1886 ( 
.A1(n_1724),
.A2(n_1589),
.B(n_855),
.C(n_860),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1771),
.A2(n_863),
.B1(n_848),
.B2(n_999),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1830),
.B(n_1),
.Y(n_1888)
);

INVx4_ASAP7_75t_L g1889 ( 
.A(n_1752),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1681),
.A2(n_970),
.B(n_1026),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1848),
.B(n_8),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1710),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1856),
.B(n_9),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1854),
.A2(n_999),
.B1(n_1021),
.B2(n_1011),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1820),
.A2(n_1057),
.B(n_970),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1790),
.A2(n_1057),
.B(n_970),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1853),
.B(n_9),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1666),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1676),
.A2(n_1667),
.B(n_1682),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1775),
.B(n_10),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1818),
.A2(n_1011),
.B1(n_1027),
.B2(n_1021),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1755),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1694),
.B(n_11),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1675),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1741),
.B(n_1770),
.C(n_1778),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1699),
.B(n_12),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1732),
.B(n_474),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1825),
.Y(n_1908)
);

AOI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1780),
.A2(n_1011),
.B1(n_1027),
.B2(n_1021),
.Y(n_1909)
);

CKINVDCx10_ASAP7_75t_R g1910 ( 
.A(n_1712),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1687),
.A2(n_970),
.B(n_1011),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1691),
.A2(n_970),
.B(n_1011),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1734),
.A2(n_970),
.B(n_1021),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1786),
.A2(n_1843),
.B1(n_1733),
.B2(n_1764),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1834),
.A2(n_1027),
.B1(n_1021),
.B2(n_15),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1795),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1726),
.B(n_13),
.Y(n_1917)
);

AO21x1_ASAP7_75t_L g1918 ( 
.A1(n_1672),
.A2(n_13),
.B(n_14),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1707),
.B(n_475),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1834),
.A2(n_1027),
.B1(n_16),
.B2(n_14),
.Y(n_1920)
);

A2O1A1Ixp33_ASAP7_75t_L g1921 ( 
.A1(n_1718),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1819),
.A2(n_603),
.B(n_602),
.Y(n_1922)
);

AOI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1748),
.A2(n_478),
.B(n_477),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1708),
.B(n_17),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1678),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1743),
.Y(n_1926)
);

CKINVDCx10_ASAP7_75t_R g1927 ( 
.A(n_1709),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1689),
.A2(n_1684),
.B(n_1765),
.Y(n_1928)
);

OR2x6_ASAP7_75t_L g1929 ( 
.A(n_1825),
.B(n_479),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1678),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1684),
.A2(n_610),
.B(n_609),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1776),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1765),
.A2(n_612),
.B(n_482),
.Y(n_1933)
);

NAND2x1p5_ASAP7_75t_L g1934 ( 
.A(n_1683),
.B(n_1788),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1835),
.B(n_1837),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1726),
.B(n_18),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1683),
.B(n_20),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1678),
.Y(n_1938)
);

NAND2xp33_ASAP7_75t_L g1939 ( 
.A(n_1825),
.B(n_22),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1761),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1847),
.B(n_21),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1769),
.Y(n_1942)
);

O2A1O1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1776),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1943)
);

O2A1O1Ixp5_ASAP7_75t_L g1944 ( 
.A1(n_1808),
.A2(n_27),
.B(n_24),
.C(n_25),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1729),
.B(n_24),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1804),
.A2(n_599),
.B(n_598),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1815),
.A2(n_601),
.B(n_600),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1759),
.Y(n_1948)
);

NOR3xp33_ASAP7_75t_L g1949 ( 
.A(n_1774),
.B(n_25),
.C(n_27),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1735),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1705),
.B(n_28),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1779),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1716),
.B(n_1811),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1758),
.A2(n_1706),
.B(n_1686),
.C(n_1750),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1756),
.B(n_31),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1817),
.A2(n_611),
.B(n_485),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1829),
.B(n_480),
.Y(n_1957)
);

O2A1O1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1772),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1731),
.A2(n_36),
.B(n_32),
.C(n_35),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1773),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1770),
.B(n_35),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1680),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1749),
.B(n_37),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1671),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1781),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1791),
.A2(n_608),
.B(n_488),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1741),
.B(n_1798),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1778),
.B(n_37),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1802),
.B(n_486),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_L g1970 ( 
.A(n_1841),
.B(n_38),
.C(n_39),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1700),
.A2(n_1739),
.B(n_1702),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1749),
.B(n_38),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1813),
.B(n_39),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1769),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1677),
.B(n_40),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1713),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1680),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1805),
.B(n_491),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1685),
.B(n_40),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1754),
.A2(n_493),
.B(n_492),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1680),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1695),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1721),
.B(n_41),
.Y(n_1983)
);

AO32x2_ASAP7_75t_L g1984 ( 
.A1(n_1842),
.A2(n_43),
.A3(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1698),
.A2(n_607),
.B(n_496),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1730),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1723),
.B(n_42),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1725),
.B(n_44),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1744),
.B(n_45),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1782),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1762),
.B(n_45),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1768),
.B(n_46),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1797),
.B(n_46),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1803),
.B(n_47),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1737),
.B(n_47),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1806),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1841),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1692),
.Y(n_1998)
);

O2A1O1Ixp33_ASAP7_75t_L g1999 ( 
.A1(n_1763),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1827),
.B(n_52),
.Y(n_2000)
);

AOI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1703),
.A2(n_497),
.B(n_494),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1828),
.A2(n_1766),
.B1(n_1821),
.B2(n_1812),
.Y(n_2002)
);

AO21x2_ASAP7_75t_L g2003 ( 
.A1(n_1767),
.A2(n_500),
.B(n_499),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1711),
.A2(n_503),
.B(n_502),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1822),
.A2(n_56),
.B1(n_53),
.B2(n_54),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1833),
.B(n_53),
.Y(n_2006)
);

O2A1O1Ixp5_ASAP7_75t_SL g2007 ( 
.A1(n_1784),
.A2(n_57),
.B(n_54),
.C(n_56),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1831),
.B(n_57),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1832),
.B(n_58),
.Y(n_2009)
);

O2A1O1Ixp33_ASAP7_75t_SL g2010 ( 
.A1(n_1796),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1720),
.A2(n_605),
.B(n_506),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1800),
.Y(n_2012)
);

AO22x1_ASAP7_75t_L g2013 ( 
.A1(n_1836),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1823),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1824),
.B(n_62),
.Y(n_2015)
);

AOI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1727),
.A2(n_508),
.B(n_505),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1740),
.A2(n_513),
.B(n_510),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1757),
.B(n_1826),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1839),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_2019)
);

BUFx12f_ASAP7_75t_L g2020 ( 
.A(n_1730),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1742),
.A2(n_604),
.B(n_515),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1746),
.A2(n_594),
.B(n_516),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1730),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1846),
.B(n_63),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1801),
.B(n_65),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1801),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1693),
.A2(n_593),
.B(n_517),
.Y(n_2027)
);

NAND2xp33_ASAP7_75t_L g2028 ( 
.A(n_1787),
.B(n_66),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1787),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1760),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1863),
.B(n_1807),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1898),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1873),
.A2(n_1794),
.B(n_1783),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1883),
.B(n_1692),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1967),
.A2(n_1860),
.B(n_1935),
.Y(n_2035)
);

O2A1O1Ixp5_ASAP7_75t_SL g2036 ( 
.A1(n_1887),
.A2(n_1849),
.B(n_1851),
.C(n_1788),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1890),
.A2(n_1845),
.B(n_1816),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1869),
.B(n_1777),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1885),
.A2(n_1855),
.B(n_1838),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1857),
.A2(n_1747),
.B(n_1690),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1905),
.A2(n_1851),
.B(n_1722),
.Y(n_2041)
);

AO21x2_ASAP7_75t_L g2042 ( 
.A1(n_1861),
.A2(n_1792),
.B(n_1787),
.Y(n_2042)
);

NOR2xp67_ASAP7_75t_L g2043 ( 
.A(n_1899),
.B(n_1701),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1904),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1866),
.A2(n_1751),
.B(n_1745),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1971),
.A2(n_1751),
.B(n_1745),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1930),
.Y(n_2047)
);

NAND2x1p5_ASAP7_75t_L g2048 ( 
.A(n_1925),
.B(n_1792),
.Y(n_2048)
);

INVx3_ASAP7_75t_L g2049 ( 
.A(n_1883),
.Y(n_2049)
);

BUFx12f_ASAP7_75t_L g2050 ( 
.A(n_1878),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1886),
.A2(n_1792),
.B(n_67),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1870),
.B(n_68),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1983),
.B(n_1917),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1940),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1953),
.B(n_69),
.Y(n_2055)
);

NAND2x1_ASAP7_75t_L g2056 ( 
.A(n_1871),
.B(n_514),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1908),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1858),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1865),
.B(n_70),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1895),
.A2(n_520),
.B(n_518),
.Y(n_2060)
);

OAI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1876),
.A2(n_71),
.B(n_72),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1911),
.A2(n_522),
.B(n_521),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1976),
.B(n_71),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_1923),
.A2(n_526),
.B(n_523),
.Y(n_2064)
);

BUFx2_ASAP7_75t_L g2065 ( 
.A(n_2029),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1954),
.A2(n_72),
.B(n_74),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1936),
.B(n_527),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1913),
.A2(n_529),
.B(n_528),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1862),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_2069)
);

OAI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2002),
.A2(n_75),
.B(n_78),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1970),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1930),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_SL g2073 ( 
.A(n_2003),
.B(n_534),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_1912),
.A2(n_2001),
.B(n_1980),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1964),
.B(n_79),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1896),
.A2(n_536),
.B(n_535),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1982),
.B(n_81),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1875),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1996),
.B(n_537),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1968),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2080)
);

OAI21x1_ASAP7_75t_L g2081 ( 
.A1(n_1928),
.A2(n_540),
.B(n_539),
.Y(n_2081)
);

OA22x2_ASAP7_75t_L g2082 ( 
.A1(n_2005),
.A2(n_87),
.B1(n_82),
.B2(n_86),
.Y(n_2082)
);

NOR2x1_ASAP7_75t_SL g2083 ( 
.A(n_2003),
.B(n_543),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_SL g2084 ( 
.A1(n_1932),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1961),
.B(n_88),
.Y(n_2085)
);

AO31x2_ASAP7_75t_L g2086 ( 
.A1(n_1918),
.A2(n_547),
.A3(n_550),
.B(n_546),
.Y(n_2086)
);

NOR2x1_ASAP7_75t_SL g2087 ( 
.A(n_2018),
.B(n_551),
.Y(n_2087)
);

OAI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1958),
.A2(n_90),
.B(n_91),
.Y(n_2088)
);

OAI21x1_ASAP7_75t_L g2089 ( 
.A1(n_1946),
.A2(n_556),
.B(n_553),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1947),
.A2(n_558),
.B(n_557),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1926),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1930),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1963),
.B(n_90),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_2020),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_SL g2095 ( 
.A1(n_1999),
.A2(n_92),
.B(n_93),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1944),
.A2(n_92),
.B(n_93),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1922),
.A2(n_562),
.B(n_559),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_1938),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1921),
.A2(n_94),
.B(n_95),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1972),
.B(n_95),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1948),
.Y(n_2101)
);

AO21x2_ASAP7_75t_L g2102 ( 
.A1(n_1933),
.A2(n_96),
.B(n_97),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1956),
.A2(n_566),
.B(n_565),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1914),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1888),
.B(n_100),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_1864),
.A2(n_568),
.B(n_567),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_1960),
.Y(n_2107)
);

INVxp67_ASAP7_75t_L g2108 ( 
.A(n_1872),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1965),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1871),
.B(n_1907),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1908),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1897),
.B(n_101),
.Y(n_2112)
);

AOI221x1_ASAP7_75t_L g2113 ( 
.A1(n_1949),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.C(n_104),
.Y(n_2113)
);

OAI21x1_ASAP7_75t_L g2114 ( 
.A1(n_1985),
.A2(n_571),
.B(n_569),
.Y(n_2114)
);

INVx5_ASAP7_75t_L g2115 ( 
.A(n_1929),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_2004),
.A2(n_574),
.B(n_572),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1990),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1910),
.Y(n_2118)
);

OAI21x1_ASAP7_75t_SL g2119 ( 
.A1(n_1902),
.A2(n_1943),
.B(n_2030),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_2011),
.A2(n_576),
.B(n_575),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_1998),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_SL g2122 ( 
.A1(n_1931),
.A2(n_103),
.B(n_104),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1951),
.B(n_577),
.Y(n_2123)
);

A2O1A1Ixp33_ASAP7_75t_L g2124 ( 
.A1(n_1882),
.A2(n_108),
.B(n_105),
.C(n_106),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_2016),
.A2(n_579),
.B(n_578),
.Y(n_2125)
);

AO21x1_ASAP7_75t_L g2126 ( 
.A1(n_1950),
.A2(n_2019),
.B(n_2028),
.Y(n_2126)
);

OAI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1881),
.A2(n_105),
.B(n_106),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1859),
.A2(n_582),
.B(n_580),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2012),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_SL g2130 ( 
.A1(n_1955),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2014),
.B(n_584),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1903),
.B(n_109),
.Y(n_2132)
);

INVx5_ASAP7_75t_L g2133 ( 
.A(n_1929),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_1868),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1906),
.B(n_111),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_SL g2136 ( 
.A1(n_1959),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_2017),
.A2(n_2021),
.B(n_2027),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_1891),
.A2(n_112),
.B(n_113),
.Y(n_2138)
);

O2A1O1Ixp5_ASAP7_75t_SL g2139 ( 
.A1(n_1975),
.A2(n_119),
.B(n_116),
.C(n_118),
.Y(n_2139)
);

AOI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2006),
.A2(n_1939),
.B1(n_1997),
.B2(n_1920),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2026),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1893),
.B(n_116),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1900),
.B(n_585),
.Y(n_2143)
);

CKINVDCx20_ASAP7_75t_R g2144 ( 
.A(n_1942),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_1966),
.A2(n_589),
.B(n_588),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1945),
.B(n_118),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1941),
.B(n_1969),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_2054),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2107),
.B(n_1962),
.Y(n_2149)
);

INVx3_ASAP7_75t_SL g2150 ( 
.A(n_2118),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2141),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2053),
.B(n_1892),
.Y(n_2152)
);

BUFx4_ASAP7_75t_SL g2153 ( 
.A(n_2144),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2121),
.Y(n_2154)
);

AOI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_2037),
.A2(n_2022),
.B(n_2013),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_SL g2156 ( 
.A(n_2131),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2035),
.A2(n_1978),
.B1(n_1957),
.B2(n_1937),
.Y(n_2157)
);

OR2x6_ASAP7_75t_L g2158 ( 
.A(n_2039),
.B(n_1957),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_2107),
.B(n_1924),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_2094),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2061),
.A2(n_2010),
.B(n_1894),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2078),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2091),
.B(n_1877),
.Y(n_2163)
);

AO32x1_ASAP7_75t_L g2164 ( 
.A1(n_2104),
.A2(n_2069),
.A3(n_1952),
.B1(n_1984),
.B2(n_2101),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_2115),
.B(n_1867),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_2058),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2109),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_2050),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_2121),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2117),
.B(n_2007),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2065),
.B(n_1916),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_2061),
.A2(n_2024),
.B(n_2015),
.Y(n_2172)
);

INVx5_ASAP7_75t_L g2173 ( 
.A(n_2115),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2137),
.A2(n_1995),
.B(n_1989),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2129),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2032),
.Y(n_2176)
);

A2O1A1Ixp33_ASAP7_75t_SL g2177 ( 
.A1(n_2127),
.A2(n_1874),
.B(n_1919),
.C(n_1973),
.Y(n_2177)
);

BUFx2_ASAP7_75t_SL g2178 ( 
.A(n_2115),
.Y(n_2178)
);

INVx5_ASAP7_75t_L g2179 ( 
.A(n_2133),
.Y(n_2179)
);

INVx8_ASAP7_75t_L g2180 ( 
.A(n_2133),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_2066),
.A2(n_1979),
.B(n_1915),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2134),
.B(n_2025),
.Y(n_2182)
);

NAND2x1p5_ASAP7_75t_L g2183 ( 
.A(n_2133),
.B(n_2043),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2147),
.B(n_1934),
.Y(n_2184)
);

A2O1A1Ixp33_ASAP7_75t_L g2185 ( 
.A1(n_2070),
.A2(n_1901),
.B(n_1879),
.C(n_1909),
.Y(n_2185)
);

NAND2xp33_ASAP7_75t_L g2186 ( 
.A(n_2071),
.B(n_1974),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2031),
.B(n_1884),
.Y(n_2187)
);

O2A1O1Ixp33_ASAP7_75t_L g2188 ( 
.A1(n_2088),
.A2(n_1987),
.B(n_1991),
.C(n_1988),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2038),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2044),
.Y(n_2190)
);

O2A1O1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_2124),
.A2(n_1992),
.B(n_1994),
.C(n_1993),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2085),
.B(n_2000),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_2123),
.B(n_2023),
.Y(n_2193)
);

INVx4_ASAP7_75t_L g2194 ( 
.A(n_2047),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2057),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2068),
.A2(n_1925),
.B(n_1880),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2108),
.B(n_1889),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2099),
.B(n_1889),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_2047),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2040),
.A2(n_2008),
.B(n_2009),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2043),
.B(n_1998),
.Y(n_2201)
);

O2A1O1Ixp5_ASAP7_75t_L g2202 ( 
.A1(n_2099),
.A2(n_1984),
.B(n_1927),
.C(n_1925),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2067),
.B(n_1984),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2042),
.Y(n_2204)
);

OAI22xp5_ASAP7_75t_SL g2205 ( 
.A1(n_2130),
.A2(n_1977),
.B1(n_1981),
.B2(n_1938),
.Y(n_2205)
);

AOI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2097),
.A2(n_2110),
.B(n_2096),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2084),
.B(n_1938),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2084),
.B(n_1977),
.Y(n_2208)
);

BUFx10_ASAP7_75t_L g2209 ( 
.A(n_2131),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2057),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2059),
.B(n_1977),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_2126),
.A2(n_1986),
.B1(n_1981),
.B2(n_122),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_2042),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2049),
.B(n_1981),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2075),
.Y(n_2215)
);

OA21x2_ASAP7_75t_L g2216 ( 
.A1(n_2074),
.A2(n_1986),
.B(n_119),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2071),
.B(n_1986),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_2055),
.B(n_120),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2049),
.B(n_120),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2077),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2052),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2111),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2047),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_2096),
.A2(n_2040),
.B(n_2102),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2136),
.B(n_123),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2166),
.B(n_2041),
.Y(n_2226)
);

HB1xp67_ASAP7_75t_L g2227 ( 
.A(n_2148),
.Y(n_2227)
);

INVx6_ASAP7_75t_L g2228 ( 
.A(n_2173),
.Y(n_2228)
);

INVx8_ASAP7_75t_L g2229 ( 
.A(n_2180),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2163),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2167),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2162),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2198),
.A2(n_2140),
.B1(n_2130),
.B2(n_2080),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2175),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_2153),
.Y(n_2235)
);

CKINVDCx20_ASAP7_75t_R g2236 ( 
.A(n_2150),
.Y(n_2236)
);

AOI21xp33_ASAP7_75t_L g2237 ( 
.A1(n_2177),
.A2(n_2138),
.B(n_2102),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2180),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_SL g2239 ( 
.A1(n_2198),
.A2(n_2119),
.B1(n_2082),
.B2(n_2095),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2186),
.A2(n_2140),
.B1(n_2122),
.B2(n_2080),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2158),
.A2(n_2136),
.B1(n_2056),
.B2(n_2106),
.Y(n_2241)
);

BUFx10_ASAP7_75t_L g2242 ( 
.A(n_2168),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2151),
.Y(n_2243)
);

BUFx2_ASAP7_75t_L g2244 ( 
.A(n_2149),
.Y(n_2244)
);

NAND2x1p5_ASAP7_75t_L g2245 ( 
.A(n_2173),
.B(n_2051),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2189),
.B(n_2086),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2149),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_2160),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2176),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_SL g2250 ( 
.A1(n_2205),
.A2(n_2083),
.B1(n_2073),
.B2(n_2087),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_SL g2251 ( 
.A1(n_2224),
.A2(n_2100),
.B1(n_2093),
.B2(n_2051),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_L g2252 ( 
.A1(n_2172),
.A2(n_2143),
.B1(n_2105),
.B2(n_2142),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2163),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2181),
.A2(n_2146),
.B1(n_2135),
.B2(n_2132),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2159),
.Y(n_2255)
);

INVx6_ASAP7_75t_L g2256 ( 
.A(n_2173),
.Y(n_2256)
);

AOI21xp33_ASAP7_75t_L g2257 ( 
.A1(n_2188),
.A2(n_2112),
.B(n_2063),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2204),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2195),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_SL g2260 ( 
.A1(n_2225),
.A2(n_2156),
.B1(n_2206),
.B2(n_2218),
.Y(n_2260)
);

BUFx8_ASAP7_75t_L g2261 ( 
.A(n_2219),
.Y(n_2261)
);

BUFx2_ASAP7_75t_SL g2262 ( 
.A(n_2156),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2190),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2213),
.Y(n_2264)
);

CKINVDCx6p67_ASAP7_75t_R g2265 ( 
.A(n_2180),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2187),
.B(n_2086),
.Y(n_2266)
);

INVx4_ASAP7_75t_L g2267 ( 
.A(n_2173),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_2171),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2158),
.A2(n_2081),
.B1(n_2090),
.B2(n_2089),
.Y(n_2269)
);

BUFx10_ASAP7_75t_L g2270 ( 
.A(n_2197),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2158),
.A2(n_2128),
.B1(n_2034),
.B2(n_2045),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2157),
.A2(n_2034),
.B1(n_2079),
.B2(n_2103),
.Y(n_2272)
);

CKINVDCx6p67_ASAP7_75t_R g2273 ( 
.A(n_2179),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_L g2274 ( 
.A1(n_2200),
.A2(n_2114),
.B1(n_2120),
.B2(n_2116),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2230),
.B(n_2152),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2258),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2253),
.B(n_2203),
.Y(n_2277)
);

O2A1O1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_2237),
.A2(n_2257),
.B(n_2225),
.C(n_2200),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2231),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2255),
.B(n_2182),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2233),
.A2(n_2212),
.B1(n_2208),
.B2(n_2207),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2240),
.A2(n_2208),
.B1(n_2207),
.B2(n_2217),
.Y(n_2282)
);

BUFx10_ASAP7_75t_L g2283 ( 
.A(n_2228),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2244),
.B(n_2216),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2227),
.B(n_2221),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2263),
.B(n_2187),
.Y(n_2286)
);

O2A1O1Ixp5_ASAP7_75t_L g2287 ( 
.A1(n_2237),
.A2(n_2202),
.B(n_2155),
.C(n_2165),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2257),
.A2(n_2174),
.B(n_2161),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2264),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2267),
.B(n_2179),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2239),
.A2(n_2217),
.B1(n_2185),
.B2(n_2192),
.Y(n_2291)
);

OA21x2_ASAP7_75t_L g2292 ( 
.A1(n_2266),
.A2(n_2170),
.B(n_2113),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2266),
.B(n_2170),
.Y(n_2293)
);

OA21x2_ASAP7_75t_L g2294 ( 
.A1(n_2246),
.A2(n_2201),
.B(n_2033),
.Y(n_2294)
);

OA21x2_ASAP7_75t_L g2295 ( 
.A1(n_2274),
.A2(n_2201),
.B(n_2064),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2247),
.B(n_2216),
.Y(n_2296)
);

O2A1O1Ixp5_ASAP7_75t_L g2297 ( 
.A1(n_2226),
.A2(n_2184),
.B(n_2196),
.C(n_2215),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2234),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2247),
.B(n_2211),
.Y(n_2299)
);

INVxp67_ASAP7_75t_L g2300 ( 
.A(n_2268),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2228),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2279),
.Y(n_2302)
);

CKINVDCx20_ASAP7_75t_R g2303 ( 
.A(n_2300),
.Y(n_2303)
);

NAND2xp33_ASAP7_75t_R g2304 ( 
.A(n_2301),
.B(n_2235),
.Y(n_2304)
);

AO31x2_ASAP7_75t_L g2305 ( 
.A1(n_2288),
.A2(n_2267),
.A3(n_2249),
.B(n_2232),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_2283),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2291),
.A2(n_2260),
.B1(n_2252),
.B2(n_2251),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2279),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2291),
.A2(n_2260),
.B1(n_2241),
.B2(n_2250),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2275),
.B(n_2262),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2286),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_R g2312 ( 
.A(n_2292),
.B(n_2248),
.Y(n_2312)
);

OA21x2_ASAP7_75t_L g2313 ( 
.A1(n_2307),
.A2(n_2297),
.B(n_2287),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2308),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_2307),
.A2(n_2293),
.B(n_2296),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2311),
.B(n_2275),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2302),
.B(n_2293),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2305),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2305),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2305),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_2313),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2313),
.A2(n_2309),
.B(n_2278),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2315),
.A2(n_2281),
.B1(n_2282),
.B2(n_2254),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2320),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2314),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2316),
.B(n_2299),
.Y(n_2326)
);

OR2x2_ASAP7_75t_L g2327 ( 
.A(n_2315),
.B(n_2299),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2314),
.B(n_2305),
.Y(n_2328)
);

INVx1_ASAP7_75t_SL g2329 ( 
.A(n_2313),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2313),
.B(n_2280),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2325),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2328),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2330),
.B(n_2310),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2328),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2321),
.Y(n_2335)
);

OAI22xp33_ASAP7_75t_L g2336 ( 
.A1(n_2322),
.A2(n_2312),
.B1(n_2315),
.B2(n_2281),
.Y(n_2336)
);

INVxp67_ASAP7_75t_L g2337 ( 
.A(n_2329),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2328),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2324),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2326),
.B(n_2306),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2324),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2327),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2336),
.B(n_2236),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_2335),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2342),
.B(n_2315),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2335),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2333),
.B(n_2323),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2339),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2340),
.B(n_2323),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2341),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2331),
.Y(n_2351)
);

NOR2xp67_ASAP7_75t_L g2352 ( 
.A(n_2345),
.B(n_2337),
.Y(n_2352)
);

AND3x2_ASAP7_75t_L g2353 ( 
.A(n_2344),
.B(n_2337),
.C(n_2334),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2346),
.B(n_2332),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2349),
.B(n_2338),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_2353),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2355),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2352),
.Y(n_2358)
);

AND2x4_ASAP7_75t_SL g2359 ( 
.A(n_2354),
.B(n_2242),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2357),
.B(n_2358),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2356),
.Y(n_2361)
);

INVxp67_ASAP7_75t_SL g2362 ( 
.A(n_2359),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2359),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2357),
.B(n_2347),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_L g2365 ( 
.A(n_2356),
.B(n_2336),
.C(n_2343),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2365),
.A2(n_2347),
.B1(n_2343),
.B2(n_2349),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2364),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2360),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2361),
.B(n_2348),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2362),
.B(n_2351),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2363),
.A2(n_2350),
.B1(n_2334),
.B2(n_2320),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2365),
.B(n_2242),
.Y(n_2372)
);

OR2x2_ASAP7_75t_L g2373 ( 
.A(n_2364),
.B(n_2317),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2364),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2364),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2367),
.B(n_2303),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2374),
.B(n_2317),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2369),
.Y(n_2378)
);

AO22x1_ASAP7_75t_L g2379 ( 
.A1(n_2368),
.A2(n_2261),
.B1(n_2312),
.B2(n_2319),
.Y(n_2379)
);

OA21x2_ASAP7_75t_L g2380 ( 
.A1(n_2366),
.A2(n_2319),
.B(n_2320),
.Y(n_2380)
);

OAI211xp5_ASAP7_75t_L g2381 ( 
.A1(n_2372),
.A2(n_2318),
.B(n_2179),
.C(n_2301),
.Y(n_2381)
);

BUFx2_ASAP7_75t_L g2382 ( 
.A(n_2375),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2370),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2371),
.B(n_2373),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2370),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2366),
.B(n_2318),
.Y(n_2386)
);

OAI211xp5_ASAP7_75t_L g2387 ( 
.A1(n_2366),
.A2(n_2179),
.B(n_2301),
.C(n_2229),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2370),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2376),
.A2(n_2285),
.B(n_2282),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2382),
.B(n_2298),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2377),
.Y(n_2391)
);

AND2x2_ASAP7_75t_SL g2392 ( 
.A(n_2384),
.B(n_2290),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2378),
.B(n_2298),
.Y(n_2393)
);

AOI221xp5_ASAP7_75t_L g2394 ( 
.A1(n_2387),
.A2(n_2378),
.B1(n_2386),
.B2(n_2381),
.C(n_2383),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2385),
.B(n_2280),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2388),
.Y(n_2396)
);

OAI221xp5_ASAP7_75t_SL g2397 ( 
.A1(n_2379),
.A2(n_2265),
.B1(n_2301),
.B2(n_2220),
.C(n_2271),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2380),
.A2(n_2304),
.B1(n_2270),
.B2(n_2178),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2380),
.B(n_2276),
.Y(n_2399)
);

INVx1_ASAP7_75t_SL g2400 ( 
.A(n_2376),
.Y(n_2400)
);

INVx1_ASAP7_75t_SL g2401 ( 
.A(n_2376),
.Y(n_2401)
);

INVx1_ASAP7_75t_SL g2402 ( 
.A(n_2376),
.Y(n_2402)
);

AOI32xp33_ASAP7_75t_L g2403 ( 
.A1(n_2376),
.A2(n_2284),
.A3(n_2296),
.B1(n_2290),
.B2(n_2238),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2392),
.B(n_2270),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2398),
.B(n_2283),
.Y(n_2405)
);

INVxp67_ASAP7_75t_L g2406 ( 
.A(n_2391),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2395),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2400),
.B(n_2401),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2402),
.B(n_2261),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2389),
.B(n_2277),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2396),
.B(n_2284),
.Y(n_2411)
);

INVx1_ASAP7_75t_SL g2412 ( 
.A(n_2393),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2394),
.B(n_2276),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_SL g2414 ( 
.A(n_2397),
.B(n_2229),
.Y(n_2414)
);

OAI221xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2403),
.A2(n_2273),
.B1(n_2191),
.B2(n_2238),
.C(n_2272),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_2390),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2399),
.B(n_2277),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_L g2418 ( 
.A(n_2406),
.B(n_124),
.C(n_125),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2409),
.A2(n_2229),
.B(n_2290),
.Y(n_2419)
);

NOR3xp33_ASAP7_75t_L g2420 ( 
.A(n_2408),
.B(n_2290),
.C(n_124),
.Y(n_2420)
);

HB1xp67_ASAP7_75t_L g2421 ( 
.A(n_2404),
.Y(n_2421)
);

NOR3xp33_ASAP7_75t_L g2422 ( 
.A(n_2407),
.B(n_125),
.C(n_127),
.Y(n_2422)
);

OAI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2405),
.A2(n_2139),
.B(n_2125),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2411),
.Y(n_2424)
);

OAI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2414),
.A2(n_2256),
.B1(n_2228),
.B2(n_2289),
.Y(n_2425)
);

HB1xp67_ASAP7_75t_L g2426 ( 
.A(n_2412),
.Y(n_2426)
);

NAND4xp25_ASAP7_75t_L g2427 ( 
.A(n_2414),
.B(n_2193),
.C(n_129),
.D(n_127),
.Y(n_2427)
);

NOR5xp2_ASAP7_75t_L g2428 ( 
.A(n_2415),
.B(n_130),
.C(n_128),
.D(n_129),
.E(n_131),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2413),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2416),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2410),
.B(n_2292),
.Y(n_2431)
);

AND3x4_ASAP7_75t_L g2432 ( 
.A(n_2417),
.B(n_2283),
.C(n_2279),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2408),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2408),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2409),
.B(n_128),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2409),
.B(n_131),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2408),
.Y(n_2437)
);

OA22x2_ASAP7_75t_L g2438 ( 
.A1(n_2409),
.A2(n_2289),
.B1(n_2199),
.B2(n_2194),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2408),
.B(n_2292),
.Y(n_2439)
);

OAI211xp5_ASAP7_75t_L g2440 ( 
.A1(n_2427),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2440)
);

NAND4xp25_ASAP7_75t_L g2441 ( 
.A(n_2434),
.B(n_134),
.C(n_132),
.D(n_133),
.Y(n_2441)
);

AOI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2425),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_2433),
.B(n_2283),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2420),
.B(n_135),
.Y(n_2444)
);

O2A1O1Ixp33_ASAP7_75t_L g2445 ( 
.A1(n_2426),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_2445)
);

AOI211x1_ASAP7_75t_L g2446 ( 
.A1(n_2419),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2437),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2421),
.B(n_2292),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2424),
.B(n_139),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2435),
.B(n_2436),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2430),
.B(n_2214),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2418),
.Y(n_2452)
);

NAND3xp33_ASAP7_75t_L g2453 ( 
.A(n_2422),
.B(n_140),
.C(n_141),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2439),
.B(n_142),
.Y(n_2454)
);

AOI322xp5_ASAP7_75t_L g2455 ( 
.A1(n_2429),
.A2(n_2269),
.A3(n_2223),
.B1(n_2164),
.B2(n_2243),
.C1(n_2259),
.C2(n_2092),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2432),
.Y(n_2456)
);

INVxp67_ASAP7_75t_L g2457 ( 
.A(n_2431),
.Y(n_2457)
);

OAI321xp33_ASAP7_75t_L g2458 ( 
.A1(n_2428),
.A2(n_2048),
.A3(n_2183),
.B1(n_2245),
.B2(n_2098),
.C(n_2092),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2438),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_SL g2460 ( 
.A(n_2423),
.B(n_2183),
.C(n_143),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2433),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2433),
.Y(n_2462)
);

AND2x2_ASAP7_75t_SL g2463 ( 
.A(n_2428),
.B(n_2194),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2433),
.B(n_143),
.Y(n_2464)
);

NAND3xp33_ASAP7_75t_SL g2465 ( 
.A(n_2420),
.B(n_144),
.C(n_145),
.Y(n_2465)
);

AOI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2420),
.A2(n_2256),
.B1(n_2199),
.B2(n_2092),
.Y(n_2466)
);

OAI211xp5_ASAP7_75t_L g2467 ( 
.A1(n_2427),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2467)
);

NOR3xp33_ASAP7_75t_L g2468 ( 
.A(n_2433),
.B(n_146),
.C(n_147),
.Y(n_2468)
);

NAND3xp33_ASAP7_75t_L g2469 ( 
.A(n_2420),
.B(n_148),
.C(n_149),
.Y(n_2469)
);

AND4x1_ASAP7_75t_L g2470 ( 
.A(n_2435),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2433),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2434),
.A2(n_2256),
.B1(n_2098),
.B2(n_2072),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2433),
.B(n_2294),
.Y(n_2473)
);

NAND4xp25_ASAP7_75t_L g2474 ( 
.A(n_2427),
.B(n_152),
.C(n_150),
.D(n_151),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2434),
.A2(n_2072),
.B1(n_2098),
.B2(n_2223),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2433),
.B(n_151),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2463),
.B(n_2294),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_L g2478 ( 
.A(n_2446),
.B(n_2461),
.C(n_2462),
.D(n_2471),
.Y(n_2478)
);

NOR2x1_ASAP7_75t_L g2479 ( 
.A(n_2441),
.B(n_152),
.Y(n_2479)
);

NOR3x1_ASAP7_75t_L g2480 ( 
.A(n_2469),
.B(n_154),
.C(n_155),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2442),
.B(n_154),
.C(n_155),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2464),
.B(n_156),
.Y(n_2482)
);

AOI211xp5_ASAP7_75t_L g2483 ( 
.A1(n_2440),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2483)
);

NAND4xp25_ASAP7_75t_L g2484 ( 
.A(n_2447),
.B(n_160),
.C(n_158),
.D(n_159),
.Y(n_2484)
);

INVxp67_ASAP7_75t_SL g2485 ( 
.A(n_2445),
.Y(n_2485)
);

NAND4xp25_ASAP7_75t_L g2486 ( 
.A(n_2450),
.B(n_162),
.C(n_160),
.D(n_161),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2470),
.B(n_161),
.Y(n_2487)
);

NOR3xp33_ASAP7_75t_L g2488 ( 
.A(n_2444),
.B(n_162),
.C(n_163),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2476),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2465),
.B(n_164),
.C(n_165),
.Y(n_2490)
);

AOI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2472),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2449),
.B(n_166),
.Y(n_2492)
);

AND3x2_ASAP7_75t_L g2493 ( 
.A(n_2468),
.B(n_168),
.C(n_169),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2458),
.B(n_2072),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2466),
.B(n_169),
.Y(n_2495)
);

AOI221x1_ASAP7_75t_L g2496 ( 
.A1(n_2454),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.C(n_173),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2453),
.B(n_171),
.C(n_172),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2448),
.B(n_174),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2451),
.B(n_174),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_L g2500 ( 
.A(n_2467),
.B(n_175),
.C(n_176),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2474),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2473),
.Y(n_2502)
);

OAI21xp33_ASAP7_75t_L g2503 ( 
.A1(n_2466),
.A2(n_2459),
.B(n_2452),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2443),
.B(n_175),
.Y(n_2504)
);

NOR4xp25_ASAP7_75t_L g2505 ( 
.A(n_2457),
.B(n_178),
.C(n_176),
.D(n_177),
.Y(n_2505)
);

O2A1O1Ixp5_ASAP7_75t_SL g2506 ( 
.A1(n_2456),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2475),
.B(n_179),
.Y(n_2507)
);

AOI211xp5_ASAP7_75t_L g2508 ( 
.A1(n_2460),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2508)
);

NAND4xp75_ASAP7_75t_L g2509 ( 
.A(n_2455),
.B(n_182),
.C(n_180),
.D(n_181),
.Y(n_2509)
);

OA211x2_ASAP7_75t_L g2510 ( 
.A1(n_2465),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2510)
);

OAI222xp33_ASAP7_75t_L g2511 ( 
.A1(n_2461),
.A2(n_2245),
.B1(n_185),
.B2(n_186),
.C1(n_187),
.C2(n_188),
.Y(n_2511)
);

NAND4xp25_ASAP7_75t_L g2512 ( 
.A(n_2446),
.B(n_187),
.C(n_183),
.D(n_186),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2442),
.B(n_188),
.C(n_189),
.Y(n_2513)
);

AOI222xp33_ASAP7_75t_L g2514 ( 
.A1(n_2443),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.C1(n_193),
.C2(n_194),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_SL g2515 ( 
.A(n_2483),
.B(n_190),
.C(n_191),
.Y(n_2515)
);

AOI211xp5_ASAP7_75t_L g2516 ( 
.A1(n_2505),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2516)
);

NAND3xp33_ASAP7_75t_L g2517 ( 
.A(n_2514),
.B(n_196),
.C(n_197),
.Y(n_2517)
);

NAND4xp25_ASAP7_75t_L g2518 ( 
.A(n_2508),
.B(n_199),
.C(n_197),
.D(n_198),
.Y(n_2518)
);

AOI21xp33_ASAP7_75t_L g2519 ( 
.A1(n_2503),
.A2(n_199),
.B(n_200),
.Y(n_2519)
);

NOR3x1_ASAP7_75t_L g2520 ( 
.A(n_2500),
.B(n_200),
.C(n_201),
.Y(n_2520)
);

NAND3xp33_ASAP7_75t_SL g2521 ( 
.A(n_2490),
.B(n_2488),
.C(n_2506),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_SL g2522 ( 
.A(n_2478),
.B(n_201),
.Y(n_2522)
);

NAND3xp33_ASAP7_75t_SL g2523 ( 
.A(n_2487),
.B(n_202),
.C(n_203),
.Y(n_2523)
);

AOI21xp33_ASAP7_75t_SL g2524 ( 
.A1(n_2498),
.A2(n_202),
.B(n_203),
.Y(n_2524)
);

NOR3xp33_ASAP7_75t_L g2525 ( 
.A(n_2485),
.B(n_204),
.C(n_205),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2493),
.B(n_204),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2479),
.B(n_2294),
.Y(n_2527)
);

OAI221xp5_ASAP7_75t_SL g2528 ( 
.A1(n_2501),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.C(n_208),
.Y(n_2528)
);

NOR3xp33_ASAP7_75t_L g2529 ( 
.A(n_2482),
.B(n_206),
.C(n_208),
.Y(n_2529)
);

NOR3xp33_ASAP7_75t_L g2530 ( 
.A(n_2492),
.B(n_2489),
.C(n_2497),
.Y(n_2530)
);

NAND4xp75_ASAP7_75t_L g2531 ( 
.A(n_2510),
.B(n_211),
.C(n_209),
.D(n_210),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2512),
.B(n_210),
.Y(n_2532)
);

NAND4xp25_ASAP7_75t_SL g2533 ( 
.A(n_2481),
.B(n_214),
.C(n_211),
.D(n_213),
.Y(n_2533)
);

NAND3x1_ASAP7_75t_L g2534 ( 
.A(n_2504),
.B(n_2499),
.C(n_2507),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2480),
.B(n_2294),
.Y(n_2535)
);

OAI21xp33_ASAP7_75t_L g2536 ( 
.A1(n_2494),
.A2(n_2145),
.B(n_2062),
.Y(n_2536)
);

AOI322xp5_ASAP7_75t_L g2537 ( 
.A1(n_2495),
.A2(n_213),
.A3(n_214),
.B1(n_215),
.B2(n_216),
.C1(n_217),
.C2(n_219),
.Y(n_2537)
);

OAI211xp5_ASAP7_75t_SL g2538 ( 
.A1(n_2502),
.A2(n_219),
.B(n_216),
.C(n_217),
.Y(n_2538)
);

NOR2xp67_ASAP7_75t_L g2539 ( 
.A(n_2484),
.B(n_220),
.Y(n_2539)
);

NAND3xp33_ASAP7_75t_L g2540 ( 
.A(n_2491),
.B(n_220),
.C(n_221),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2496),
.B(n_221),
.Y(n_2541)
);

AOI211xp5_ASAP7_75t_L g2542 ( 
.A1(n_2513),
.A2(n_2511),
.B(n_2486),
.C(n_2477),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2509),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.C(n_225),
.Y(n_2543)
);

NOR3xp33_ASAP7_75t_L g2544 ( 
.A(n_2478),
.B(n_222),
.C(n_223),
.Y(n_2544)
);

NOR3xp33_ASAP7_75t_L g2545 ( 
.A(n_2478),
.B(n_224),
.C(n_225),
.Y(n_2545)
);

NOR3xp33_ASAP7_75t_L g2546 ( 
.A(n_2478),
.B(n_227),
.C(n_228),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2498),
.Y(n_2547)
);

NOR3xp33_ASAP7_75t_L g2548 ( 
.A(n_2478),
.B(n_227),
.C(n_228),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2498),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2485),
.A2(n_229),
.B(n_230),
.Y(n_2550)
);

NAND2xp33_ASAP7_75t_R g2551 ( 
.A(n_2493),
.B(n_229),
.Y(n_2551)
);

OAI211xp5_ASAP7_75t_L g2552 ( 
.A1(n_2503),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2500),
.A2(n_2295),
.B1(n_2154),
.B2(n_2169),
.Y(n_2553)
);

AND4x1_ASAP7_75t_L g2554 ( 
.A(n_2505),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2554)
);

NAND4xp25_ASAP7_75t_SL g2555 ( 
.A(n_2508),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2555)
);

A2O1A1Ixp33_ASAP7_75t_L g2556 ( 
.A1(n_2487),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_2556)
);

OAI211xp5_ASAP7_75t_L g2557 ( 
.A1(n_2503),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_2557)
);

OAI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2503),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.C(n_243),
.Y(n_2558)
);

NAND3xp33_ASAP7_75t_SL g2559 ( 
.A(n_2483),
.B(n_240),
.C(n_241),
.Y(n_2559)
);

AOI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2485),
.A2(n_242),
.B(n_243),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2493),
.B(n_244),
.Y(n_2561)
);

AOI211xp5_ASAP7_75t_L g2562 ( 
.A1(n_2505),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_2562)
);

OR2x2_ASAP7_75t_L g2563 ( 
.A(n_2505),
.B(n_245),
.Y(n_2563)
);

NOR2x1_ASAP7_75t_L g2564 ( 
.A(n_2484),
.B(n_246),
.Y(n_2564)
);

OAI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2503),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.C(n_251),
.Y(n_2565)
);

O2A1O1Ixp33_ASAP7_75t_L g2566 ( 
.A1(n_2498),
.A2(n_251),
.B(n_248),
.C(n_249),
.Y(n_2566)
);

NAND4xp25_ASAP7_75t_L g2567 ( 
.A(n_2508),
.B(n_254),
.C(n_252),
.D(n_253),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2512),
.B(n_253),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2505),
.B(n_255),
.Y(n_2569)
);

AOI211x1_ASAP7_75t_L g2570 ( 
.A1(n_2494),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2493),
.B(n_256),
.Y(n_2571)
);

OAI311xp33_ASAP7_75t_L g2572 ( 
.A1(n_2503),
.A2(n_258),
.A3(n_260),
.B1(n_261),
.C1(n_262),
.Y(n_2572)
);

NOR5xp2_ASAP7_75t_L g2573 ( 
.A(n_2503),
.B(n_258),
.C(n_261),
.D(n_262),
.E(n_263),
.Y(n_2573)
);

NOR3x1_ASAP7_75t_L g2574 ( 
.A(n_2500),
.B(n_263),
.C(n_264),
.Y(n_2574)
);

NAND4xp75_ASAP7_75t_L g2575 ( 
.A(n_2510),
.B(n_267),
.C(n_265),
.D(n_266),
.Y(n_2575)
);

AOI211xp5_ASAP7_75t_SL g2576 ( 
.A1(n_2503),
.A2(n_268),
.B(n_265),
.C(n_267),
.Y(n_2576)
);

NAND4xp75_ASAP7_75t_L g2577 ( 
.A(n_2520),
.B(n_271),
.C(n_268),
.D(n_269),
.Y(n_2577)
);

INVx2_ASAP7_75t_SL g2578 ( 
.A(n_2554),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2526),
.Y(n_2579)
);

OAI22xp5_ASAP7_75t_SL g2580 ( 
.A1(n_2570),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_2580)
);

HB1xp67_ASAP7_75t_L g2581 ( 
.A(n_2531),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2561),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_R g2583 ( 
.A(n_2551),
.B(n_272),
.Y(n_2583)
);

AOI222xp33_ASAP7_75t_L g2584 ( 
.A1(n_2515),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.C1(n_277),
.C2(n_278),
.Y(n_2584)
);

AOI211xp5_ASAP7_75t_L g2585 ( 
.A1(n_2519),
.A2(n_278),
.B(n_275),
.C(n_277),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2576),
.B(n_279),
.Y(n_2586)
);

NOR2x1_ASAP7_75t_L g2587 ( 
.A(n_2575),
.B(n_281),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2571),
.Y(n_2588)
);

OAI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2522),
.A2(n_2295),
.B1(n_2169),
.B2(n_2154),
.Y(n_2589)
);

NAND3xp33_ASAP7_75t_L g2590 ( 
.A(n_2544),
.B(n_281),
.C(n_282),
.Y(n_2590)
);

INVxp33_ASAP7_75t_L g2591 ( 
.A(n_2532),
.Y(n_2591)
);

AOI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2545),
.A2(n_2295),
.B1(n_2209),
.B2(n_2222),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2547),
.Y(n_2593)
);

CKINVDCx16_ASAP7_75t_R g2594 ( 
.A(n_2522),
.Y(n_2594)
);

CKINVDCx6p67_ASAP7_75t_R g2595 ( 
.A(n_2569),
.Y(n_2595)
);

AOI211xp5_ASAP7_75t_L g2596 ( 
.A1(n_2572),
.A2(n_286),
.B(n_283),
.C(n_284),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2564),
.B(n_2295),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2541),
.Y(n_2598)
);

XNOR2xp5_ASAP7_75t_L g2599 ( 
.A(n_2534),
.B(n_283),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2516),
.B(n_2562),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2539),
.B(n_286),
.Y(n_2601)
);

NOR3xp33_ASAP7_75t_L g2602 ( 
.A(n_2523),
.B(n_287),
.C(n_288),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2563),
.Y(n_2603)
);

O2A1O1Ixp33_ASAP7_75t_L g2604 ( 
.A1(n_2556),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2604)
);

AOI22xp5_ASAP7_75t_L g2605 ( 
.A1(n_2546),
.A2(n_2209),
.B1(n_2210),
.B2(n_2076),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2524),
.B(n_289),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2568),
.Y(n_2607)
);

OAI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2558),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2521),
.A2(n_290),
.B(n_291),
.Y(n_2609)
);

NAND3xp33_ASAP7_75t_L g2610 ( 
.A(n_2548),
.B(n_292),
.C(n_294),
.Y(n_2610)
);

NOR3xp33_ASAP7_75t_L g2611 ( 
.A(n_2565),
.B(n_295),
.C(n_296),
.Y(n_2611)
);

BUFx2_ASAP7_75t_L g2612 ( 
.A(n_2518),
.Y(n_2612)
);

OAI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2517),
.A2(n_2060),
.B(n_2036),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2552),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2540),
.A2(n_2046),
.B1(n_298),
.B2(n_296),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2537),
.B(n_297),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2557),
.Y(n_2617)
);

OAI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2543),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.C(n_300),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2525),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2550),
.Y(n_2620)
);

NOR2x1_ASAP7_75t_L g2621 ( 
.A(n_2533),
.B(n_301),
.Y(n_2621)
);

AOI21xp33_ASAP7_75t_SL g2622 ( 
.A1(n_2566),
.A2(n_301),
.B(n_302),
.Y(n_2622)
);

INVxp67_ASAP7_75t_L g2623 ( 
.A(n_2555),
.Y(n_2623)
);

NAND2xp33_ASAP7_75t_R g2624 ( 
.A(n_2560),
.B(n_303),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2559),
.A2(n_306),
.B1(n_303),
.B2(n_305),
.Y(n_2625)
);

AOI211xp5_ASAP7_75t_L g2626 ( 
.A1(n_2538),
.A2(n_305),
.B(n_307),
.C(n_308),
.Y(n_2626)
);

OAI211xp5_ASAP7_75t_SL g2627 ( 
.A1(n_2542),
.A2(n_307),
.B(n_308),
.C(n_310),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2574),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2529),
.B(n_310),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2567),
.Y(n_2630)
);

OAI211xp5_ASAP7_75t_L g2631 ( 
.A1(n_2530),
.A2(n_311),
.B(n_312),
.C(n_313),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_2549),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2535),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_2633)
);

OAI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2553),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2527),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2573),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2528),
.B(n_315),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2536),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_2638)
);

NOR2x1p5_ASAP7_75t_L g2639 ( 
.A(n_2531),
.B(n_317),
.Y(n_2639)
);

OAI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2539),
.A2(n_318),
.B(n_319),
.Y(n_2640)
);

OAI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2539),
.A2(n_320),
.B(n_321),
.Y(n_2641)
);

XOR2x1_ASAP7_75t_L g2642 ( 
.A(n_2639),
.B(n_320),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2581),
.B(n_321),
.Y(n_2643)
);

NAND2x1p5_ASAP7_75t_L g2644 ( 
.A(n_2587),
.B(n_322),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2609),
.B(n_322),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_2624),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2578),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2577),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2625),
.A2(n_323),
.B1(n_324),
.B2(n_326),
.Y(n_2649)
);

NAND4xp75_ASAP7_75t_L g2650 ( 
.A(n_2640),
.B(n_327),
.C(n_328),
.D(n_329),
.Y(n_2650)
);

NOR2x1p5_ASAP7_75t_L g2651 ( 
.A(n_2586),
.B(n_327),
.Y(n_2651)
);

NOR2x1_ASAP7_75t_L g2652 ( 
.A(n_2599),
.B(n_328),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2606),
.B(n_329),
.Y(n_2653)
);

NOR3xp33_ASAP7_75t_L g2654 ( 
.A(n_2594),
.B(n_330),
.C(n_331),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2601),
.B(n_330),
.Y(n_2655)
);

NOR2x1_ASAP7_75t_L g2656 ( 
.A(n_2631),
.B(n_331),
.Y(n_2656)
);

XNOR2xp5_ASAP7_75t_L g2657 ( 
.A(n_2596),
.B(n_332),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2580),
.Y(n_2658)
);

AOI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2602),
.A2(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_2659)
);

NOR2xp67_ASAP7_75t_L g2660 ( 
.A(n_2636),
.B(n_333),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2616),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2601),
.B(n_335),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2621),
.Y(n_2663)
);

INVxp33_ASAP7_75t_L g2664 ( 
.A(n_2583),
.Y(n_2664)
);

NAND3xp33_ASAP7_75t_L g2665 ( 
.A(n_2584),
.B(n_336),
.C(n_337),
.Y(n_2665)
);

NOR2x1_ASAP7_75t_L g2666 ( 
.A(n_2641),
.B(n_336),
.Y(n_2666)
);

NOR2x1_ASAP7_75t_L g2667 ( 
.A(n_2635),
.B(n_337),
.Y(n_2667)
);

AND2x4_ASAP7_75t_L g2668 ( 
.A(n_2623),
.B(n_2628),
.Y(n_2668)
);

NAND2x1p5_ASAP7_75t_L g2669 ( 
.A(n_2620),
.B(n_338),
.Y(n_2669)
);

OAI211xp5_ASAP7_75t_L g2670 ( 
.A1(n_2633),
.A2(n_339),
.B(n_340),
.C(n_341),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2637),
.Y(n_2671)
);

OAI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2590),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_2672)
);

NAND4xp75_ASAP7_75t_L g2673 ( 
.A(n_2614),
.B(n_342),
.C(n_343),
.D(n_344),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2632),
.B(n_344),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2610),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2626),
.B(n_346),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2629),
.Y(n_2677)
);

NOR2x1_ASAP7_75t_L g2678 ( 
.A(n_2627),
.B(n_346),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2618),
.B(n_347),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2603),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2600),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2595),
.B(n_2617),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2597),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2604),
.Y(n_2684)
);

NAND2x1p5_ASAP7_75t_L g2685 ( 
.A(n_2598),
.B(n_348),
.Y(n_2685)
);

AND2x2_ASAP7_75t_SL g2686 ( 
.A(n_2612),
.B(n_348),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2579),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2585),
.Y(n_2688)
);

AOI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2611),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_2689)
);

NAND4xp75_ASAP7_75t_L g2690 ( 
.A(n_2619),
.B(n_349),
.C(n_351),
.D(n_352),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2608),
.B(n_353),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2638),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_2692)
);

NOR2x1_ASAP7_75t_L g2693 ( 
.A(n_2582),
.B(n_2588),
.Y(n_2693)
);

XNOR2xp5_ASAP7_75t_L g2694 ( 
.A(n_2591),
.B(n_354),
.Y(n_2694)
);

NOR2x1_ASAP7_75t_L g2695 ( 
.A(n_2630),
.B(n_355),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2593),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2655),
.Y(n_2697)
);

NOR2x2_ASAP7_75t_L g2698 ( 
.A(n_2650),
.B(n_2622),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2674),
.B(n_2607),
.Y(n_2699)
);

NAND4xp25_ASAP7_75t_SL g2700 ( 
.A(n_2689),
.B(n_2659),
.C(n_2670),
.D(n_2678),
.Y(n_2700)
);

NOR3xp33_ASAP7_75t_SL g2701 ( 
.A(n_2658),
.B(n_2645),
.C(n_2665),
.Y(n_2701)
);

NOR4xp25_ASAP7_75t_L g2702 ( 
.A(n_2663),
.B(n_2634),
.C(n_2615),
.D(n_2589),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_2643),
.B(n_2605),
.Y(n_2703)
);

NAND4xp75_ASAP7_75t_L g2704 ( 
.A(n_2660),
.B(n_2613),
.C(n_2592),
.D(n_360),
.Y(n_2704)
);

OAI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2657),
.A2(n_358),
.B(n_359),
.Y(n_2705)
);

AND3x4_ASAP7_75t_L g2706 ( 
.A(n_2656),
.B(n_362),
.C(n_363),
.Y(n_2706)
);

NOR3xp33_ASAP7_75t_L g2707 ( 
.A(n_2680),
.B(n_362),
.C(n_363),
.Y(n_2707)
);

NOR4xp25_ASAP7_75t_L g2708 ( 
.A(n_2646),
.B(n_364),
.C(n_366),
.D(n_367),
.Y(n_2708)
);

NOR4xp25_ASAP7_75t_L g2709 ( 
.A(n_2648),
.B(n_366),
.C(n_367),
.D(n_368),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2662),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2669),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2668),
.B(n_368),
.Y(n_2712)
);

NAND4xp25_ASAP7_75t_L g2713 ( 
.A(n_2679),
.B(n_369),
.C(n_370),
.D(n_371),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_L g2714 ( 
.A(n_2693),
.B(n_369),
.C(n_370),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2668),
.B(n_371),
.Y(n_2715)
);

NOR2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2642),
.B(n_372),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2690),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2685),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2651),
.B(n_373),
.Y(n_2719)
);

NAND3xp33_ASAP7_75t_SL g2720 ( 
.A(n_2644),
.B(n_373),
.C(n_374),
.Y(n_2720)
);

NAND2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2695),
.B(n_374),
.Y(n_2721)
);

NOR3xp33_ASAP7_75t_L g2722 ( 
.A(n_2687),
.B(n_2681),
.C(n_2682),
.Y(n_2722)
);

NOR3x1_ASAP7_75t_L g2723 ( 
.A(n_2673),
.B(n_375),
.C(n_376),
.Y(n_2723)
);

NAND5xp2_ASAP7_75t_L g2724 ( 
.A(n_2664),
.B(n_375),
.C(n_376),
.D(n_377),
.E(n_378),
.Y(n_2724)
);

NAND3xp33_ASAP7_75t_L g2725 ( 
.A(n_2654),
.B(n_377),
.C(n_379),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2653),
.B(n_380),
.Y(n_2726)
);

XNOR2xp5_ASAP7_75t_L g2727 ( 
.A(n_2686),
.B(n_380),
.Y(n_2727)
);

AOI32xp33_ASAP7_75t_L g2728 ( 
.A1(n_2652),
.A2(n_381),
.A3(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_2728)
);

AND2x2_ASAP7_75t_SL g2729 ( 
.A(n_2676),
.B(n_381),
.Y(n_2729)
);

NOR3xp33_ASAP7_75t_SL g2730 ( 
.A(n_2684),
.B(n_384),
.C(n_385),
.Y(n_2730)
);

NOR5xp2_ASAP7_75t_L g2731 ( 
.A(n_2661),
.B(n_386),
.C(n_387),
.D(n_389),
.E(n_390),
.Y(n_2731)
);

NOR2x1_ASAP7_75t_L g2732 ( 
.A(n_2667),
.B(n_386),
.Y(n_2732)
);

OAI211xp5_ASAP7_75t_SL g2733 ( 
.A1(n_2666),
.A2(n_390),
.B(n_391),
.C(n_392),
.Y(n_2733)
);

OAI221xp5_ASAP7_75t_L g2734 ( 
.A1(n_2649),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.C(n_395),
.Y(n_2734)
);

AOI211xp5_ASAP7_75t_SL g2735 ( 
.A1(n_2675),
.A2(n_393),
.B(n_394),
.C(n_395),
.Y(n_2735)
);

INVx2_ASAP7_75t_SL g2736 ( 
.A(n_2694),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2691),
.B(n_396),
.Y(n_2737)
);

NAND3xp33_ASAP7_75t_SL g2738 ( 
.A(n_2683),
.B(n_398),
.C(n_399),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2672),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2732),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2736),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2727),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2721),
.Y(n_2743)
);

AND3x4_ASAP7_75t_L g2744 ( 
.A(n_2722),
.B(n_2688),
.C(n_2671),
.Y(n_2744)
);

BUFx2_ASAP7_75t_L g2745 ( 
.A(n_2719),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2701),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2697),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_2699),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2710),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2711),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2716),
.Y(n_2751)
);

CKINVDCx16_ASAP7_75t_R g2752 ( 
.A(n_2720),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2712),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2730),
.Y(n_2754)
);

NOR2xp67_ASAP7_75t_L g2755 ( 
.A(n_2724),
.B(n_2738),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2715),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2718),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2705),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2706),
.Y(n_2759)
);

O2A1O1Ixp5_ASAP7_75t_SL g2760 ( 
.A1(n_2739),
.A2(n_2677),
.B(n_2692),
.C(n_2647),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2735),
.Y(n_2761)
);

OAI221xp5_ASAP7_75t_L g2762 ( 
.A1(n_2728),
.A2(n_2696),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_2762)
);

BUFx2_ASAP7_75t_L g2763 ( 
.A(n_2698),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2717),
.Y(n_2764)
);

BUFx2_ASAP7_75t_L g2765 ( 
.A(n_2737),
.Y(n_2765)
);

AOI221xp5_ASAP7_75t_SL g2766 ( 
.A1(n_2713),
.A2(n_398),
.B1(n_401),
.B2(n_402),
.C(n_403),
.Y(n_2766)
);

INVx1_ASAP7_75t_SL g2767 ( 
.A(n_2729),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2703),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2759),
.Y(n_2769)
);

INVx1_ASAP7_75t_SL g2770 ( 
.A(n_2740),
.Y(n_2770)
);

AOI322xp5_ASAP7_75t_L g2771 ( 
.A1(n_2761),
.A2(n_2714),
.A3(n_2726),
.B1(n_2707),
.B2(n_2723),
.C1(n_2700),
.C2(n_2702),
.Y(n_2771)
);

AOI222xp33_ASAP7_75t_L g2772 ( 
.A1(n_2763),
.A2(n_2733),
.B1(n_2725),
.B2(n_2734),
.C1(n_2704),
.C2(n_2731),
.Y(n_2772)
);

NOR2x1_ASAP7_75t_L g2773 ( 
.A(n_2743),
.B(n_2709),
.Y(n_2773)
);

OAI211xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2751),
.A2(n_2708),
.B(n_404),
.C(n_405),
.Y(n_2774)
);

AOI32xp33_ASAP7_75t_L g2775 ( 
.A1(n_2767),
.A2(n_403),
.A3(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_2775)
);

AOI221xp5_ASAP7_75t_L g2776 ( 
.A1(n_2762),
.A2(n_408),
.B1(n_409),
.B2(n_411),
.C(n_412),
.Y(n_2776)
);

O2A1O1Ixp33_ASAP7_75t_L g2777 ( 
.A1(n_2753),
.A2(n_408),
.B(n_411),
.C(n_412),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2741),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2745),
.Y(n_2779)
);

NOR3xp33_ASAP7_75t_L g2780 ( 
.A(n_2752),
.B(n_414),
.C(n_415),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2748),
.Y(n_2781)
);

AOI322xp5_ASAP7_75t_L g2782 ( 
.A1(n_2766),
.A2(n_416),
.A3(n_417),
.B1(n_418),
.B2(n_419),
.C1(n_420),
.C2(n_421),
.Y(n_2782)
);

AOI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2746),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_2783)
);

AOI322xp5_ASAP7_75t_L g2784 ( 
.A1(n_2756),
.A2(n_2742),
.A3(n_2754),
.B1(n_2764),
.B2(n_2768),
.C1(n_2750),
.C2(n_2757),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2759),
.Y(n_2785)
);

INVxp67_ASAP7_75t_L g2786 ( 
.A(n_2748),
.Y(n_2786)
);

INVxp67_ASAP7_75t_L g2787 ( 
.A(n_2748),
.Y(n_2787)
);

OAI211xp5_ASAP7_75t_L g2788 ( 
.A1(n_2747),
.A2(n_421),
.B(n_422),
.C(n_423),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2781),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2779),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2786),
.A2(n_2744),
.B1(n_2749),
.B2(n_2755),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2780),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2774),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2773),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2769),
.Y(n_2795)
);

OAI22x1_ASAP7_75t_L g2796 ( 
.A1(n_2787),
.A2(n_2770),
.B1(n_2785),
.B2(n_2758),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2788),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2776),
.A2(n_2759),
.B1(n_2765),
.B2(n_2760),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2777),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2772),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_2800)
);

OAI221xp5_ASAP7_75t_R g2801 ( 
.A1(n_2798),
.A2(n_2784),
.B1(n_2771),
.B2(n_2783),
.C(n_2782),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2790),
.A2(n_2778),
.B1(n_2775),
.B2(n_427),
.Y(n_2802)
);

NAND3xp33_ASAP7_75t_SL g2803 ( 
.A(n_2791),
.B(n_425),
.C(n_426),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2800),
.B(n_425),
.Y(n_2804)
);

AOI22xp33_ASAP7_75t_L g2805 ( 
.A1(n_2794),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2805)
);

NOR3xp33_ASAP7_75t_L g2806 ( 
.A(n_2795),
.B(n_428),
.C(n_429),
.Y(n_2806)
);

CKINVDCx20_ASAP7_75t_R g2807 ( 
.A(n_2789),
.Y(n_2807)
);

XNOR2x1_ASAP7_75t_L g2808 ( 
.A(n_2796),
.B(n_429),
.Y(n_2808)
);

OR2x6_ASAP7_75t_L g2809 ( 
.A(n_2804),
.B(n_2797),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2808),
.B(n_2793),
.Y(n_2810)
);

XNOR2x1_ASAP7_75t_L g2811 ( 
.A(n_2802),
.B(n_2792),
.Y(n_2811)
);

OA21x2_ASAP7_75t_L g2812 ( 
.A1(n_2806),
.A2(n_2799),
.B(n_431),
.Y(n_2812)
);

OAI22x1_ASAP7_75t_L g2813 ( 
.A1(n_2801),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_2813)
);

NAND3xp33_ASAP7_75t_L g2814 ( 
.A(n_2807),
.B(n_2805),
.C(n_2803),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_SL g2815 ( 
.A1(n_2813),
.A2(n_430),
.B1(n_433),
.B2(n_434),
.Y(n_2815)
);

OAI22xp5_ASAP7_75t_SL g2816 ( 
.A1(n_2814),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_2816)
);

XNOR2xp5_ASAP7_75t_L g2817 ( 
.A(n_2811),
.B(n_435),
.Y(n_2817)
);

OAI21xp33_ASAP7_75t_L g2818 ( 
.A1(n_2810),
.A2(n_436),
.B(n_437),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2812),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2819),
.A2(n_2809),
.B(n_2815),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2817),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_2821)
);

NOR3xp33_ASAP7_75t_L g2822 ( 
.A(n_2820),
.B(n_2818),
.C(n_2816),
.Y(n_2822)
);

AOI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2822),
.A2(n_2821),
.B1(n_440),
.B2(n_441),
.Y(n_2823)
);

OAI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2822),
.A2(n_439),
.B1(n_440),
.B2(n_442),
.Y(n_2824)
);

NOR2xp67_ASAP7_75t_L g2825 ( 
.A(n_2823),
.B(n_442),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2825),
.Y(n_2826)
);

AOI221xp5_ASAP7_75t_L g2827 ( 
.A1(n_2826),
.A2(n_2824),
.B1(n_444),
.B2(n_445),
.C(n_446),
.Y(n_2827)
);

AOI221x1_ASAP7_75t_L g2828 ( 
.A1(n_2827),
.A2(n_443),
.B1(n_444),
.B2(n_446),
.C(n_447),
.Y(n_2828)
);

AOI211xp5_ASAP7_75t_L g2829 ( 
.A1(n_2828),
.A2(n_447),
.B(n_448),
.C(n_449),
.Y(n_2829)
);


endmodule