module real_jpeg_3150_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_48),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_54),
.B1(n_56),
.B2(n_78),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_78),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_78),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_68),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_5),
.B(n_27),
.C(n_74),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_5),
.B(n_73),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_32),
.C(n_35),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_110),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_44),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_5),
.B(n_39),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_110),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_54),
.B1(n_56),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_67),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_14),
.A2(n_26),
.B1(n_59),
.B2(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_14),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_15),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_53),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_53),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_115),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_21),
.B(n_115),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_83),
.C(n_92),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_22),
.B(n_83),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_49),
.B1(n_81),
.B2(n_82),
.Y(n_22)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_24),
.B(n_40),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_25),
.Y(n_175)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_27),
.A2(n_29),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_27),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_30),
.A2(n_37),
.B1(n_39),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_30),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_30),
.B(n_158),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_34),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_34),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_34),
.A2(n_176),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_34),
.A2(n_119),
.B1(n_155),
.B2(n_196),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_35),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_35),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_39),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_41),
.A2(n_44),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_41),
.A2(n_110),
.B(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_43),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_42),
.A2(n_43),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_42),
.A2(n_43),
.B1(n_113),
.B2(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_42),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_42),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_42),
.A2(n_43),
.B1(n_188),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_43),
.A2(n_152),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_43),
.B(n_166),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_44),
.A2(n_165),
.B(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_45),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_69),
.B2(n_70),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_51),
.B(n_69),
.C(n_81),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_60),
.A3(n_62),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_110),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_54),
.A2(n_109),
.B(n_110),
.C(n_134),
.Y(n_171)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_58),
.B(n_99),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_59),
.B(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_59),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_76),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_71),
.A2(n_72),
.B1(n_103),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_72),
.A2(n_76),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_72),
.A2(n_102),
.B1(n_103),
.B2(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_77),
.Y(n_104)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_91),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_92),
.A2(n_93),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.C(n_105),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_243)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_103),
.A2(n_104),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_105),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_138),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_119),
.A2(n_157),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_137),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_239),
.B(n_253),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_182),
.B(n_238),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_167),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_143),
.B(n_167),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.C(n_159),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_144),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_148),
.C(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_159),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_168),
.B(n_179),
.C(n_181),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_177),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_173),
.C(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_233),
.B(n_237),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_223),
.B(n_232),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_205),
.B(n_222),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_199),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_197),
.B2(n_198),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_216),
.B(n_221),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_214),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_219),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_229),
.C(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_248),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);


endmodule