module fake_jpeg_24440_n_260 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_18),
.B1(n_15),
.B2(n_27),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_26),
.B(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_15),
.B1(n_17),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_54),
.B1(n_18),
.B2(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_0),
.B(n_1),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_54),
.B1(n_57),
.B2(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_64),
.B1(n_73),
.B2(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_28),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_70),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_24),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_49),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_36),
.B1(n_19),
.B2(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_83),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_43),
.A3(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_85),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_56),
.C(n_45),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_56),
.B1(n_47),
.B2(n_46),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_95),
.B1(n_78),
.B2(n_64),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_52),
.A3(n_34),
.B1(n_35),
.B2(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_52),
.C(n_35),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_97),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_47),
.B1(n_49),
.B2(n_23),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_29),
.B1(n_28),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_70),
.B1(n_29),
.B2(n_71),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_118),
.B(n_121),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_123),
.B(n_101),
.C(n_85),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_124),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_60),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_122),
.B1(n_93),
.B2(n_95),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_68),
.B1(n_60),
.B2(n_75),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_67),
.B(n_74),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_77),
.B1(n_76),
.B2(n_69),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_0),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_83),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_87),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_138),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_99),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_108),
.B(n_124),
.C(n_122),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_144),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_86),
.B1(n_123),
.B2(n_111),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_93),
.C(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_110),
.C(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_79),
.B1(n_92),
.B2(n_66),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_86),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_92),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_125),
.B1(n_117),
.B2(n_107),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_151),
.B1(n_170),
.B2(n_140),
.Y(n_171)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_109),
.B1(n_119),
.B2(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_168),
.C(n_169),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_137),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_100),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_23),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_120),
.B1(n_109),
.B2(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_166),
.B1(n_140),
.B2(n_142),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_111),
.B(n_115),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_131),
.B(n_136),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_89),
.C(n_90),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_89),
.C(n_90),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_149),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_178),
.B1(n_182),
.B2(n_170),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_142),
.B(n_130),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_180),
.B(n_190),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_138),
.C(n_144),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_187),
.C(n_188),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_142),
.B1(n_141),
.B2(n_134),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_22),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_128),
.B1(n_71),
.B2(n_79),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_67),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.Y(n_191)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_71),
.B1(n_65),
.B2(n_66),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_150),
.B1(n_152),
.B2(n_164),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_65),
.C(n_67),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_1),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_12),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_165),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_194),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_201),
.B(n_181),
.C(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_165),
.C(n_160),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_205),
.C(n_174),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_12),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_22),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_210),
.C(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_177),
.C(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_216),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_175),
.B(n_184),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_196),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

AO221x1_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_202),
.B1(n_206),
.B2(n_4),
.C(n_5),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_173),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_194),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_222),
.C(n_230),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_195),
.C(n_205),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_212),
.B(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_193),
.C(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_2),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_217),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_207),
.B1(n_216),
.B2(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_238),
.C(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_212),
.C(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_11),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_224),
.A3(n_228),
.B1(n_222),
.B2(n_230),
.C1(n_9),
.C2(n_11),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_246),
.B(n_238),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_11),
.C(n_10),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_245),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_237),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_2),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_249),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_252),
.B(n_3),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_10),
.B(n_9),
.C(n_5),
.Y(n_252)
);

OAI321xp33_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_244),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_3),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_256),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_258)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_257),
.A3(n_254),
.B1(n_8),
.B2(n_4),
.C(n_3),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_8),
.Y(n_260)
);


endmodule