module fake_jpeg_13393_n_572 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_572);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_572;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_45),
.Y(n_127)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_27),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g167 ( 
.A(n_75),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_85),
.Y(n_117)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_86),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_32),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_107),
.Y(n_176)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

BUFx12f_ASAP7_75t_SL g96 ( 
.A(n_31),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_96),
.A2(n_16),
.B(n_17),
.Y(n_142)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_103),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_39),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_114),
.B(n_137),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_24),
.B1(n_47),
.B2(n_45),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_21),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_127),
.B(n_159),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_63),
.A2(n_64),
.B1(n_80),
.B2(n_86),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_132),
.A2(n_99),
.B1(n_83),
.B2(n_102),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_41),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_41),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_109),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_15),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_63),
.B(n_29),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_148),
.B(n_157),
.Y(n_217)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_149),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_29),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_56),
.B(n_42),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_100),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_42),
.B(n_46),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_40),
.Y(n_188)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_89),
.B(n_46),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_170),
.B(n_47),
.Y(n_233)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_98),
.A2(n_49),
.B1(n_43),
.B2(n_47),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_62),
.B1(n_108),
.B2(n_105),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_182),
.B(n_183),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_209),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_188),
.A2(n_227),
.B(n_229),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_224),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_19),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_210),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_197),
.Y(n_252)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_192),
.Y(n_279)
);

FAx1_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_73),
.CI(n_71),
.CON(n_193),
.SN(n_193)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_193),
.A2(n_213),
.B(n_231),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_79),
.B1(n_95),
.B2(n_72),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_195),
.A2(n_199),
.B1(n_232),
.B2(n_235),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_198),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_218),
.Y(n_253)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

CKINVDCx9p33_ASAP7_75t_R g205 ( 
.A(n_153),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_205),
.Y(n_261)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_40),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_61),
.C(n_104),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_212),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_116),
.B(n_57),
.C(n_58),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_223),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_126),
.C(n_115),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_124),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_21),
.B1(n_38),
.B2(n_20),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_117),
.B(n_20),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_177),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_236),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_38),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_176),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_156),
.B(n_15),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_33),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_135),
.B(n_33),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_233),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_174),
.A2(n_33),
.B1(n_43),
.B2(n_49),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_87),
.B1(n_82),
.B2(n_69),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_171),
.A2(n_43),
.B1(n_90),
.B2(n_102),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_240),
.B(n_163),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_110),
.B1(n_88),
.B2(n_59),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_161),
.B(n_0),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_237),
.B(n_3),
.Y(n_277)
);

HAxp5_ASAP7_75t_SL g238 ( 
.A(n_142),
.B(n_0),
.CON(n_238),
.SN(n_238)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_238),
.B(n_179),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_146),
.B(n_0),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_242),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_244),
.Y(n_292)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_111),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_238),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_199),
.A2(n_169),
.B1(n_132),
.B2(n_128),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_257),
.A2(n_270),
.B1(n_283),
.B2(n_286),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_140),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_223),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_193),
.A2(n_131),
.B1(n_178),
.B2(n_164),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_281),
.B1(n_293),
.B2(n_239),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_268),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_269),
.A2(n_221),
.B(n_196),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_188),
.A2(n_128),
.B1(n_178),
.B2(n_131),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_277),
.B(n_198),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_205),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_285),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_211),
.A2(n_164),
.B1(n_154),
.B2(n_138),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_189),
.A2(n_154),
.B1(n_151),
.B2(n_158),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_216),
.B(n_166),
.C(n_118),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_295),
.C(n_239),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_190),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_214),
.A2(n_147),
.B1(n_158),
.B2(n_133),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_193),
.A2(n_158),
.B1(n_133),
.B2(n_166),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_291),
.B1(n_207),
.B2(n_181),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_235),
.A2(n_210),
.B1(n_194),
.B2(n_217),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_229),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_229),
.B(n_166),
.C(n_118),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_299),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_308),
.C(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_291),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_201),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_300),
.B(n_301),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_249),
.B(n_236),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_206),
.B1(n_225),
.B2(n_184),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_303),
.A2(n_316),
.B1(n_266),
.B2(n_261),
.Y(n_368)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_227),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_245),
.B(n_227),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_277),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_312),
.B(n_321),
.Y(n_353)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_203),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_267),
.C(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_244),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_288),
.C(n_270),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_323),
.Y(n_370)
);

AO22x1_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_204),
.B1(n_200),
.B2(n_186),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_324),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_253),
.B(n_196),
.Y(n_321)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_246),
.A2(n_204),
.A3(n_212),
.B1(n_208),
.B2(n_180),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_251),
.B(n_192),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_326),
.B(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_200),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_292),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_330),
.B(n_331),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_224),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_275),
.B(n_185),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_332),
.B(n_334),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_268),
.B(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_336),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_264),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_252),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_337),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_5),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_339),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_6),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_323),
.A2(n_269),
.B(n_248),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_340),
.B(n_329),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_267),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_358),
.C(n_377),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_SL g399 ( 
.A1(n_345),
.A2(n_354),
.B(n_360),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_319),
.B1(n_314),
.B2(n_296),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_347),
.A2(n_356),
.B1(n_352),
.B2(n_346),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_336),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_278),
.B(n_286),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_281),
.B1(n_265),
.B2(n_257),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_282),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_255),
.B(n_258),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_311),
.B(n_318),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_297),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_368),
.A2(n_371),
.B1(n_333),
.B2(n_276),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_309),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_303),
.A2(n_266),
.B1(n_263),
.B2(n_256),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_304),
.A2(n_272),
.B(n_258),
.C(n_294),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_294),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_380),
.A2(n_383),
.B(n_401),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_361),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_381),
.B(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_357),
.B(n_338),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_385),
.B(n_388),
.Y(n_423)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_357),
.B(n_308),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_389),
.A2(n_392),
.B1(n_406),
.B2(n_409),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_390),
.B(n_391),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_327),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_299),
.B1(n_324),
.B2(n_300),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_394),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_395),
.B(n_343),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_279),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_402),
.Y(n_414)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

INVx13_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_407),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_333),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_279),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_259),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_404),
.Y(n_418)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_259),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_365),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_356),
.A2(n_370),
.B1(n_350),
.B2(n_341),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_336),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_351),
.C(n_358),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_370),
.A2(n_333),
.B1(n_325),
.B2(n_322),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_370),
.A2(n_350),
.B1(n_340),
.B2(n_346),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_410),
.A2(n_373),
.B1(n_349),
.B2(n_366),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_367),
.B(n_259),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_411),
.B(n_365),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_250),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_383),
.A2(n_360),
.B(n_362),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_417),
.B(n_287),
.Y(n_470)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_421),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_351),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_432),
.C(n_433),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_345),
.B(n_354),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_424),
.A2(n_436),
.B(n_401),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_368),
.B1(n_371),
.B2(n_349),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_431),
.Y(n_448)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_407),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_384),
.B(n_377),
.C(n_369),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_373),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_440),
.C(n_378),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_376),
.B(n_366),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_389),
.A2(n_372),
.B1(n_359),
.B2(n_276),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_412),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_273),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_273),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_408),
.C(n_394),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_381),
.B(n_264),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_444),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_445),
.A2(n_382),
.B1(n_379),
.B2(n_409),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_449),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_470),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_395),
.C(n_406),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_453),
.C(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_452),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_393),
.C(n_397),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_378),
.Y(n_454)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_387),
.C(n_386),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_458),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_463),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_461),
.A2(n_443),
.B(n_415),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_423),
.B(n_404),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g486 ( 
.A(n_462),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_419),
.Y(n_463)
);

FAx1_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_398),
.CI(n_287),
.CON(n_464),
.SN(n_464)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_472),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_417),
.C(n_434),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_438),
.C(n_443),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_436),
.A2(n_271),
.B1(n_247),
.B2(n_250),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_468),
.A2(n_439),
.B1(n_427),
.B2(n_430),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_434),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_469),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_418),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_466),
.Y(n_476)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_271),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_473),
.B(n_421),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_413),
.B(n_7),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_426),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_454),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_475),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_476),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_453),
.Y(n_477)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_477),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_428),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_481),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_452),
.B1(n_472),
.B2(n_463),
.Y(n_503)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_489),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_448),
.A2(n_431),
.B1(n_445),
.B2(n_416),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_492),
.B1(n_457),
.B2(n_460),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_448),
.A2(n_416),
.B1(n_420),
.B2(n_438),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_447),
.A2(n_430),
.B1(n_438),
.B2(n_437),
.Y(n_493)
);

XNOR2x1_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_490),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_496),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_467),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_473),
.B(n_459),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_446),
.B(n_425),
.C(n_437),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_450),
.C(n_456),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_490),
.B(n_488),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_493),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_502),
.A2(n_488),
.B1(n_480),
.B2(n_489),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_503),
.A2(n_491),
.B1(n_485),
.B2(n_478),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_505),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_484),
.A2(n_456),
.B1(n_465),
.B2(n_464),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_492),
.A2(n_451),
.B1(n_464),
.B2(n_461),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_506),
.A2(n_478),
.B1(n_485),
.B2(n_487),
.Y(n_527)
);

BUFx12_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_508),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_470),
.C(n_474),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_516),
.C(n_517),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_514),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_425),
.C(n_415),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_483),
.B(n_7),
.C(n_9),
.Y(n_517)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_502),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_522),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_482),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_521),
.A2(n_515),
.B1(n_508),
.B2(n_504),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_495),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_527),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_525),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_510),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_531),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_507),
.Y(n_543)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_500),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_499),
.A2(n_486),
.B1(n_494),
.B2(n_10),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_533),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_506),
.A2(n_499),
.B1(n_513),
.B2(n_512),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_523),
.A2(n_510),
.B1(n_515),
.B2(n_508),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_534),
.A2(n_541),
.B1(n_543),
.B2(n_7),
.Y(n_553)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_536),
.Y(n_551)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_519),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_539),
.B(n_540),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_533),
.B(n_511),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_509),
.B1(n_517),
.B2(n_507),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_530),
.A2(n_521),
.B(n_528),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_528),
.B(n_522),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_537),
.Y(n_547)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_548),
.A2(n_544),
.B(n_545),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_520),
.C(n_529),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_552),
.Y(n_559)
);

AOI31xp67_ASAP7_75t_L g550 ( 
.A1(n_534),
.A2(n_518),
.A3(n_524),
.B(n_494),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_550),
.B(n_551),
.C(n_538),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_7),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_553),
.B(n_556),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_546),
.B(n_9),
.Y(n_555)
);

CKINVDCx14_ASAP7_75t_R g558 ( 
.A(n_555),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_9),
.C(n_10),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g563 ( 
.A1(n_557),
.A2(n_560),
.B(n_554),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_564),
.Y(n_567)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_561),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_555),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_558),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_566),
.A2(n_562),
.B(n_556),
.Y(n_568)
);

AOI322xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_558),
.A3(n_567),
.B1(n_12),
.B2(n_13),
.C1(n_10),
.C2(n_11),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_11),
.B(n_13),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_13),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_13),
.Y(n_572)
);


endmodule