module fake_jpeg_25308_n_309 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_12),
.Y(n_38)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_11),
.B1(n_14),
.B2(n_20),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_11),
.B1(n_28),
.B2(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_25),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_41),
.C(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_44),
.B1(n_38),
.B2(n_39),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_38),
.B1(n_30),
.B2(n_40),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_91),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_38),
.C(n_50),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_32),
.C(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_74),
.B1(n_36),
.B2(n_30),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_93),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_49),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_33),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_100),
.B(n_26),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_11),
.B1(n_33),
.B2(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_53),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_77),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_135),
.C(n_118),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_97),
.B1(n_88),
.B2(n_84),
.Y(n_138)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_120),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_76),
.B(n_1),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_77),
.B1(n_37),
.B2(n_42),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_29),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_121),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_26),
.Y(n_118)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_29),
.B(n_13),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_129),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_74),
.B1(n_72),
.B2(n_78),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_82),
.B1(n_84),
.B2(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_133),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_57),
.B(n_59),
.C(n_74),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_26),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_78),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_127),
.B1(n_131),
.B2(n_42),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_86),
.C(n_90),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_139),
.B(n_171),
.C(n_19),
.Y(n_200)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_143),
.Y(n_179)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_148),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_162),
.B(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_21),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_154),
.B(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_103),
.B1(n_72),
.B2(n_78),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_118),
.B1(n_132),
.B2(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_109),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_62),
.B1(n_52),
.B2(n_56),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_134),
.B1(n_110),
.B2(n_106),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_55),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_26),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_114),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_19),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_121),
.B(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_115),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_122),
.B(n_112),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_186),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_193),
.B1(n_198),
.B2(n_35),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_117),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_178),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_105),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_138),
.B1(n_153),
.B2(n_141),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_105),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_151),
.Y(n_205)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_113),
.B1(n_120),
.B2(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_143),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_153),
.B(n_137),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_133),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_152),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_18),
.B1(n_21),
.B2(n_30),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_157),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_137),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_171),
.C(n_161),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_160),
.C(n_140),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_183),
.C(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_223),
.B1(n_176),
.B2(n_179),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_168),
.B(n_165),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_168),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_199),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_149),
.B(n_18),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_35),
.B1(n_28),
.B2(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_230),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_174),
.B1(n_182),
.B2(n_190),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_244),
.B1(n_225),
.B2(n_239),
.Y(n_258)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

XOR2x1_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_184),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_212),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_194),
.B1(n_195),
.B2(n_175),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_241),
.B1(n_28),
.B2(n_43),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_195),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_181),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_198),
.B1(n_184),
.B2(n_35),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_17),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_224),
.B1(n_210),
.B2(n_202),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_203),
.C(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_249),
.C(n_254),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_247),
.B(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_213),
.C(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

BUFx12_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_221),
.C(n_206),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_253),
.Y(n_265)
);

BUFx12_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

OAI322xp33_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_215),
.A3(n_17),
.B1(n_15),
.B2(n_19),
.C1(n_23),
.C2(n_20),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_28),
.CI(n_15),
.CON(n_260),
.SN(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_259),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_242),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_7),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_237),
.C(n_225),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_270),
.C(n_19),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_15),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_251),
.C(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_15),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_247),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_278),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_247),
.B1(n_251),
.B2(n_43),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_20),
.Y(n_275)
);

NOR2x1_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_43),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_20),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_17),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_282),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_23),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_23),
.C(n_15),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_262),
.B(n_268),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_6),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_10),
.C2(n_7),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_289),
.B1(n_282),
.B2(n_276),
.Y(n_295)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_261),
.C(n_270),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_15),
.C(n_17),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_6),
.Y(n_294)
);

AOI31xp33_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_296),
.A3(n_298),
.B(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_0),
.C(n_3),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_3),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_285),
.B(n_298),
.Y(n_301)
);

XOR2x2_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

OAI311xp33_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_286),
.A3(n_294),
.B1(n_7),
.C1(n_8),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_303),
.B(n_297),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_0),
.A3(n_4),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_304),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_8),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_9),
.B(n_0),
.Y(n_309)
);


endmodule