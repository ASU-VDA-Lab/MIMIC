module fake_jpeg_29256_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_62),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_46),
.B1(n_37),
.B2(n_40),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_42),
.B2(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_37),
.B1(n_43),
.B2(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_76),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_47),
.B(n_51),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_79),
.Y(n_84)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_39),
.B1(n_18),
.B2(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_42),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_19),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_89),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_17),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_90),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_7),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_5),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_6),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_80),
.C(n_72),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_71),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_92),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_99),
.B1(n_86),
.B2(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_102),
.B1(n_85),
.B2(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_82),
.B(n_94),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_22),
.B1(n_9),
.B2(n_11),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_23),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_87),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.C1(n_20),
.C2(n_21),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_25),
.C(n_26),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_27),
.B(n_30),
.C(n_31),
.D(n_7),
.Y(n_108)
);


endmodule