module fake_jpeg_480_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_59),
.Y(n_146)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_68),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_29),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_30),
.B1(n_52),
.B2(n_50),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_16),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_109),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_72),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_74),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_76),
.Y(n_204)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_78),
.Y(n_151)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_80),
.Y(n_179)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_125),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_0),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_90),
.A2(n_97),
.B(n_105),
.Y(n_158)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_0),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_100),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_101),
.B(n_103),
.Y(n_205)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_1),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_21),
.B(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_52),
.B1(n_50),
.B2(n_41),
.Y(n_149)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_22),
.Y(n_117)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_34),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_127),
.A2(n_150),
.B1(n_172),
.B2(n_71),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_43),
.B1(n_35),
.B2(n_34),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g275 ( 
.A1(n_133),
.A2(n_173),
.B(n_189),
.C(n_135),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_134),
.A2(n_149),
.B1(n_206),
.B2(n_73),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_57),
.B(n_56),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_139),
.B(n_141),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_57),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_152),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_38),
.B1(n_41),
.B2(n_24),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_56),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_79),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_159),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_84),
.B(n_54),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_48),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_181),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_67),
.B(n_36),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_163),
.B(n_164),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_104),
.B(n_36),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_80),
.B(n_24),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_169),
.B(n_178),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_48),
.B1(n_46),
.B2(n_28),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_80),
.B(n_46),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_60),
.B(n_43),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_5),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_88),
.B(n_121),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_6),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_61),
.B(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_69),
.A2(n_40),
.B1(n_8),
.B2(n_9),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_92),
.B(n_7),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_136),
.A2(n_128),
.A3(n_148),
.B1(n_158),
.B2(n_129),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_211),
.B(n_217),
.Y(n_318)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_213),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_127),
.A2(n_111),
.B1(n_75),
.B2(n_108),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_214),
.A2(n_215),
.B1(n_223),
.B2(n_243),
.Y(n_301)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_216),
.Y(n_303)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_221),
.B(n_231),
.Y(n_332)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_158),
.A2(n_64),
.B1(n_100),
.B2(n_89),
.Y(n_223)
);

AO22x2_ASAP7_75t_L g224 ( 
.A1(n_133),
.A2(n_115),
.B1(n_98),
.B2(n_85),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_224),
.A2(n_275),
.B(n_214),
.C(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_226),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_140),
.A2(n_83),
.B1(n_76),
.B2(n_78),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_227),
.A2(n_229),
.B1(n_250),
.B2(n_258),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_40),
.B1(n_8),
.B2(n_10),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_228),
.A2(n_254),
.B1(n_268),
.B2(n_271),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_156),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_10),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_131),
.A2(n_177),
.B1(n_132),
.B2(n_168),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_233),
.A2(n_256),
.B1(n_257),
.B2(n_277),
.Y(n_327)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_142),
.Y(n_238)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_239),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_152),
.A2(n_126),
.B1(n_145),
.B2(n_175),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_240),
.A2(n_253),
.B1(n_262),
.B2(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_241),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_166),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_11),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_244),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_251),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_138),
.A2(n_16),
.B1(n_11),
.B2(n_15),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_252),
.B(n_260),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_187),
.A2(n_15),
.B1(n_210),
.B2(n_208),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_205),
.A2(n_146),
.B1(n_179),
.B2(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_197),
.B(n_154),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_269),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g256 ( 
.A1(n_210),
.A2(n_208),
.B1(n_207),
.B2(n_204),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_166),
.A2(n_207),
.B1(n_204),
.B2(n_198),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_192),
.A2(n_170),
.B1(n_126),
.B2(n_146),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_258),
.Y(n_291)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_144),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_259),
.B(n_261),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_160),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_145),
.A2(n_198),
.B1(n_182),
.B2(n_144),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_130),
.A2(n_143),
.B1(n_203),
.B2(n_195),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_265),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_267),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_179),
.A2(n_200),
.B1(n_191),
.B2(n_130),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_195),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_270),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_160),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_216),
.Y(n_287)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_276),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_191),
.A2(n_200),
.B1(n_153),
.B2(n_194),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_275),
.A2(n_278),
.B1(n_224),
.B2(n_253),
.Y(n_317)
);

AO22x1_ASAP7_75t_SL g276 ( 
.A1(n_194),
.A2(n_167),
.B1(n_153),
.B2(n_173),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_135),
.A2(n_186),
.B1(n_189),
.B2(n_161),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_135),
.A2(n_186),
.B1(n_189),
.B2(n_161),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_186),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_244),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_150),
.A2(n_134),
.B1(n_149),
.B2(n_181),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_280),
.A2(n_235),
.B1(n_238),
.B2(n_248),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_287),
.B(n_308),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_246),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_292),
.C(n_296),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_322),
.B(n_311),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_242),
.C(n_221),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_245),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_217),
.B1(n_212),
.B2(n_211),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_299),
.A2(n_310),
.B1(n_316),
.B2(n_322),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_234),
.A2(n_231),
.B(n_244),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_286),
.B(n_312),
.Y(n_342)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_281),
.A2(n_263),
.A3(n_264),
.B1(n_218),
.B2(n_232),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_269),
.A2(n_233),
.B1(n_231),
.B2(n_255),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_224),
.A2(n_265),
.B1(n_239),
.B2(n_236),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_237),
.B(n_251),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_323),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_222),
.B(n_225),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_321),
.B(n_330),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_224),
.A2(n_256),
.B1(n_259),
.B2(n_220),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_213),
.B(n_252),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_219),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_314),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_261),
.B(n_273),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_327),
.B1(n_301),
.B2(n_300),
.Y(n_347)
);

OAI21xp33_ASAP7_75t_SL g336 ( 
.A1(n_311),
.A2(n_275),
.B(n_276),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_336),
.A2(n_350),
.B(n_368),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_316),
.A2(n_275),
.B1(n_249),
.B2(n_226),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_230),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_341),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_270),
.B1(n_267),
.B2(n_247),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_344),
.B1(n_347),
.B2(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_247),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_360),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_289),
.A2(n_317),
.B1(n_327),
.B2(n_331),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_345),
.A2(n_358),
.B1(n_344),
.B2(n_349),
.Y(n_405)
);

BUFx12f_ASAP7_75t_SL g346 ( 
.A(n_291),
.Y(n_346)
);

NAND2x1_ASAP7_75t_SL g403 ( 
.A(n_346),
.B(n_348),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_325),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_328),
.Y(n_351)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_351),
.Y(n_375)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_295),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_284),
.A2(n_292),
.B1(n_318),
.B2(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_318),
.A2(n_299),
.B1(n_332),
.B2(n_293),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_359),
.A2(n_293),
.B1(n_315),
.B2(n_285),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_332),
.C(n_318),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_342),
.C(n_334),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_290),
.B(n_330),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_366),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_298),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_307),
.B(n_332),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_369),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_289),
.A2(n_306),
.B(n_314),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_329),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_290),
.B(n_326),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_373),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_372),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_333),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_356),
.C(n_335),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_368),
.A2(n_315),
.B(n_313),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_387),
.B(n_341),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_302),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_381),
.B(n_361),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_403),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_337),
.A2(n_303),
.B(n_285),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_373),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_402),
.Y(n_408)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_352),
.Y(n_394)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_345),
.A2(n_304),
.B1(n_324),
.B2(n_309),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_396),
.B1(n_401),
.B2(n_336),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_343),
.A2(n_309),
.B1(n_302),
.B2(n_283),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_372),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_372),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_343),
.A2(n_282),
.B1(n_283),
.B2(n_305),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_398),
.A2(n_357),
.B1(n_371),
.B2(n_369),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_347),
.A2(n_282),
.B1(n_305),
.B2(n_297),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_303),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_405),
.A2(n_297),
.B1(n_364),
.B2(n_380),
.Y(n_434)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_407),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_428),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_413),
.C(n_424),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_416),
.B(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_359),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_354),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_432),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_403),
.A2(n_346),
.B(n_339),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_400),
.Y(n_418)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_418),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_358),
.B(n_350),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_426),
.B1(n_429),
.B2(n_388),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_399),
.A2(n_344),
.B(n_350),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_367),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_379),
.A2(n_344),
.B1(n_358),
.B2(n_350),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_425),
.A2(n_427),
.B1(n_430),
.B2(n_382),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_379),
.A2(n_338),
.B1(n_353),
.B2(n_363),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_353),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_338),
.A3(n_348),
.B1(n_365),
.B2(n_354),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_405),
.A2(n_340),
.B1(n_348),
.B2(n_366),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_374),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_431),
.A2(n_434),
.B1(n_401),
.B2(n_432),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_403),
.A2(n_346),
.B(n_348),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_355),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_385),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_399),
.B(n_380),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_435),
.A2(n_441),
.B(n_411),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_437),
.A2(n_444),
.B1(n_454),
.B2(n_459),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_438),
.A2(n_446),
.B(n_420),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_393),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_457),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_415),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_453),
.C(n_458),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_431),
.A2(n_387),
.B(n_386),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_395),
.B1(n_404),
.B2(n_385),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_449),
.B(n_433),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_393),
.C(n_383),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_451),
.C(n_423),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_396),
.C(n_398),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_390),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_429),
.A2(n_406),
.B1(n_375),
.B2(n_376),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_389),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_389),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_375),
.B1(n_376),
.B2(n_394),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_470),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_445),
.A2(n_444),
.B1(n_454),
.B2(n_438),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_461),
.A2(n_477),
.B1(n_478),
.B2(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_462),
.B(n_476),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_464),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_416),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_465),
.Y(n_481)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_455),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_430),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_408),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_428),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_475),
.C(n_442),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_422),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_452),
.B(n_408),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_445),
.A2(n_422),
.B1(n_412),
.B2(n_434),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_443),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_486),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_461),
.A2(n_446),
.B1(n_441),
.B2(n_435),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_483),
.A2(n_465),
.B1(n_464),
.B2(n_407),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_451),
.C(n_450),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_486),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_448),
.C(n_457),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_489),
.A2(n_471),
.B1(n_488),
.B2(n_483),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_449),
.C(n_436),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_491),
.C(n_463),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_436),
.C(n_422),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_482),
.A2(n_472),
.B(n_470),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_493),
.B(n_499),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_494),
.A2(n_504),
.B1(n_481),
.B2(n_414),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_500),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_485),
.A2(n_460),
.B(n_473),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_501),
.B(n_417),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_498),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_452),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_479),
.A2(n_447),
.B(n_477),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_474),
.B(n_469),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_468),
.C(n_471),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_492),
.C(n_480),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_490),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_507),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_487),
.Y(n_509)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_509),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_480),
.C(n_414),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_513),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_497),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

AOI322xp5_ASAP7_75t_L g515 ( 
.A1(n_510),
.A2(n_496),
.A3(n_417),
.B1(n_419),
.B2(n_504),
.C1(n_495),
.C2(n_397),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_511),
.B1(n_507),
.B2(n_392),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_505),
.A2(n_419),
.B(n_384),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_517),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_384),
.Y(n_518)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_518),
.Y(n_525)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_510),
.B(n_508),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_524),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_520),
.B(n_518),
.Y(n_526)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_526),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_529),
.Y(n_531)
);

AOI21xp33_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_530),
.B(n_519),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_527),
.B1(n_521),
.B2(n_525),
.Y(n_533)
);


endmodule