module fake_jpeg_22469_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_22),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_40),
.B1(n_49),
.B2(n_17),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_43),
.B1(n_16),
.B2(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_14),
.B1(n_24),
.B2(n_21),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_16),
.B1(n_15),
.B2(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_19),
.B1(n_27),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_60),
.Y(n_84)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_59),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_16),
.B1(n_19),
.B2(n_26),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_51),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_67),
.B1(n_38),
.B2(n_25),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_51),
.B1(n_56),
.B2(n_68),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_43),
.B(n_50),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_77),
.B(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_85),
.B1(n_55),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_81),
.B1(n_57),
.B2(n_54),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_36),
.B(n_31),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_64),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_49),
.B1(n_48),
.B2(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_94),
.B1(n_46),
.B2(n_29),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_97),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_93),
.B(n_84),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_64),
.B1(n_67),
.B2(n_61),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_64),
.A3(n_30),
.B1(n_35),
.B2(n_34),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_103),
.Y(n_122)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_52),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_44),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_80),
.A3(n_70),
.B1(n_75),
.B2(n_86),
.C1(n_83),
.C2(n_73),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_72),
.B(n_83),
.C(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_114),
.B1(n_119),
.B2(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_76),
.C(n_73),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_103),
.C(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_20),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_48),
.B(n_52),
.C(n_44),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_123),
.B1(n_99),
.B2(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_88),
.B1(n_96),
.B2(n_58),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_97),
.B1(n_95),
.B2(n_90),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_108),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_0),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_135),
.C(n_136),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_138),
.B1(n_22),
.B2(n_20),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_35),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_34),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_29),
.B1(n_44),
.B2(n_33),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_22),
.B1(n_34),
.B2(n_33),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_145),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_120),
.B(n_107),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_147),
.B(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_112),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_116),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_153),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_116),
.B(n_33),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_116),
.A3(n_22),
.B1(n_20),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_133),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_155),
.B1(n_137),
.B2(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_135),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_160),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_136),
.B(n_6),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_164),
.C(n_7),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_6),
.C(n_10),
.D(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_155),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_5),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_152),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_153),
.B(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_174),
.C(n_178),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_149),
.B1(n_148),
.B2(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_154),
.C(n_156),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_178),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_0),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_149),
.C(n_1),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_185),
.C(n_9),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_184),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_4),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_0),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_7),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_176),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_192),
.B(n_193),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_177),
.B1(n_8),
.B2(n_3),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_4),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.C(n_8),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_182),
.B(n_11),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_11),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_193),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_2),
.B(n_195),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_193),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_2),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_2),
.B(n_203),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);


endmodule