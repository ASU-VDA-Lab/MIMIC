module real_jpeg_31269_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_86),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_0),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_0),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_0),
.B(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_2),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_2),
.B(n_166),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_2),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_2),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_3),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_3),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_3),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_3),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_3),
.B(n_310),
.Y(n_309)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_6),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_9),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_9),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_9),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_141),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_9),
.B(n_166),
.Y(n_165)
);

NAND2x1p5_ASAP7_75t_L g198 ( 
.A(n_9),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_10),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_10),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_10),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_10),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_11),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_11),
.B(n_108),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_11),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_11),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_91),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_12),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_12),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_13),
.Y(n_401)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_16),
.Y(n_298)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_16),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_17),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_17),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_17),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_17),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_17),
.B(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_17),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_93),
.B(n_274),
.C(n_428),
.D(n_437),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_236),
.C(n_264),
.Y(n_24)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_205),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_171),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_27),
.B(n_171),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_99),
.C(n_132),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_29),
.B(n_100),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_70),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_30),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_44),
.B(n_69),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_31),
.B(n_45),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_34),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_39),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_39),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_104),
.C(n_105),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_40),
.A2(n_41),
.B1(n_287),
.B2(n_288),
.Y(n_379)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_41),
.B(n_198),
.C(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_58),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_52),
.B(n_57),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_47),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_47),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_47),
.A2(n_150),
.B1(n_329),
.B2(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_96),
.C(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_50),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_56),
.Y(n_233)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_57),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_58),
.Y(n_355)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_61),
.A2(n_97),
.B1(n_165),
.B2(n_261),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_L g437 ( 
.A(n_61),
.B(n_179),
.C(n_261),
.Y(n_437)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_88),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_71),
.B(n_173),
.C(n_174),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.C(n_84),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_72),
.B(n_169),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.C(n_79),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_79),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_73),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_73),
.A2(n_137),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_73),
.B(n_187),
.C(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_75),
.B(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_82),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_82),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_83),
.A2(n_84),
.B1(n_85),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_93),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_84),
.A2(n_85),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_85),
.B(n_218),
.C(n_222),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_96),
.B(n_123),
.C(n_126),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_120),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_119),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_119),
.C(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_107),
.B(n_110),
.C(n_113),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_107),
.A2(n_165),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_107),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_107),
.B(n_235),
.C(n_261),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_109)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_140),
.C(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_110),
.A2(n_118),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_117),
.Y(n_340)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_123),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_123),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_123),
.B(n_333),
.C(n_336),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_123),
.A2(n_200),
.B1(n_336),
.B2(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_125),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_128),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_132),
.B(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_151),
.C(n_167),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_134),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_147),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_135),
.B(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_139),
.A2(n_147),
.B1(n_148),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_139),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_140),
.A2(n_196),
.B1(n_197),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_140),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_197),
.C(n_229),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_140),
.B(n_144),
.Y(n_344)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_151),
.A2(n_152),
.B1(n_167),
.B2(n_168),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.C(n_165),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_153),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_159),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_154),
.B(n_156),
.Y(n_305)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_155),
.Y(n_321)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_159),
.B(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_160),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g331 ( 
.A(n_160),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_162),
.B(n_165),
.Y(n_300)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_190),
.C(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

XOR2x1_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_179),
.A2(n_220),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_188),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_200),
.C(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_197),
.B(n_379),
.Y(n_378)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_207),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_209),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_215),
.C(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_224),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_234),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g429 ( 
.A1(n_237),
.A2(n_265),
.B(n_430),
.C(n_434),
.D(n_435),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_262),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_238),
.B(n_262),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_257),
.B2(n_258),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_255),
.C(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_266),
.B(n_267),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_269),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_357),
.B(n_419),
.C(n_420),
.D(n_427),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_347),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_277),
.B(n_347),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.C(n_322),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g384 ( 
.A(n_279),
.B(n_283),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_303),
.Y(n_283)
);

AO22x2_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_294),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_290),
.B1(n_294),
.B2(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_352),
.C(n_353),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_312),
.Y(n_303)
);

XOR2x2_ASAP7_75t_L g380 ( 
.A(n_304),
.B(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_306),
.A2(n_307),
.B1(n_312),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_319),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_314),
.B1(n_319),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_384),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_341),
.C(n_345),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.C(n_332),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_333),
.B(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_345),
.Y(n_361)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_354),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_385),
.B(n_418),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_383),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_383),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.C(n_380),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_SL g387 ( 
.A(n_363),
.B(n_380),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_375),
.C(n_377),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_364),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.C(n_371),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_378),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_415),
.Y(n_388)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_397),
.C(n_412),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.C(n_409),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_425),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.C(n_424),
.Y(n_421)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.C(n_433),
.Y(n_430)
);


endmodule