module fake_netlist_1_6950_n_1369 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1369);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1369;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g338 ( .A(n_298), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_199), .Y(n_339) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_92), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_269), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_156), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_49), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_260), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_307), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_101), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_161), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_7), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_139), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_140), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_163), .Y(n_352) );
NOR2xp67_ASAP7_75t_L g353 ( .A(n_71), .B(n_159), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_261), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_1), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_46), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_327), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_152), .Y(n_358) );
CKINVDCx16_ASAP7_75t_R g359 ( .A(n_33), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_34), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_214), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_11), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_278), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_283), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_336), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_282), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_319), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_32), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_228), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_169), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_78), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_219), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_258), .B(n_225), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_21), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_58), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_7), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_243), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_59), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_81), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_277), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_16), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_276), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_247), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_32), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_176), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_312), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_244), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_223), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_206), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_204), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_184), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_313), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_170), .Y(n_396) );
CKINVDCx14_ASAP7_75t_R g397 ( .A(n_52), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_136), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_270), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_149), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_193), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_227), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_154), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_187), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_188), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_218), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_210), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_63), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_165), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_232), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_5), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_56), .B(n_191), .Y(n_412) );
BUFx8_ASAP7_75t_SL g413 ( .A(n_302), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_19), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_41), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_162), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_189), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_245), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_288), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_289), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_45), .Y(n_421) );
INVxp33_ASAP7_75t_SL g422 ( .A(n_242), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_74), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_92), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_162), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_161), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_10), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_186), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_182), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_54), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_190), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_96), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_238), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_68), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_140), .B(n_284), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_100), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_65), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_80), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_23), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_133), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_259), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_205), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_1), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_220), .Y(n_444) );
INVxp33_ASAP7_75t_L g445 ( .A(n_286), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_217), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_201), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_263), .Y(n_448) );
BUFx5_ASAP7_75t_L g449 ( .A(n_267), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_123), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_275), .Y(n_451) );
INVxp33_ASAP7_75t_SL g452 ( .A(n_231), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_209), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_139), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_142), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_167), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_81), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_60), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_297), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_134), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_271), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_36), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_133), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_274), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_123), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_265), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_70), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_180), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_196), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_117), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_303), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_155), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_83), .Y(n_474) );
INVxp33_ASAP7_75t_SL g475 ( .A(n_268), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_68), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_40), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_53), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_6), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_43), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_337), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_43), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_234), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_121), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_154), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_324), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_118), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_226), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_49), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_86), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_122), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_251), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_27), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_175), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_90), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_317), .Y(n_496) );
INVxp33_ASAP7_75t_SL g497 ( .A(n_95), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_66), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_299), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_249), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_301), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_230), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_79), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_266), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_8), .Y(n_505) );
CKINVDCx14_ASAP7_75t_R g506 ( .A(n_221), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_183), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_240), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_156), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_77), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_246), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_106), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_148), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_166), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_160), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_213), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_300), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_60), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_413), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_365), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_365), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_365), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_445), .B(n_0), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_356), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_347), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_417), .B(n_2), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_397), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_417), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_365), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_417), .B(n_6), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_449), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_449), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_485), .B(n_9), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_389), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_445), .B(n_9), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_397), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_438), .B(n_12), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_389), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_389), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_372), .B(n_13), .Y(n_540) );
INVx6_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
AND2x6_ASAP7_75t_L g542 ( .A(n_446), .B(n_385), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_413), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_408), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_449), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_389), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_502), .B(n_13), .Y(n_547) );
BUFx8_ASAP7_75t_L g548 ( .A(n_449), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_449), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_515), .B(n_14), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_449), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_420), .B(n_15), .Y(n_552) );
BUFx3_ASAP7_75t_L g553 ( .A(n_446), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_354), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_340), .B(n_17), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_372), .B(n_18), .Y(n_557) );
INVx5_ASAP7_75t_L g558 ( .A(n_541), .Y(n_558) );
OR2x6_ASAP7_75t_L g559 ( .A(n_524), .B(n_353), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_523), .A2(n_497), .B1(n_362), .B2(n_414), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_526), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_553), .B(n_339), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_526), .B(n_385), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_520), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_531), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_531), .Y(n_567) );
INVx4_ASAP7_75t_L g568 ( .A(n_526), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_532), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_526), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_528), .B(n_393), .Y(n_571) );
BUFx3_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_530), .A2(n_343), .B1(n_349), .B2(n_348), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_532), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_530), .A2(n_350), .B1(n_355), .B2(n_351), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_520), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_553), .B(n_368), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_548), .Y(n_579) );
INVx4_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_545), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_523), .B(n_506), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_545), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_528), .B(n_393), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_535), .B(n_506), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_430), .B1(n_359), .B2(n_406), .Y(n_587) );
INVx8_ASAP7_75t_L g588 ( .A(n_540), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_548), .B(n_404), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
INVx4_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_520), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_519), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_541), .B(n_395), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_525), .B(n_391), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_555), .B(n_361), .Y(n_596) );
NAND2xp33_ASAP7_75t_R g597 ( .A(n_556), .B(n_357), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_541), .B(n_395), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_525), .B(n_418), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_540), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_520), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_540), .B(n_418), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
NAND2xp33_ASAP7_75t_L g604 ( .A(n_579), .B(n_542), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_596), .B(n_552), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_582), .B(n_557), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_582), .B(n_557), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_562), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_582), .B(n_543), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_557), .B1(n_533), .B2(n_536), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_586), .B(n_563), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_572), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_586), .B(n_537), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_572), .B(n_369), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_562), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_572), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_560), .A2(n_527), .B1(n_524), .B2(n_536), .C(n_415), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_562), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_578), .B(n_366), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_579), .B(n_369), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_562), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_568), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_570), .Y(n_624) );
OR2x6_ASAP7_75t_L g625 ( .A(n_588), .B(n_550), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_570), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_590), .B(n_415), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_570), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_578), .B(n_568), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_593), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_588), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_597), .A2(n_448), .B1(n_394), .B2(n_554), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_588), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_570), .Y(n_634) );
NOR2x1p5_ASAP7_75t_L g635 ( .A(n_560), .B(n_400), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_588), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_568), .B(n_410), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_580), .B(n_410), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_589), .B(n_357), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_580), .B(n_492), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_588), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_583), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_580), .B(n_492), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_583), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_564), .B(n_422), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_583), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_574), .A2(n_376), .B1(n_381), .B2(n_352), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_587), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_600), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_590), .B(n_496), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_599), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_576), .B(n_501), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_576), .B(n_501), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_587), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_600), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_600), .B(n_452), .Y(n_659) );
NOR2x1p5_ASAP7_75t_L g660 ( .A(n_600), .B(n_383), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_600), .A2(n_424), .B1(n_454), .B2(n_443), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_595), .B(n_603), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_603), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_603), .A2(n_467), .B1(n_472), .B2(n_455), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_566), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_602), .A2(n_479), .B1(n_503), .B2(n_476), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_591), .B(n_475), .Y(n_667) );
O2A1O1Ixp5_ASAP7_75t_L g668 ( .A1(n_602), .A2(n_547), .B(n_451), .C(n_367), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_566), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_SL g670 ( .A1(n_567), .A2(n_402), .B(n_435), .C(n_549), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_591), .B(n_345), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_591), .B(n_363), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_591), .B(n_382), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_567), .A2(n_542), .B1(n_551), .B2(n_549), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_569), .A2(n_542), .B1(n_551), .B2(n_358), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_575), .Y(n_677) );
AND2x6_ASAP7_75t_SL g678 ( .A(n_559), .B(n_360), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_577), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_581), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_594), .B(n_542), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_558), .B(n_399), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_638), .B(n_558), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_654), .B(n_598), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_606), .A2(n_598), .B(n_584), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_609), .Y(n_686) );
INVx4_ASAP7_75t_L g687 ( .A(n_633), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_609), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_585), .B(n_571), .C(n_380), .Y(n_689) );
NAND2x2_ASAP7_75t_L g690 ( .A(n_635), .B(n_559), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_615), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_638), .B(n_558), .Y(n_692) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_607), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_611), .B(n_559), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_624), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_608), .A2(n_559), .B1(n_542), .B2(n_585), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_627), .B(n_375), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_652), .A2(n_374), .B(n_341), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_608), .A2(n_436), .B1(n_478), .B2(n_423), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_633), .B(n_613), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_614), .B(n_518), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_625), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_608), .A2(n_436), .B1(n_478), .B2(n_423), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_625), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_631), .B(n_558), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_651), .B(n_493), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_642), .B(n_493), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_607), .A2(n_344), .B(n_338), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_624), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_627), .B(n_377), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_616), .A2(n_364), .B(n_346), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_626), .Y(n_713) );
BUFx10_ASAP7_75t_L g714 ( .A(n_660), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_644), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_626), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_612), .A2(n_398), .B(n_403), .C(n_387), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_616), .A2(n_371), .B(n_370), .Y(n_718) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_625), .Y(n_719) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_632), .B(n_512), .Y(n_720) );
BUFx3_ASAP7_75t_L g721 ( .A(n_669), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_657), .A2(n_416), .B(n_425), .C(n_411), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_605), .B(n_512), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_619), .A2(n_378), .B(n_373), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_621), .B(n_426), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_625), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_619), .A2(n_384), .B(n_379), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_622), .A2(n_388), .B(n_386), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_678), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_650), .B(n_421), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_628), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_662), .A2(n_427), .B(n_434), .C(n_432), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_669), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_618), .B(n_487), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_659), .B(n_437), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_628), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_665), .A2(n_439), .B(n_450), .C(n_440), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_622), .Y(n_738) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_680), .Y(n_739) );
INVx3_ASAP7_75t_L g740 ( .A(n_623), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_637), .A2(n_392), .B(n_390), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_665), .B(n_457), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_634), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_648), .B(n_458), .Y(n_744) );
AOI21x1_ASAP7_75t_L g745 ( .A1(n_681), .A2(n_565), .B(n_561), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_653), .B(n_460), .Y(n_746) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_680), .Y(n_747) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_623), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_677), .A2(n_462), .B(n_465), .C(n_463), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_640), .A2(n_405), .B(n_401), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_677), .Y(n_751) );
NOR3xp33_ASAP7_75t_SL g752 ( .A(n_666), .B(n_466), .C(n_459), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_652), .B(n_474), .Y(n_753) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_655), .A2(n_477), .B1(n_482), .B2(n_480), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_647), .A2(n_409), .B(n_407), .Y(n_755) );
INVxp67_ASAP7_75t_L g756 ( .A(n_656), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_661), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_664), .B(n_484), .Y(n_758) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_658), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_667), .B(n_489), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_639), .B(n_468), .Y(n_761) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_658), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_634), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_647), .B(n_490), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_649), .A2(n_428), .B(n_419), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_649), .A2(n_431), .B(n_429), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_636), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_641), .B(n_469), .Y(n_768) );
BUFx3_ASAP7_75t_L g769 ( .A(n_645), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_629), .A2(n_441), .B(n_433), .Y(n_770) );
O2A1O1Ixp33_ASAP7_75t_L g771 ( .A1(n_670), .A2(n_509), .B(n_510), .C(n_505), .Y(n_771) );
O2A1O1Ixp5_ASAP7_75t_L g772 ( .A1(n_668), .A2(n_494), .B(n_499), .C(n_483), .Y(n_772) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_663), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_620), .B(n_544), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_643), .B(n_470), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_663), .A2(n_447), .B(n_444), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_646), .B(n_491), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g778 ( .A(n_671), .B(n_471), .Y(n_778) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_675), .A2(n_498), .B1(n_491), .B2(n_473), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_674), .A2(n_412), .B(n_498), .C(n_456), .Y(n_780) );
O2A1O1Ixp5_ASAP7_75t_L g781 ( .A1(n_672), .A2(n_494), .B(n_499), .C(n_483), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_673), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_604), .B(n_481), .Y(n_783) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_679), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_604), .A2(n_461), .B(n_453), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_682), .B(n_464), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_679), .B(n_504), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_630), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_606), .A2(n_488), .B(n_486), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_609), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_606), .A2(n_508), .B(n_507), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_654), .B(n_514), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_638), .B(n_511), .Y(n_793) );
AO21x2_ASAP7_75t_L g794 ( .A1(n_670), .A2(n_517), .B(n_516), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_654), .A2(n_473), .B1(n_495), .B2(n_342), .Y(n_795) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_660), .B(n_342), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_660), .B(n_342), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_609), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_606), .A2(n_592), .B(n_573), .Y(n_799) );
AO21x1_ASAP7_75t_L g800 ( .A1(n_606), .A2(n_592), .B(n_573), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_610), .B(n_342), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_654), .B(n_473), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g803 ( .A1(n_654), .A2(n_495), .B(n_513), .C(n_473), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_633), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_654), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_654), .B(n_495), .Y(n_806) );
O2A1O1Ixp33_ASAP7_75t_L g807 ( .A1(n_651), .A2(n_601), .B(n_592), .C(n_513), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_609), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g809 ( .A1(n_654), .A2(n_513), .B(n_495), .C(n_442), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_606), .A2(n_601), .B(n_577), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_654), .B(n_513), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_606), .A2(n_601), .B(n_577), .Y(n_812) );
BUFx3_ASAP7_75t_L g813 ( .A(n_630), .Y(n_813) );
AO32x1_ASAP7_75t_L g814 ( .A1(n_665), .A2(n_529), .A3(n_534), .B1(n_522), .B2(n_521), .Y(n_814) );
NAND3xp33_ASAP7_75t_SL g815 ( .A(n_630), .B(n_19), .C(n_20), .Y(n_815) );
AO32x2_ASAP7_75t_L g816 ( .A1(n_779), .A2(n_795), .A3(n_754), .B1(n_800), .B2(n_814), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_707), .B(n_22), .Y(n_817) );
O2A1O1Ixp33_ASAP7_75t_L g818 ( .A1(n_732), .A2(n_24), .B(n_22), .C(n_23), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_805), .Y(n_819) );
O2A1O1Ixp33_ASAP7_75t_L g820 ( .A1(n_717), .A2(n_26), .B(n_24), .C(n_25), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_753), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_810), .A2(n_577), .B(n_442), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_695), .A2(n_442), .B1(n_500), .B2(n_396), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_700), .B(n_28), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_812), .A2(n_577), .B(n_442), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_721), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_720), .A2(n_500), .B1(n_396), .B2(n_521), .Y(n_827) );
AOI21x1_ASAP7_75t_L g828 ( .A1(n_745), .A2(n_500), .B(n_396), .Y(n_828) );
BUFx10_ASAP7_75t_L g829 ( .A(n_797), .Y(n_829) );
NOR2x1_ASAP7_75t_SL g830 ( .A(n_703), .B(n_521), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_753), .Y(n_831) );
BUFx2_ASAP7_75t_L g832 ( .A(n_813), .Y(n_832) );
INVx6_ASAP7_75t_L g833 ( .A(n_714), .Y(n_833) );
AO31x2_ASAP7_75t_L g834 ( .A1(n_780), .A2(n_522), .A3(n_529), .B(n_521), .Y(n_834) );
OA21x2_ASAP7_75t_L g835 ( .A1(n_809), .A2(n_522), .B(n_521), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_799), .A2(n_577), .B(n_522), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_L g837 ( .A1(n_689), .A2(n_31), .B(n_29), .C(n_30), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_774), .A2(n_522), .B(n_529), .C(n_521), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_684), .A2(n_529), .B1(n_534), .B2(n_522), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_685), .A2(n_534), .B(n_529), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_714), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_L g842 ( .A1(n_737), .A2(n_31), .B(n_29), .C(n_30), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_764), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_691), .A2(n_534), .B1(n_538), .B2(n_529), .Y(n_844) );
AO31x2_ASAP7_75t_L g845 ( .A1(n_803), .A2(n_538), .A3(n_539), .B(n_534), .Y(n_845) );
BUFx3_ASAP7_75t_L g846 ( .A(n_788), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_797), .B(n_35), .Y(n_847) );
BUFx10_ASAP7_75t_L g848 ( .A(n_760), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_751), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_723), .B(n_708), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_757), .B(n_35), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_734), .B(n_36), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_756), .B(n_37), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_690), .A2(n_538), .B1(n_539), .B2(n_534), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_806), .A2(n_539), .B(n_538), .Y(n_855) );
AO32x2_ASAP7_75t_L g856 ( .A1(n_779), .A2(n_546), .A3(n_539), .B1(n_538), .B2(n_39), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_784), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g858 ( .A1(n_772), .A2(n_546), .B(n_539), .Y(n_858) );
O2A1O1Ixp33_ASAP7_75t_L g859 ( .A1(n_749), .A2(n_39), .B(n_37), .C(n_38), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_700), .B(n_42), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_751), .Y(n_861) );
INVx2_ASAP7_75t_SL g862 ( .A(n_796), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_704), .B(n_42), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_758), .A2(n_546), .B1(n_45), .B2(n_44), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_751), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_730), .B(n_46), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_770), .A2(n_171), .B(n_168), .Y(n_867) );
AO31x2_ASAP7_75t_L g868 ( .A1(n_795), .A2(n_50), .A3(n_47), .B(n_48), .Y(n_868) );
BUFx6f_ASAP7_75t_L g869 ( .A(n_693), .Y(n_869) );
INVx3_ASAP7_75t_L g870 ( .A(n_687), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_715), .B(n_50), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_789), .A2(n_173), .B(n_172), .Y(n_872) );
O2A1O1Ixp33_ASAP7_75t_L g873 ( .A1(n_722), .A2(n_55), .B(n_51), .C(n_54), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_811), .A2(n_177), .B(n_174), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_702), .B(n_55), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_703), .A2(n_58), .B1(n_56), .B2(n_57), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_764), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_705), .A2(n_61), .B1(n_57), .B2(n_59), .Y(n_878) );
AOI221x1_ASAP7_75t_L g879 ( .A1(n_815), .A2(n_62), .B1(n_64), .B2(n_65), .C(n_66), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_771), .A2(n_70), .B(n_67), .C(n_69), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_733), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_792), .A2(n_179), .B(n_178), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_802), .A2(n_185), .B(n_181), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_711), .B(n_72), .Y(n_884) );
O2A1O1Ixp33_ASAP7_75t_L g885 ( .A1(n_744), .A2(n_75), .B(n_73), .C(n_74), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_742), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_733), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_705), .A2(n_76), .B1(n_73), .B2(n_75), .Y(n_888) );
INVx3_ASAP7_75t_SL g889 ( .A(n_729), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_719), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_760), .A2(n_82), .B1(n_79), .B2(n_80), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_775), .A2(n_194), .B(n_192), .Y(n_892) );
A2O1A1Ixp33_ASAP7_75t_L g893 ( .A1(n_791), .A2(n_84), .B(n_82), .C(n_83), .Y(n_893) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_693), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_777), .A2(n_197), .B(n_195), .Y(n_895) );
A2O1A1Ixp33_ASAP7_75t_L g896 ( .A1(n_709), .A2(n_87), .B(n_85), .C(n_86), .Y(n_896) );
OAI211xp5_ASAP7_75t_L g897 ( .A1(n_697), .A2(n_89), .B(n_85), .C(n_88), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_793), .A2(n_200), .B(n_198), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_735), .A2(n_91), .B1(n_89), .B2(n_90), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_725), .B(n_91), .Y(n_900) );
O2A1O1Ixp33_ASAP7_75t_SL g901 ( .A1(n_742), .A2(n_233), .B(n_335), .C(n_334), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_725), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_801), .A2(n_93), .A3(n_94), .B(n_96), .Y(n_903) );
A2O1A1Ixp33_ASAP7_75t_L g904 ( .A1(n_712), .A2(n_97), .B(n_98), .C(n_99), .Y(n_904) );
AO31x2_ASAP7_75t_L g905 ( .A1(n_785), .A2(n_97), .A3(n_98), .B(n_99), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_746), .A2(n_100), .B1(n_102), .B2(n_103), .C(n_104), .Y(n_906) );
INVx4_ASAP7_75t_L g907 ( .A(n_726), .Y(n_907) );
OAI21xp5_ASAP7_75t_L g908 ( .A1(n_694), .A2(n_103), .B(n_104), .Y(n_908) );
A2O1A1Ixp33_ASAP7_75t_L g909 ( .A1(n_718), .A2(n_105), .B(n_106), .C(n_107), .Y(n_909) );
O2A1O1Ixp33_ASAP7_75t_SL g910 ( .A1(n_786), .A2(n_241), .B(n_333), .C(n_332), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_724), .A2(n_108), .B(n_109), .C(n_110), .Y(n_911) );
AOI22x1_ASAP7_75t_L g912 ( .A1(n_776), .A2(n_239), .B1(n_331), .B2(n_330), .Y(n_912) );
O2A1O1Ixp33_ASAP7_75t_SL g913 ( .A1(n_786), .A2(n_237), .B(n_329), .C(n_328), .Y(n_913) );
O2A1O1Ixp33_ASAP7_75t_SL g914 ( .A1(n_738), .A2(n_235), .B(n_326), .C(n_325), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_752), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_782), .Y(n_916) );
AO31x2_ASAP7_75t_L g917 ( .A1(n_727), .A2(n_111), .A3(n_112), .B(n_113), .Y(n_917) );
AOI31xp67_ASAP7_75t_L g918 ( .A1(n_814), .A2(n_236), .A3(n_323), .B(n_322), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_804), .B(n_112), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_699), .A2(n_203), .B(n_202), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_740), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_921) );
A2O1A1Ixp33_ASAP7_75t_L g922 ( .A1(n_728), .A2(n_114), .B(n_115), .C(n_116), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_740), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_733), .Y(n_924) );
INVx3_ASAP7_75t_L g925 ( .A(n_804), .Y(n_925) );
OA21x2_ASAP7_75t_L g926 ( .A1(n_781), .A2(n_208), .B(n_207), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_741), .A2(n_212), .B(n_211), .Y(n_927) );
OR2x2_ASAP7_75t_L g928 ( .A(n_739), .B(n_119), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_794), .A2(n_120), .B1(n_122), .B2(n_124), .Y(n_929) );
INVx3_ASAP7_75t_L g930 ( .A(n_748), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_686), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_739), .B(n_124), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_747), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_794), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_934) );
A2O1A1Ixp33_ASAP7_75t_L g935 ( .A1(n_750), .A2(n_125), .B(n_126), .C(n_127), .Y(n_935) );
A2O1A1Ixp33_ASAP7_75t_L g936 ( .A1(n_755), .A2(n_128), .B(n_129), .C(n_130), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_688), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_696), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_761), .A2(n_256), .B(n_320), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_748), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_940) );
AO21x1_ASAP7_75t_L g941 ( .A1(n_807), .A2(n_257), .B(n_318), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_710), .Y(n_942) );
O2A1O1Ixp33_ASAP7_75t_L g943 ( .A1(n_768), .A2(n_131), .B(n_132), .C(n_134), .Y(n_943) );
AOI21xp5_ASAP7_75t_L g944 ( .A1(n_713), .A2(n_255), .B(n_316), .Y(n_944) );
OR2x6_ASAP7_75t_L g945 ( .A(n_701), .B(n_131), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g946 ( .A1(n_765), .A2(n_254), .B(n_315), .Y(n_946) );
INVxp67_ASAP7_75t_L g947 ( .A(n_748), .Y(n_947) );
OAI21xp5_ASAP7_75t_L g948 ( .A1(n_766), .A2(n_253), .B(n_314), .Y(n_948) );
OAI221xp5_ASAP7_75t_L g949 ( .A1(n_778), .A2(n_132), .B1(n_135), .B2(n_136), .C(n_137), .Y(n_949) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_759), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g951 ( .A1(n_716), .A2(n_135), .B1(n_137), .B2(n_138), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_706), .B(n_141), .Y(n_952) );
AOI21xp5_ASAP7_75t_L g953 ( .A1(n_731), .A2(n_262), .B(n_311), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_736), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_743), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_763), .B(n_141), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_767), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_790), .A2(n_264), .B(n_309), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_769), .B(n_142), .Y(n_959) );
O2A1O1Ixp33_ASAP7_75t_L g960 ( .A1(n_683), .A2(n_692), .B(n_798), .C(n_808), .Y(n_960) );
INVxp67_ASAP7_75t_L g961 ( .A(n_787), .Y(n_961) );
OAI21xp5_ASAP7_75t_L g962 ( .A1(n_783), .A2(n_252), .B(n_308), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_762), .A2(n_250), .B(n_306), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g964 ( .A1(n_762), .A2(n_248), .B(n_305), .Y(n_964) );
A2O1A1Ixp33_ASAP7_75t_L g965 ( .A1(n_773), .A2(n_143), .B(n_144), .C(n_145), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_773), .A2(n_143), .B1(n_144), .B2(n_146), .C(n_147), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_773), .B(n_146), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_805), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_819), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_968), .Y(n_970) );
OR2x6_ASAP7_75t_L g971 ( .A(n_945), .B(n_149), .Y(n_971) );
AND2x4_ASAP7_75t_L g972 ( .A(n_886), .B(n_150), .Y(n_972) );
INVx1_ASAP7_75t_SL g973 ( .A(n_950), .Y(n_973) );
AO21x2_ASAP7_75t_L g974 ( .A1(n_858), .A2(n_273), .B(n_304), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_824), .B(n_150), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_821), .B(n_151), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_860), .B(n_153), .Y(n_977) );
BUFx8_ASAP7_75t_L g978 ( .A(n_832), .Y(n_978) );
INVx2_ASAP7_75t_L g979 ( .A(n_957), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_931), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_855), .A2(n_843), .B(n_831), .Y(n_981) );
A2O1A1Ixp33_ASAP7_75t_L g982 ( .A1(n_877), .A2(n_157), .B(n_158), .C(n_159), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_956), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_937), .Y(n_984) );
BUFx12f_ASAP7_75t_L g985 ( .A(n_833), .Y(n_985) );
INVx3_ASAP7_75t_L g986 ( .A(n_907), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_847), .Y(n_987) );
BUFx10_ASAP7_75t_L g988 ( .A(n_833), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_847), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_951), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_951), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_938), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_902), .B(n_164), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g994 ( .A1(n_827), .A2(n_215), .B(n_216), .C(n_222), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_871), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_848), .B(n_224), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_916), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_942), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_852), .B(n_229), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_866), .A2(n_279), .B1(n_280), .B2(n_281), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_945), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_869), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_954), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_955), .Y(n_1004) );
INVx3_ASAP7_75t_L g1005 ( .A(n_907), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_863), .B(n_285), .Y(n_1006) );
AOI21x1_ASAP7_75t_L g1007 ( .A1(n_932), .A2(n_287), .B(n_290), .Y(n_1007) );
NOR2x1_ASAP7_75t_R g1008 ( .A(n_846), .B(n_292), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_851), .B(n_293), .Y(n_1009) );
A2O1A1Ixp33_ASAP7_75t_L g1010 ( .A1(n_820), .A2(n_294), .B(n_295), .C(n_296), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_870), .B(n_890), .Y(n_1011) );
A2O1A1Ixp33_ASAP7_75t_L g1012 ( .A1(n_884), .A2(n_837), .B(n_818), .C(n_873), .Y(n_1012) );
OA21x2_ASAP7_75t_L g1013 ( .A1(n_823), .A2(n_962), .B(n_867), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_908), .Y(n_1014) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_869), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_915), .Y(n_1016) );
BUFx4f_ASAP7_75t_SL g1017 ( .A(n_841), .Y(n_1017) );
AOI21xp33_ASAP7_75t_L g1018 ( .A1(n_823), .A2(n_919), .B(n_885), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_900), .B(n_826), .Y(n_1019) );
A2O1A1Ixp33_ASAP7_75t_L g1020 ( .A1(n_943), .A2(n_859), .B(n_842), .C(n_952), .Y(n_1020) );
AOI21x1_ASAP7_75t_L g1021 ( .A1(n_926), .A2(n_839), .B(n_920), .Y(n_1021) );
A2O1A1Ixp33_ASAP7_75t_L g1022 ( .A1(n_959), .A2(n_880), .B(n_967), .C(n_934), .Y(n_1022) );
INVx4_ASAP7_75t_L g1023 ( .A(n_870), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_853), .B(n_923), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_864), .A2(n_906), .B1(n_891), .B2(n_899), .C(n_934), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_961), .B(n_849), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_928), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_890), .B(n_862), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_905), .Y(n_1029) );
AO21x2_ASAP7_75t_L g1030 ( .A1(n_872), .A2(n_927), .B(n_946), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_861), .B(n_865), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_881), .B(n_887), .Y(n_1032) );
INVx6_ASAP7_75t_L g1033 ( .A(n_829), .Y(n_1033) );
AO31x2_ASAP7_75t_L g1034 ( .A1(n_879), .A2(n_830), .A3(n_893), .B(n_874), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_905), .Y(n_1035) );
AO21x2_ASAP7_75t_L g1036 ( .A1(n_948), .A2(n_929), .B(n_901), .Y(n_1036) );
A2O1A1Ixp33_ASAP7_75t_L g1037 ( .A1(n_929), .A2(n_960), .B(n_897), .C(n_935), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_905), .Y(n_1038) );
OAI211xp5_ASAP7_75t_SL g1039 ( .A1(n_854), .A2(n_966), .B(n_949), .C(n_909), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_856), .Y(n_1040) );
OAI21xp5_ASAP7_75t_L g1041 ( .A1(n_882), .A2(n_892), .B(n_895), .Y(n_1041) );
CKINVDCx11_ASAP7_75t_R g1042 ( .A(n_894), .Y(n_1042) );
INVx3_ASAP7_75t_L g1043 ( .A(n_894), .Y(n_1043) );
NAND4xp25_ASAP7_75t_SL g1044 ( .A(n_921), .B(n_911), .C(n_904), .D(n_922), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_917), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_924), .B(n_925), .Y(n_1046) );
OAI21xp5_ASAP7_75t_L g1047 ( .A1(n_939), .A2(n_896), .B(n_936), .Y(n_1047) );
AOI21xp5_ASAP7_75t_L g1048 ( .A1(n_910), .A2(n_913), .B(n_914), .Y(n_1048) );
NAND3xp33_ASAP7_75t_L g1049 ( .A(n_965), .B(n_940), .C(n_878), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_925), .B(n_947), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_917), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_930), .B(n_933), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_876), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_888), .A2(n_912), .B1(n_844), .B2(n_835), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_917), .Y(n_1055) );
AOI22xp33_ASAP7_75t_SL g1056 ( .A1(n_926), .A2(n_835), .B1(n_856), .B2(n_816), .Y(n_1056) );
NAND4xp25_ASAP7_75t_L g1057 ( .A(n_898), .B(n_964), .C(n_963), .D(n_958), .Y(n_1057) );
OA21x2_ASAP7_75t_L g1058 ( .A1(n_883), .A2(n_953), .B(n_944), .Y(n_1058) );
OA21x2_ASAP7_75t_L g1059 ( .A1(n_816), .A2(n_834), .B(n_918), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_903), .Y(n_1060) );
AO21x1_ASAP7_75t_L g1061 ( .A1(n_816), .A2(n_903), .B(n_868), .Y(n_1061) );
INVx2_ASAP7_75t_SL g1062 ( .A(n_868), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_834), .B(n_845), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1064 ( .A1(n_845), .A2(n_836), .B(n_840), .Y(n_1064) );
AOI21xp5_ASAP7_75t_L g1065 ( .A1(n_845), .A2(n_836), .B(n_840), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_819), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_819), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_886), .B(n_805), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_886), .B(n_821), .Y(n_1069) );
AO21x2_ASAP7_75t_L g1070 ( .A1(n_840), .A2(n_858), .B(n_828), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_950), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_886), .B(n_805), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_822), .A2(n_825), .B(n_836), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_819), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_819), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_819), .Y(n_1076) );
A2O1A1Ixp33_ASAP7_75t_L g1077 ( .A1(n_875), .A2(n_850), .B(n_817), .C(n_886), .Y(n_1077) );
OR2x6_ASAP7_75t_L g1078 ( .A(n_945), .B(n_857), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_886), .B(n_821), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_848), .B(n_698), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_889), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_819), .Y(n_1082) );
OAI21x1_ASAP7_75t_SL g1083 ( .A1(n_908), .A2(n_830), .B(n_821), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1084 ( .A1(n_836), .A2(n_840), .B(n_825), .Y(n_1084) );
AOI21xp33_ASAP7_75t_L g1085 ( .A1(n_823), .A2(n_794), .B(n_850), .Y(n_1085) );
AO31x2_ASAP7_75t_L g1086 ( .A1(n_941), .A2(n_800), .A3(n_838), .B(n_825), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_819), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_819), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1040), .Y(n_1089) );
AOI21xp5_ASAP7_75t_SL g1090 ( .A1(n_971), .A2(n_1013), .B(n_972), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1068), .B(n_1072), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1068), .B(n_1072), .Y(n_1092) );
INVx4_ASAP7_75t_SL g1093 ( .A(n_971), .Y(n_1093) );
AO21x2_ASAP7_75t_L g1094 ( .A1(n_1064), .A2(n_1065), .B(n_1063), .Y(n_1094) );
CKINVDCx8_ASAP7_75t_R g1095 ( .A(n_1081), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_969), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g1097 ( .A1(n_1077), .A2(n_1012), .B(n_1022), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_970), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1023), .B(n_1078), .Y(n_1099) );
AOI21xp5_ASAP7_75t_SL g1100 ( .A1(n_1013), .A2(n_972), .B(n_1008), .Y(n_1100) );
INVx4_ASAP7_75t_R g1101 ( .A(n_1071), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1066), .Y(n_1102) );
OA21x2_ASAP7_75t_L g1103 ( .A1(n_1084), .A2(n_1061), .B(n_1035), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1069), .B(n_1079), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1067), .Y(n_1105) );
OA21x2_ASAP7_75t_L g1106 ( .A1(n_1029), .A2(n_1038), .B(n_1073), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1074), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1075), .Y(n_1108) );
OR2x6_ASAP7_75t_L g1109 ( .A(n_1078), .B(n_1001), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1076), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_980), .B(n_984), .Y(n_1111) );
BUFx3_ASAP7_75t_L g1112 ( .A(n_985), .Y(n_1112) );
OA21x2_ASAP7_75t_L g1113 ( .A1(n_1045), .A2(n_1055), .B(n_1051), .Y(n_1113) );
AND2x4_ASAP7_75t_L g1114 ( .A(n_1023), .B(n_986), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_992), .B(n_998), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1079), .B(n_979), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1117 ( .A(n_973), .B(n_975), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1082), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1003), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1087), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1088), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1004), .Y(n_1122) );
OR2x6_ASAP7_75t_L g1123 ( .A(n_1083), .B(n_990), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1080), .B(n_983), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_1026), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_991), .B(n_997), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1027), .B(n_977), .Y(n_1127) );
OR2x6_ASAP7_75t_L g1128 ( .A(n_987), .B(n_989), .Y(n_1128) );
AO21x2_ASAP7_75t_L g1129 ( .A1(n_1085), .A2(n_1070), .B(n_1036), .Y(n_1129) );
OA21x2_ASAP7_75t_L g1130 ( .A1(n_1085), .A2(n_1014), .B(n_1062), .Y(n_1130) );
AO21x2_ASAP7_75t_L g1131 ( .A1(n_1070), .A2(n_1036), .B(n_1021), .Y(n_1131) );
AO21x2_ASAP7_75t_L g1132 ( .A1(n_1018), .A2(n_1037), .B(n_1030), .Y(n_1132) );
INVxp67_ASAP7_75t_SL g1133 ( .A(n_1026), .Y(n_1133) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_1052), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_986), .B(n_1005), .Y(n_1135) );
OR2x2_ASAP7_75t_SL g1136 ( .A(n_1009), .B(n_1033), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_976), .B(n_993), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_993), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1060), .B(n_1019), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1019), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_995), .B(n_1006), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1005), .B(n_1011), .Y(n_1142) );
OA21x2_ASAP7_75t_L g1143 ( .A1(n_1047), .A2(n_1041), .B(n_1054), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1024), .B(n_1050), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1145 ( .A(n_1043), .B(n_1011), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_982), .B(n_1052), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1046), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1043), .B(n_1031), .Y(n_1148) );
BUFx3_ASAP7_75t_L g1149 ( .A(n_1042), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1046), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1031), .B(n_981), .Y(n_1151) );
AO21x2_ASAP7_75t_L g1152 ( .A1(n_1020), .A2(n_974), .B(n_1010), .Y(n_1152) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_1017), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1032), .B(n_999), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_1025), .A2(n_1044), .B1(n_1039), .B2(n_1053), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1032), .B(n_999), .Y(n_1156) );
OR2x6_ASAP7_75t_L g1157 ( .A(n_1002), .B(n_1015), .Y(n_1157) );
OA21x2_ASAP7_75t_L g1158 ( .A1(n_1007), .A2(n_1049), .B(n_1057), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1028), .B(n_1025), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1044), .B(n_1049), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1028), .Y(n_1161) );
BUFx4f_ASAP7_75t_SL g1162 ( .A(n_988), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1059), .B(n_1056), .Y(n_1163) );
AND2x4_ASAP7_75t_L g1164 ( .A(n_1034), .B(n_974), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g1165 ( .A1(n_1000), .A2(n_996), .B1(n_1057), .B2(n_1016), .C(n_994), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1034), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1034), .Y(n_1167) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_1058), .B(n_1086), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1068), .B(n_1072), .Y(n_1169) );
AOI21xp5_ASAP7_75t_L g1170 ( .A1(n_1048), .A2(n_1030), .B(n_1073), .Y(n_1170) );
OR2x6_ASAP7_75t_L g1171 ( .A(n_971), .B(n_1078), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1172 ( .A(n_978), .Y(n_1172) );
BUFx3_ASAP7_75t_L g1173 ( .A(n_985), .Y(n_1173) );
AO21x2_ASAP7_75t_L g1174 ( .A1(n_1064), .A2(n_1065), .B(n_1063), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1068), .B(n_1072), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1089), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1116), .B(n_1126), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1116), .B(n_1126), .Y(n_1178) );
BUFx3_ASAP7_75t_L g1179 ( .A(n_1114), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1139), .B(n_1125), .Y(n_1180) );
INVx1_ASAP7_75t_SL g1181 ( .A(n_1162), .Y(n_1181) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_1171), .Y(n_1182) );
BUFx3_ASAP7_75t_L g1183 ( .A(n_1114), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1113), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1139), .B(n_1133), .Y(n_1185) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1106), .Y(n_1186) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_1093), .B(n_1123), .Y(n_1187) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_1112), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1113), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1111), .B(n_1115), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1111), .Y(n_1191) );
INVxp67_ASAP7_75t_SL g1192 ( .A(n_1134), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1115), .B(n_1119), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1159), .B(n_1104), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1151), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1163), .B(n_1154), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1127), .B(n_1140), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1154), .B(n_1156), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1103), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1103), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1127), .B(n_1136), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1156), .B(n_1160), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1160), .B(n_1097), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1166), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1132), .B(n_1148), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1147), .Y(n_1206) );
INVx5_ASAP7_75t_SL g1207 ( .A(n_1171), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1208 ( .A(n_1112), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1132), .B(n_1148), .Y(n_1209) );
INVx4_ASAP7_75t_L g1210 ( .A(n_1093), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1171), .B(n_1117), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1132), .B(n_1091), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1150), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1091), .B(n_1092), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1092), .B(n_1169), .Y(n_1215) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_1099), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1144), .B(n_1155), .Y(n_1217) );
NAND2x1_ASAP7_75t_L g1218 ( .A(n_1090), .B(n_1100), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1169), .B(n_1175), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1118), .B(n_1120), .Y(n_1220) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_1099), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1096), .B(n_1098), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1121), .B(n_1102), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1155), .B(n_1124), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1105), .B(n_1107), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1108), .B(n_1110), .Y(n_1226) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_1093), .Y(n_1227) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_1123), .Y(n_1228) );
AND2x4_ASAP7_75t_SL g1229 ( .A(n_1172), .B(n_1135), .Y(n_1229) );
BUFx2_ASAP7_75t_L g1230 ( .A(n_1123), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1122), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1141), .B(n_1143), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1143), .B(n_1137), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1167), .B(n_1094), .Y(n_1234) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_1157), .Y(n_1235) );
INVx1_ASAP7_75t_SL g1236 ( .A(n_1188), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1204), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1188), .B(n_1173), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1196), .B(n_1143), .Y(n_1239) );
INVx1_ASAP7_75t_SL g1240 ( .A(n_1208), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1177), .B(n_1138), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1196), .B(n_1094), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1184), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1177), .B(n_1161), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1232), .B(n_1094), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1232), .B(n_1174), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1184), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1195), .B(n_1174), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1233), .B(n_1174), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1233), .B(n_1168), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1189), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1178), .B(n_1109), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1186), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1189), .Y(n_1254) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1218), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1198), .B(n_1130), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1198), .B(n_1130), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1212), .B(n_1205), .Y(n_1258) );
INVx4_ASAP7_75t_L g1259 ( .A(n_1210), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1180), .B(n_1109), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1212), .B(n_1130), .Y(n_1261) );
INVx1_ASAP7_75t_SL g1262 ( .A(n_1229), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1178), .B(n_1109), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1264 ( .A(n_1180), .B(n_1109), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1209), .B(n_1129), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1202), .B(n_1164), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1202), .B(n_1164), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1191), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1190), .B(n_1142), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1193), .B(n_1146), .Y(n_1270) );
INVx3_ASAP7_75t_L g1271 ( .A(n_1218), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1185), .B(n_1131), .Y(n_1272) );
INVx1_ASAP7_75t_SL g1273 ( .A(n_1229), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1176), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1185), .B(n_1170), .Y(n_1275) );
NAND2xp5_ASAP7_75t_SL g1276 ( .A(n_1210), .B(n_1149), .Y(n_1276) );
NOR4xp25_ASAP7_75t_SL g1277 ( .A(n_1227), .B(n_1165), .C(n_1153), .D(n_1152), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1243), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1268), .B(n_1203), .Y(n_1279) );
INVx2_ASAP7_75t_L g1280 ( .A(n_1253), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1258), .B(n_1234), .Y(n_1281) );
NAND2xp33_ASAP7_75t_L g1282 ( .A(n_1262), .B(n_1201), .Y(n_1282) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_1259), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1258), .B(n_1234), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1242), .B(n_1234), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1241), .B(n_1225), .Y(n_1286) );
INVx1_ASAP7_75t_SL g1287 ( .A(n_1236), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1243), .Y(n_1288) );
INVx2_ASAP7_75t_SL g1289 ( .A(n_1259), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1242), .B(n_1234), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1239), .B(n_1223), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1247), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1244), .B(n_1231), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1247), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1246), .B(n_1192), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1237), .Y(n_1296) );
INVxp67_ASAP7_75t_L g1297 ( .A(n_1238), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1237), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1256), .B(n_1199), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1251), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1251), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1257), .B(n_1200), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1254), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1257), .B(n_1200), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1270), .B(n_1231), .Y(n_1305) );
INVx1_ASAP7_75t_SL g1306 ( .A(n_1240), .Y(n_1306) );
NAND2x1p5_ASAP7_75t_L g1307 ( .A(n_1259), .B(n_1187), .Y(n_1307) );
NAND2x1_ASAP7_75t_L g1308 ( .A(n_1255), .B(n_1187), .Y(n_1308) );
INVx1_ASAP7_75t_SL g1309 ( .A(n_1273), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1245), .B(n_1220), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1249), .B(n_1194), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1274), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1272), .B(n_1211), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1278), .Y(n_1314) );
OAI31xp33_ASAP7_75t_L g1315 ( .A1(n_1283), .A2(n_1276), .A3(n_1201), .B(n_1182), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1311), .B(n_1265), .Y(n_1316) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1291), .B(n_1275), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1310), .B(n_1248), .Y(n_1318) );
XNOR2xp5_ASAP7_75t_L g1319 ( .A(n_1287), .B(n_1181), .Y(n_1319) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_1282), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1288), .Y(n_1321) );
CKINVDCx16_ASAP7_75t_R g1322 ( .A(n_1306), .Y(n_1322) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1280), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1292), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1325 ( .A(n_1279), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1299), .B(n_1266), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_1297), .A2(n_1267), .B1(n_1250), .B2(n_1217), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1294), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1302), .B(n_1261), .Y(n_1329) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_1309), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1300), .Y(n_1331) );
OAI21xp33_ASAP7_75t_L g1332 ( .A1(n_1320), .A2(n_1284), .B(n_1281), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1331), .Y(n_1333) );
INVxp67_ASAP7_75t_SL g1334 ( .A(n_1319), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1325), .B(n_1304), .Y(n_1335) );
OAI32xp33_ASAP7_75t_L g1336 ( .A1(n_1322), .A2(n_1307), .A3(n_1289), .B1(n_1295), .B2(n_1286), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1329), .B(n_1281), .Y(n_1337) );
AOI221xp5_ASAP7_75t_SL g1338 ( .A1(n_1330), .A2(n_1305), .B1(n_1290), .B2(n_1285), .C(n_1293), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1323), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1340 ( .A1(n_1338), .A2(n_1327), .B1(n_1316), .B2(n_1315), .C(n_1326), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g1341 ( .A(n_1334), .B(n_1317), .Y(n_1341) );
AOI21xp5_ASAP7_75t_L g1342 ( .A1(n_1336), .A2(n_1308), .B(n_1277), .Y(n_1342) );
AOI221x1_ASAP7_75t_L g1343 ( .A1(n_1332), .A2(n_1328), .B1(n_1324), .B2(n_1314), .C(n_1321), .Y(n_1343) );
OAI211xp5_ASAP7_75t_L g1344 ( .A1(n_1335), .A2(n_1095), .B(n_1217), .C(n_1224), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1333), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1341), .B(n_1337), .Y(n_1346) );
OAI221xp5_ASAP7_75t_SL g1347 ( .A1(n_1340), .A2(n_1313), .B1(n_1318), .B2(n_1263), .C(n_1252), .Y(n_1347) );
OAI221xp5_ASAP7_75t_SL g1348 ( .A1(n_1344), .A2(n_1313), .B1(n_1269), .B2(n_1260), .C(n_1264), .Y(n_1348) );
NAND3xp33_ASAP7_75t_SL g1349 ( .A(n_1342), .B(n_1101), .C(n_1228), .Y(n_1349) );
OAI21xp5_ASAP7_75t_L g1350 ( .A1(n_1343), .A2(n_1222), .B(n_1226), .Y(n_1350) );
AOI211xp5_ASAP7_75t_L g1351 ( .A1(n_1349), .A2(n_1345), .B(n_1271), .C(n_1255), .Y(n_1351) );
NAND3xp33_ASAP7_75t_L g1352 ( .A(n_1347), .B(n_1339), .C(n_1301), .Y(n_1352) );
NOR3xp33_ASAP7_75t_L g1353 ( .A(n_1348), .B(n_1350), .C(n_1346), .Y(n_1353) );
NAND4xp25_ASAP7_75t_L g1354 ( .A(n_1350), .B(n_1271), .C(n_1230), .D(n_1183), .Y(n_1354) );
NOR3xp33_ASAP7_75t_SL g1355 ( .A(n_1354), .B(n_1206), .C(n_1213), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1353), .B(n_1296), .Y(n_1356) );
NAND3xp33_ASAP7_75t_SL g1357 ( .A(n_1351), .B(n_1235), .C(n_1248), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1356), .B(n_1352), .Y(n_1358) );
OR4x2_ASAP7_75t_L g1359 ( .A(n_1357), .B(n_1207), .C(n_1219), .D(n_1214), .Y(n_1359) );
NAND2x1p5_ASAP7_75t_L g1360 ( .A(n_1355), .B(n_1179), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1358), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1362 ( .A(n_1360), .Y(n_1362) );
AOI22xp5_ASAP7_75t_L g1363 ( .A1(n_1362), .A2(n_1359), .B1(n_1221), .B2(n_1216), .Y(n_1363) );
XOR2xp5_ASAP7_75t_L g1364 ( .A(n_1361), .B(n_1197), .Y(n_1364) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_1364), .A2(n_1128), .B1(n_1145), .B2(n_1215), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1363), .Y(n_1366) );
AOI21xp33_ASAP7_75t_L g1367 ( .A1(n_1366), .A2(n_1157), .B(n_1158), .Y(n_1367) );
AOI21xp5_ASAP7_75t_L g1368 ( .A1(n_1367), .A2(n_1365), .B(n_1157), .Y(n_1368) );
AOI221xp5_ASAP7_75t_L g1369 ( .A1(n_1368), .A2(n_1303), .B1(n_1298), .B2(n_1312), .C(n_1235), .Y(n_1369) );
endmodule