module real_aes_4280_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_1392, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_1393, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_1391, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_1392;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_1393;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_1391;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_733;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_483;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_0), .A2(n_276), .B1(n_578), .B2(n_580), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_1), .A2(n_373), .B1(n_616), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_2), .A2(n_352), .B1(n_651), .B2(n_667), .Y(n_875) );
INVx1_ASAP7_75t_L g920 ( .A(n_3), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_4), .A2(n_326), .B1(n_593), .B2(n_594), .Y(n_932) );
INVx1_ASAP7_75t_L g1377 ( .A(n_5), .Y(n_1377) );
INVx1_ASAP7_75t_L g647 ( .A(n_6), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_7), .A2(n_302), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g1383 ( .A1(n_8), .A2(n_340), .B1(n_664), .B2(n_892), .Y(n_1383) );
INVx1_ASAP7_75t_L g824 ( .A(n_9), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_10), .A2(n_226), .B1(n_475), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_11), .A2(n_355), .B1(n_546), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_12), .A2(n_270), .B1(n_529), .B2(n_835), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1209 ( .A(n_13), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_14), .A2(n_172), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_15), .A2(n_254), .B1(n_593), .B2(n_683), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_16), .A2(n_336), .B1(n_643), .B2(n_644), .C(n_646), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g855 ( .A1(n_17), .A2(n_89), .B1(n_574), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g955 ( .A(n_18), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_19), .A2(n_280), .B1(n_626), .B2(n_634), .Y(n_807) );
INVx1_ASAP7_75t_L g923 ( .A(n_20), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_21), .A2(n_23), .B1(n_580), .B2(n_746), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_22), .A2(n_86), .B1(n_664), .B2(n_892), .Y(n_891) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_24), .B(n_450), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_25), .A2(n_162), .B1(n_626), .B2(n_631), .Y(n_1059) );
AOI21xp33_ASAP7_75t_L g1013 ( .A1(n_26), .A2(n_475), .B(n_1014), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_27), .A2(n_284), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g1353 ( .A1(n_28), .A2(n_211), .B1(n_667), .B2(n_835), .Y(n_1353) );
INVx1_ASAP7_75t_L g603 ( .A(n_29), .Y(n_603) );
INVx1_ASAP7_75t_L g918 ( .A(n_30), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_31), .A2(n_403), .B1(n_573), .B2(n_655), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_32), .A2(n_268), .B1(n_785), .B2(n_943), .Y(n_942) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_33), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_34), .A2(n_40), .B1(n_578), .B2(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g906 ( .A(n_35), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_36), .A2(n_260), .B1(n_986), .B2(n_988), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_37), .A2(n_418), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_38), .A2(n_61), .B1(n_848), .B2(n_1068), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_39), .A2(n_106), .B1(n_523), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g799 ( .A(n_41), .Y(n_799) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_42), .A2(n_601), .B(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_43), .A2(n_244), .B1(n_659), .B2(n_775), .Y(n_872) );
INVx1_ASAP7_75t_L g737 ( .A(n_44), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_45), .A2(n_182), .B1(n_542), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_46), .A2(n_145), .B1(n_659), .B2(n_968), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_47), .A2(n_291), .B1(n_692), .B2(n_1012), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_48), .A2(n_347), .B1(n_474), .B2(n_479), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_49), .A2(n_135), .B1(n_628), .B2(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g1376 ( .A(n_50), .Y(n_1376) );
CKINVDCx16_ASAP7_75t_R g718 ( .A(n_51), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_52), .A2(n_222), .B1(n_582), .B2(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_53), .B(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_54), .A2(n_356), .B1(n_576), .B2(n_748), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_55), .A2(n_193), .B1(n_1102), .B2(n_1104), .Y(n_1110) );
INVx1_ASAP7_75t_L g952 ( .A(n_56), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g1354 ( .A1(n_57), .A2(n_300), .B1(n_516), .B2(n_573), .Y(n_1354) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_58), .A2(n_350), .B1(n_470), .B2(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_59), .A2(n_69), .B1(n_578), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_60), .A2(n_271), .B1(n_573), .B2(n_593), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_62), .A2(n_160), .B1(n_628), .B2(n_629), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_63), .A2(n_389), .B1(n_515), .B2(n_523), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_64), .A2(n_289), .B1(n_576), .B2(n_748), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_65), .A2(n_273), .B1(n_685), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_66), .A2(n_411), .B1(n_608), .B2(n_661), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_67), .A2(n_421), .B1(n_662), .B2(n_777), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_68), .A2(n_405), .B1(n_619), .B2(n_925), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_70), .A2(n_390), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g489 ( .A1(n_71), .A2(n_490), .B(n_494), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_72), .B(n_717), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_73), .A2(n_170), .B1(n_982), .B2(n_1074), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_74), .A2(n_415), .B1(n_539), .B2(n_582), .Y(n_1024) );
OA22x2_ASAP7_75t_L g448 ( .A1(n_75), .A2(n_192), .B1(n_449), .B2(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g486 ( .A(n_75), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_76), .A2(n_168), .B1(n_628), .B2(n_629), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_77), .A2(n_228), .B1(n_565), .B2(n_614), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_78), .A2(n_369), .B1(n_633), .B2(n_634), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_79), .A2(n_133), .B1(n_565), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g1124 ( .A(n_80), .Y(n_1124) );
NAND2xp33_ASAP7_75t_L g708 ( .A(n_81), .B(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_82), .A2(n_179), .B1(n_1115), .B2(n_1123), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_83), .A2(n_181), .B1(n_605), .B2(n_850), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_84), .A2(n_263), .B1(n_546), .B2(n_576), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_85), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g1126 ( .A(n_87), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_88), .B(n_214), .Y(n_432) );
INVx1_ASAP7_75t_L g456 ( .A(n_88), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g487 ( .A1(n_88), .A2(n_192), .B(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_90), .A2(n_131), .B1(n_1095), .B2(n_1099), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_91), .A2(n_304), .B1(n_524), .B2(n_574), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_92), .A2(n_148), .B1(n_690), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_93), .A2(n_299), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_94), .A2(n_313), .B1(n_539), .B2(n_582), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_95), .A2(n_262), .B1(n_539), .B2(n_542), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_96), .A2(n_215), .B1(n_643), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_97), .A2(n_398), .B1(n_516), .B2(n_834), .Y(n_992) );
INVx1_ASAP7_75t_L g827 ( .A(n_98), .Y(n_827) );
INVx1_ASAP7_75t_L g1343 ( .A(n_99), .Y(n_1343) );
AOI22xp33_ASAP7_75t_SL g1363 ( .A1(n_100), .A2(n_1364), .B1(n_1385), .B2(n_1386), .Y(n_1363) );
INVx1_ASAP7_75t_L g1385 ( .A(n_100), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_101), .A2(n_266), .B1(n_516), .B2(n_667), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_102), .A2(n_123), .B1(n_664), .B2(n_892), .Y(n_994) );
AOI21xp33_ASAP7_75t_L g1031 ( .A1(n_103), .A2(n_643), .B(n_1032), .Y(n_1031) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_104), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1097 ( .A(n_105), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_105), .B(n_325), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_107), .A2(n_269), .B1(n_654), .B2(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g961 ( .A(n_108), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_109), .A2(n_371), .B1(n_1095), .B2(n_1112), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_110), .A2(n_341), .B1(n_539), .B2(n_582), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_111), .A2(n_174), .B1(n_516), .B2(n_546), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_112), .A2(n_188), .B1(n_560), .B2(n_605), .Y(n_750) );
INVx1_ASAP7_75t_L g831 ( .A(n_113), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_114), .A2(n_202), .B1(n_654), .B2(n_835), .Y(n_995) );
AO22x1_ASAP7_75t_L g1022 ( .A1(n_115), .A2(n_366), .B1(n_574), .B2(n_856), .Y(n_1022) );
AO22x2_ASAP7_75t_L g1140 ( .A1(n_116), .A2(n_346), .B1(n_1095), .B2(n_1112), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_117), .A2(n_213), .B1(n_717), .B2(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_118), .A2(n_142), .B1(n_788), .B2(n_791), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_119), .A2(n_177), .B1(n_605), .B2(n_690), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_120), .A2(n_322), .B1(n_529), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_121), .A2(n_139), .B1(n_470), .B2(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_122), .A2(n_267), .B1(n_565), .B2(n_605), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_124), .A2(n_169), .B1(n_578), .B2(n_668), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_125), .A2(n_156), .B1(n_1123), .B2(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_126), .A2(n_348), .B1(n_654), .B2(n_1083), .Y(n_1384) );
INVx1_ASAP7_75t_L g739 ( .A(n_127), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_127), .A2(n_159), .B1(n_1102), .B2(n_1104), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_128), .A2(n_134), .B1(n_573), .B2(n_655), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_129), .A2(n_150), .B1(n_651), .B2(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_130), .A2(n_380), .B1(n_856), .B2(n_1057), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_132), .B(n_428), .Y(n_1098) );
INVx1_ASAP7_75t_SL g1103 ( .A(n_132), .Y(n_1103) );
INVx1_ASAP7_75t_L g1106 ( .A(n_132), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_136), .A2(n_401), .B1(n_651), .B2(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g1034 ( .A(n_137), .B(n_491), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g977 ( .A1(n_138), .A2(n_978), .B(n_979), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_140), .B(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_141), .A2(n_240), .B1(n_668), .B2(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g1336 ( .A(n_143), .Y(n_1336) );
AO22x2_ASAP7_75t_L g945 ( .A1(n_144), .A2(n_183), .B1(n_701), .B2(n_946), .Y(n_945) );
XOR2x2_ASAP7_75t_L g936 ( .A(n_146), .B(n_937), .Y(n_936) );
AOI33xp33_ASAP7_75t_R g859 ( .A1(n_147), .A2(n_298), .A3(n_472), .B1(n_482), .B2(n_860), .B3(n_1393), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_149), .A2(n_166), .B1(n_1095), .B2(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g999 ( .A(n_151), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_151), .A2(n_419), .B1(n_1095), .B2(n_1115), .Y(n_1136) );
INVx1_ASAP7_75t_L g1064 ( .A(n_152), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_153), .A2(n_319), .B1(n_617), .B2(n_625), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_154), .A2(n_317), .B1(n_664), .B2(n_665), .Y(n_1080) );
AO22x1_ASAP7_75t_L g653 ( .A1(n_155), .A2(n_368), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_157), .A2(n_199), .B1(n_787), .B2(n_789), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_158), .A2(n_286), .B1(n_444), .B2(n_468), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_161), .A2(n_379), .B1(n_643), .B2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_163), .A2(n_399), .B1(n_690), .B2(n_982), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_164), .A2(n_197), .B1(n_546), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_165), .A2(n_312), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_167), .A2(n_232), .B1(n_562), .B2(n_608), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_171), .A2(n_351), .B1(n_600), .B2(n_601), .C(n_602), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_173), .A2(n_394), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_175), .A2(n_178), .B1(n_573), .B2(n_655), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_176), .A2(n_339), .B1(n_445), .B2(n_848), .Y(n_847) );
AOI22x1_ASAP7_75t_L g973 ( .A1(n_179), .A2(n_974), .B1(n_975), .B2(n_996), .Y(n_973) );
INVx1_ASAP7_75t_L g996 ( .A(n_179), .Y(n_996) );
INVx1_ASAP7_75t_L g980 ( .A(n_180), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_184), .B(n_491), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_185), .A2(n_272), .B1(n_608), .B2(n_871), .Y(n_870) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_186), .A2(n_354), .B1(n_539), .B2(n_582), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_187), .A2(n_408), .B1(n_651), .B2(n_667), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_189), .A2(n_205), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_190), .A2(n_382), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g467 ( .A(n_191), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_191), .B(n_258), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_191), .B(n_484), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_192), .B(n_335), .Y(n_431) );
XNOR2x1_ASAP7_75t_L g722 ( .A(n_193), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g679 ( .A(n_194), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_195), .A2(n_223), .B1(n_692), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_SL g1350 ( .A1(n_196), .A2(n_229), .B1(n_654), .B2(n_1077), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_198), .A2(n_386), .B1(n_573), .B2(n_655), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_200), .B(n_601), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_201), .A2(n_209), .B1(n_546), .B2(n_591), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_203), .A2(n_221), .B1(n_631), .B2(n_633), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_204), .A2(n_308), .B1(n_654), .B2(n_655), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_206), .A2(n_331), .B1(n_580), .B2(n_746), .Y(n_1025) );
CKINVDCx5p33_ASAP7_75t_R g1129 ( .A(n_207), .Y(n_1129) );
INVx1_ASAP7_75t_L g822 ( .A(n_208), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_210), .A2(n_230), .B1(n_622), .B2(n_659), .Y(n_820) );
INVx1_ASAP7_75t_L g1371 ( .A(n_212), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_214), .B(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_216), .A2(n_248), .B1(n_516), .B2(n_573), .Y(n_838) );
INVx1_ASAP7_75t_L g1374 ( .A(n_217), .Y(n_1374) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_218), .A2(n_392), .B1(n_654), .B2(n_835), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_219), .A2(n_296), .B1(n_787), .B2(n_892), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_220), .A2(n_374), .B1(n_829), .B2(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g715 ( .A(n_224), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_225), .A2(n_416), .B1(n_538), .B2(n_541), .Y(n_537) );
INVxp33_ASAP7_75t_SL g1131 ( .A(n_227), .Y(n_1131) );
XNOR2x1_ASAP7_75t_L g1332 ( .A(n_227), .B(n_1333), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_227), .A2(n_1360), .B1(n_1362), .B2(n_1387), .Y(n_1359) );
INVx1_ASAP7_75t_L g696 ( .A(n_231), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_233), .A2(n_278), .B1(n_539), .B2(n_582), .Y(n_742) );
INVx1_ASAP7_75t_L g1341 ( .A(n_234), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_235), .B(n_661), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_236), .A2(n_409), .B1(n_626), .B2(n_631), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_237), .A2(n_383), .B1(n_560), .B2(n_605), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_238), .A2(n_420), .B1(n_605), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_239), .A2(n_406), .B1(n_1112), .B2(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g963 ( .A(n_241), .Y(n_963) );
INVx1_ASAP7_75t_L g1346 ( .A(n_242), .Y(n_1346) );
INVx1_ASAP7_75t_L g913 ( .A(n_243), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_245), .A2(n_282), .B1(n_591), .B2(n_625), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_246), .A2(n_365), .B1(n_746), .B2(n_941), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_247), .A2(n_412), .B1(n_601), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g1051 ( .A(n_249), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_250), .A2(n_367), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_251), .A2(n_293), .B1(n_545), .B2(n_548), .Y(n_544) );
XOR2x2_ASAP7_75t_L g844 ( .A(n_252), .B(n_845), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_253), .A2(n_349), .B1(n_665), .B2(n_787), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_255), .A2(n_330), .B1(n_600), .B2(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_256), .B(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_257), .A2(n_404), .B1(n_628), .B2(n_629), .Y(n_810) );
INVx1_ASAP7_75t_L g454 ( .A(n_258), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_259), .B(n_865), .Y(n_1072) );
INVx1_ASAP7_75t_L g640 ( .A(n_261), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_261), .A2(n_657), .B1(n_663), .B2(n_666), .C1(n_1391), .C2(n_1392), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_261), .B(n_666), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_264), .A2(n_402), .B1(n_617), .B2(n_625), .Y(n_808) );
INVx1_ASAP7_75t_L g586 ( .A(n_265), .Y(n_586) );
XNOR2x1_ASAP7_75t_L g440 ( .A(n_274), .B(n_441), .Y(n_440) );
XNOR2x2_ASAP7_75t_SL g635 ( .A(n_274), .B(n_441), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_275), .A2(n_314), .B1(n_664), .B2(n_665), .Y(n_876) );
INVx1_ASAP7_75t_L g903 ( .A(n_277), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_279), .A2(n_295), .B1(n_605), .B2(n_606), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_281), .A2(n_327), .B1(n_534), .B2(n_573), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_283), .A2(n_643), .B(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g752 ( .A1(n_285), .A2(n_305), .B1(n_643), .B2(n_753), .C(n_754), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_287), .A2(n_768), .B(n_771), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_288), .A2(n_385), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_290), .A2(n_407), .B1(n_601), .B2(n_620), .Y(n_734) );
OAI21x1_ASAP7_75t_L g1017 ( .A1(n_292), .A2(n_1018), .B(n_1035), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_292), .B(n_1021), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_292), .A2(n_400), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_294), .A2(n_387), .B1(n_600), .B2(n_733), .C(n_1050), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_297), .A2(n_310), .B1(n_848), .B2(n_1053), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_301), .A2(n_370), .B1(n_516), .B2(n_667), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_303), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g772 ( .A(n_306), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_307), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g1015 ( .A(n_309), .Y(n_1015) );
INVx1_ASAP7_75t_L g504 ( .A(n_311), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_315), .A2(n_345), .B1(n_546), .B2(n_576), .Y(n_928) );
INVx1_ASAP7_75t_L g1367 ( .A(n_316), .Y(n_1367) );
INVx1_ASAP7_75t_L g960 ( .A(n_318), .Y(n_960) );
INVx1_ASAP7_75t_L g815 ( .A(n_320), .Y(n_815) );
INVx1_ASAP7_75t_L g755 ( .A(n_321), .Y(n_755) );
AO22x1_ASAP7_75t_L g1141 ( .A1(n_323), .A2(n_329), .B1(n_1102), .B2(n_1116), .Y(n_1141) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_324), .A2(n_900), .B(n_902), .Y(n_899) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_325), .Y(n_433) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_325), .B(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_328), .A2(n_333), .B1(n_633), .B2(n_634), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g1046 ( .A(n_329), .B(n_1047), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_332), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g948 ( .A(n_334), .Y(n_948) );
INVx1_ASAP7_75t_L g465 ( .A(n_335), .Y(n_465) );
INVxp67_ASAP7_75t_L g503 ( .A(n_335), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_337), .A2(n_410), .B1(n_528), .B2(n_533), .Y(n_527) );
INVx1_ASAP7_75t_L g1033 ( .A(n_338), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_342), .A2(n_378), .B1(n_664), .B2(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g428 ( .A(n_343), .Y(n_428) );
INVxp33_ASAP7_75t_SL g1210 ( .A(n_344), .Y(n_1210) );
INVx1_ASAP7_75t_L g915 ( .A(n_353), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_357), .A2(n_361), .B1(n_616), .B2(n_620), .Y(n_803) );
XNOR2x2_ASAP7_75t_L g861 ( .A(n_358), .B(n_862), .Y(n_861) );
AO221x2_ASAP7_75t_L g1206 ( .A1(n_359), .A2(n_360), .B1(n_1163), .B2(n_1207), .C(n_1208), .Y(n_1206) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_362), .A2(n_600), .B(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_363), .A2(n_381), .B1(n_445), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_364), .A2(n_376), .B1(n_600), .B2(n_619), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_372), .B(n_661), .Y(n_853) );
INVx1_ASAP7_75t_L g957 ( .A(n_375), .Y(n_957) );
XOR2xp5_ASAP7_75t_L g610 ( .A(n_377), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g1337 ( .A(n_384), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_388), .A2(n_393), .B1(n_565), .B2(n_614), .Y(n_1028) );
INVx1_ASAP7_75t_L g583 ( .A(n_391), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_395), .A2(n_414), .B1(n_717), .B2(n_733), .Y(n_804) );
AO22x2_ASAP7_75t_L g907 ( .A1(n_396), .A2(n_908), .B1(n_909), .B2(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_396), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_397), .A2(n_413), .B1(n_834), .B2(n_835), .Y(n_833) );
XOR2x2_ASAP7_75t_L g764 ( .A(n_417), .B(n_765), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_434), .B(n_1086), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx4_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .C(n_433), .Y(n_425) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_426), .B(n_1357), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_426), .B(n_1358), .Y(n_1361) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OA21x2_ASAP7_75t_L g1388 ( .A1(n_427), .A2(n_1103), .B(n_1389), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND3x4_ASAP7_75t_L g1102 ( .A(n_428), .B(n_1096), .C(n_1103), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_428), .B(n_1106), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_429), .B(n_1358), .Y(n_1357) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_430), .A2(n_510), .B(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g1358 ( .A(n_433), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_883), .B1(n_1084), .B2(n_1085), .Y(n_434) );
INVx1_ASAP7_75t_L g1084 ( .A(n_435), .Y(n_1084) );
XNOR2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_761), .Y(n_435) );
XNOR2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_636), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_552), .B1(n_553), .B2(n_635), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_513), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_473), .C(n_489), .Y(n_442) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g914 ( .A(n_445), .Y(n_914) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_446), .Y(n_643) );
BUFx3_ASAP7_75t_L g692 ( .A(n_446), .Y(n_692) );
INVx1_ASAP7_75t_L g830 ( .A(n_446), .Y(n_830) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_457), .Y(n_446) );
AND2x4_ASAP7_75t_L g476 ( .A(n_447), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g600 ( .A(n_447), .B(n_457), .Y(n_600) );
AND2x2_ASAP7_75t_L g733 ( .A(n_447), .B(n_477), .Y(n_733) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
AND2x2_ASAP7_75t_L g472 ( .A(n_448), .B(n_452), .Y(n_472) );
AND2x2_ASAP7_75t_L g501 ( .A(n_448), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g519 ( .A(n_448), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_449), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp33_ASAP7_75t_L g453 ( .A(n_450), .B(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g460 ( .A(n_450), .Y(n_460) );
NAND2xp33_ASAP7_75t_L g466 ( .A(n_450), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g488 ( .A(n_450), .Y(n_488) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_450), .Y(n_499) );
AND2x4_ASAP7_75t_L g518 ( .A(n_451), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_454), .B(n_486), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_456), .A2(n_488), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g471 ( .A(n_457), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g540 ( .A(n_457), .B(n_518), .Y(n_540) );
AND2x4_ASAP7_75t_L g616 ( .A(n_457), .B(n_472), .Y(n_616) );
AND2x4_ASAP7_75t_L g628 ( .A(n_457), .B(n_518), .Y(n_628) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
INVx2_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
AND2x2_ASAP7_75t_L g497 ( .A(n_458), .B(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g521 ( .A(n_458), .B(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g531 ( .A(n_458), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_460), .B(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g484 ( .A(n_460), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_461), .B(n_483), .C(n_512), .Y(n_511) );
AND2x4_ASAP7_75t_L g477 ( .A(n_462), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g522 ( .A(n_463), .Y(n_522) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_469), .A2(n_827), .B1(n_828), .B2(n_831), .Y(n_826) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g780 ( .A(n_470), .Y(n_780) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_471), .Y(n_605) );
INVx2_ASAP7_75t_L g869 ( .A(n_471), .Y(n_869) );
AND2x2_ASAP7_75t_L g493 ( .A(n_472), .B(n_477), .Y(n_493) );
AND2x2_ASAP7_75t_L g530 ( .A(n_472), .B(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g535 ( .A(n_472), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g579 ( .A(n_472), .B(n_531), .Y(n_579) );
AND2x2_ASAP7_75t_L g601 ( .A(n_472), .B(n_477), .Y(n_601) );
AND2x4_ASAP7_75t_L g626 ( .A(n_472), .B(n_520), .Y(n_626) );
AND2x4_ASAP7_75t_L g631 ( .A(n_472), .B(n_531), .Y(n_631) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g563 ( .A(n_476), .Y(n_563) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_476), .Y(n_614) );
BUFx3_ASAP7_75t_L g661 ( .A(n_476), .Y(n_661) );
BUFx8_ASAP7_75t_SL g871 ( .A(n_476), .Y(n_871) );
INVx2_ASAP7_75t_L g1069 ( .A(n_476), .Y(n_1069) );
AND2x4_ASAP7_75t_L g481 ( .A(n_477), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_518), .Y(n_543) );
AND2x4_ASAP7_75t_L g620 ( .A(n_477), .B(n_482), .Y(n_620) );
AND2x4_ASAP7_75t_L g629 ( .A(n_477), .B(n_518), .Y(n_629) );
INVx1_ASAP7_75t_L g1344 ( .A(n_479), .Y(n_1344) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g608 ( .A(n_480), .Y(n_608) );
INVx2_ASAP7_75t_L g848 ( .A(n_480), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_480), .A2(n_919), .B1(n_960), .B2(n_961), .Y(n_959) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_481), .Y(n_565) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_481), .Y(n_662) );
AND2x4_ASAP7_75t_L g526 ( .A(n_482), .B(n_520), .Y(n_526) );
AND2x4_ASAP7_75t_L g551 ( .A(n_482), .B(n_531), .Y(n_551) );
AND2x4_ASAP7_75t_L g633 ( .A(n_482), .B(n_531), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_482), .B(n_520), .Y(n_634) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_SL g709 ( .A(n_492), .Y(n_709) );
INVx2_ASAP7_75t_L g753 ( .A(n_492), .Y(n_753) );
INVx2_ASAP7_75t_L g770 ( .A(n_492), .Y(n_770) );
INVx2_ASAP7_75t_L g1053 ( .A(n_492), .Y(n_1053) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx3_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
INVx2_ASAP7_75t_L g819 ( .A(n_493), .Y(n_819) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_504), .B(n_505), .Y(n_494) );
INVx2_ASAP7_75t_L g606 ( .A(n_495), .Y(n_606) );
INVx2_ASAP7_75t_L g659 ( .A(n_495), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g902 ( .A1(n_495), .A2(n_903), .B(n_904), .Y(n_902) );
OAI21xp33_ASAP7_75t_L g979 ( .A1(n_495), .A2(n_980), .B(n_981), .Y(n_979) );
INVx4_ASAP7_75t_L g1012 ( .A(n_495), .Y(n_1012) );
INVx2_ASAP7_75t_L g1074 ( .A(n_495), .Y(n_1074) );
INVx5_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
BUFx4f_ASAP7_75t_L g690 ( .A(n_496), .Y(n_690) );
BUFx2_ASAP7_75t_L g850 ( .A(n_496), .Y(n_850) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
AND2x2_ASAP7_75t_L g619 ( .A(n_497), .B(n_501), .Y(n_619) );
AND2x4_ASAP7_75t_L g731 ( .A(n_497), .B(n_501), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g510 ( .A(n_499), .Y(n_510) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_507), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g775 ( .A(n_507), .Y(n_775) );
INVx4_ASAP7_75t_L g968 ( .A(n_507), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_507), .B(n_1015), .Y(n_1014) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g983 ( .A(n_508), .Y(n_983) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_509), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_527), .C(n_537), .D(n_544), .Y(n_513) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_517), .Y(n_651) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g547 ( .A(n_518), .B(n_531), .Y(n_547) );
AND2x4_ASAP7_75t_L g617 ( .A(n_518), .B(n_536), .Y(n_617) );
AND2x4_ASAP7_75t_L g625 ( .A(n_518), .B(n_531), .Y(n_625) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g536 ( .A(n_521), .Y(n_536) );
INVx1_ASAP7_75t_L g532 ( .A(n_522), .Y(n_532) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g594 ( .A(n_525), .Y(n_594) );
INVx1_ASAP7_75t_L g652 ( .A(n_525), .Y(n_652) );
INVx2_ASAP7_75t_L g683 ( .A(n_525), .Y(n_683) );
INVx5_ASAP7_75t_L g856 ( .A(n_525), .Y(n_856) );
INVx1_ASAP7_75t_L g1078 ( .A(n_525), .Y(n_1078) );
INVx6_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx12f_ASAP7_75t_L g573 ( .A(n_526), .Y(n_573) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_529), .Y(n_1082) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx8_ASAP7_75t_L g654 ( .A(n_530), .Y(n_654) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_531), .Y(n_860) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx12f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_535), .Y(n_574) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_535), .Y(n_593) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_535), .Y(n_655) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_535), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx12f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g597 ( .A(n_540), .Y(n_597) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_540), .Y(n_664) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_543), .Y(n_582) );
BUFx5_ASAP7_75t_L g665 ( .A(n_543), .Y(n_665) );
INVx1_ASAP7_75t_L g792 ( .A(n_543), .Y(n_792) );
INVx1_ASAP7_75t_L g949 ( .A(n_545), .Y(n_949) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g795 ( .A(n_546), .Y(n_795) );
BUFx12f_ASAP7_75t_L g834 ( .A(n_546), .Y(n_834) );
BUFx12f_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_547), .Y(n_667) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_547), .Y(n_748) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
INVx4_ASAP7_75t_L g668 ( .A(n_550), .Y(n_668) );
INVx2_ASAP7_75t_SL g685 ( .A(n_550), .Y(n_685) );
INVx2_ASAP7_75t_L g706 ( .A(n_550), .Y(n_706) );
INVx4_ASAP7_75t_L g835 ( .A(n_550), .Y(n_835) );
INVx1_ASAP7_75t_L g1083 ( .A(n_550), .Y(n_1083) );
INVx8_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
XNOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_584), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g843 ( .A(n_556), .B(n_844), .Y(n_843) );
XOR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_583), .Y(n_556) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .C(n_564), .D(n_566), .Y(n_558) );
INVx2_ASAP7_75t_L g1342 ( .A(n_562), .Y(n_1342) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g777 ( .A(n_563), .Y(n_777) );
INVx3_ASAP7_75t_L g921 ( .A(n_565), .Y(n_921) );
INVx2_ASAP7_75t_L g645 ( .A(n_567), .Y(n_645) );
INVx1_ASAP7_75t_L g966 ( .A(n_567), .Y(n_966) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_569), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_569), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g1032 ( .A(n_569), .B(n_1033), .Y(n_1032) );
NOR2xp67_ASAP7_75t_SL g1050 ( .A(n_569), .B(n_1051), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g622 ( .A(n_570), .Y(n_622) );
INVx2_ASAP7_75t_L g717 ( .A(n_570), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_570), .B(n_737), .Y(n_736) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_570), .Y(n_756) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .C(n_577), .D(n_581), .Y(n_571) );
BUFx3_ASAP7_75t_L g943 ( .A(n_573), .Y(n_943) );
BUFx3_ASAP7_75t_L g785 ( .A(n_574), .Y(n_785) );
BUFx3_ASAP7_75t_L g783 ( .A(n_576), .Y(n_783) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_579), .Y(n_746) );
BUFx2_ASAP7_75t_L g941 ( .A(n_580), .Y(n_941) );
BUFx2_ASAP7_75t_SL g946 ( .A(n_582), .Y(n_946) );
XNOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_609), .Y(n_584) );
XNOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_598), .Y(n_587) );
NAND4xp25_ASAP7_75t_SL g588 ( .A(n_589), .B(n_590), .C(n_592), .D(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g701 ( .A(n_597), .Y(n_701) );
INVx2_ASAP7_75t_L g788 ( .A(n_597), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_604), .C(n_607), .Y(n_598) );
INVx3_ASAP7_75t_L g916 ( .A(n_605), .Y(n_916) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_623), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .C(n_618), .D(n_621), .Y(n_612) );
INVx2_ASAP7_75t_L g919 ( .A(n_614), .Y(n_919) );
BUFx3_ASAP7_75t_L g1373 ( .A(n_614), .Y(n_1373) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .C(n_630), .D(n_632), .Y(n_623) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_633), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_719), .B1(n_758), .B2(n_759), .Y(n_636) );
INVx1_ASAP7_75t_L g758 ( .A(n_637), .Y(n_758) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_676), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_639), .B(n_669), .Y(n_638) );
AOI21x1_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B(n_656), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_648), .Y(n_641) );
BUFx2_ASAP7_75t_L g670 ( .A(n_642), .Y(n_670) );
INVx4_ASAP7_75t_L g956 ( .A(n_643), .Y(n_956) );
INVx1_ASAP7_75t_L g1368 ( .A(n_644), .Y(n_1368) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g922 ( .A1(n_645), .A2(n_923), .B(n_924), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g674 ( .A(n_650), .B(n_663), .Y(n_674) );
BUFx3_ASAP7_75t_L g951 ( .A(n_651), .Y(n_951) );
INVx1_ASAP7_75t_L g675 ( .A(n_653), .Y(n_675) );
INVx1_ASAP7_75t_L g673 ( .A(n_657), .Y(n_673) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx2_ASAP7_75t_L g823 ( .A(n_661), .Y(n_823) );
BUFx3_ASAP7_75t_L g778 ( .A(n_662), .Y(n_778) );
INVx4_ASAP7_75t_L g825 ( .A(n_662), .Y(n_825) );
NAND4xp75_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .C(n_674), .D(n_675), .Y(n_669) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
XOR2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_697), .Y(n_676) );
XNOR2x1_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_688), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .C(n_686), .D(n_687), .Y(n_681) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .C(n_693), .D(n_694), .Y(n_688) );
INVx2_ASAP7_75t_SL g773 ( .A(n_690), .Y(n_773) );
INVx2_ASAP7_75t_L g987 ( .A(n_692), .Y(n_987) );
XNOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_718), .Y(n_697) );
NAND4xp75_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .C(n_707), .D(n_711), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g760 ( .A(n_720), .Y(n_760) );
AO22x2_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_738), .B2(n_757), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
XNOR2xp5_ASAP7_75t_L g1045 ( .A(n_722), .B(n_1046), .Y(n_1045) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .C(n_727), .D(n_728), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .C(n_734), .D(n_735), .Y(n_729) );
INVx1_ASAP7_75t_L g757 ( .A(n_738), .Y(n_757) );
XNOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .C(n_749), .D(n_752), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g901 ( .A(n_753), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g925 ( .A(n_756), .Y(n_925) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_840), .B1(n_880), .B2(n_881), .Y(n_761) );
INVx2_ASAP7_75t_SL g880 ( .A(n_762), .Y(n_880) );
AO22x2_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_796), .B2(n_839), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_781), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_776), .C(n_779), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g1345 ( .A1(n_769), .A2(n_1346), .B(n_1347), .Y(n_1345) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_774), .Y(n_771) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .C(n_786), .D(n_793), .Y(n_781) );
BUFx4f_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
BUFx6f_ASAP7_75t_L g892 ( .A(n_791), .Y(n_892) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g839 ( .A(n_796), .Y(n_839) );
XNOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_811), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
XNOR2x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
OR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_806), .Y(n_800) );
NAND4xp25_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .C(n_804), .D(n_805), .Y(n_801) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .C(n_809), .D(n_810), .Y(n_806) );
NAND2x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_832), .Y(n_812) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_821), .C(n_826), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_820), .Y(n_814) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g865 ( .A(n_818), .Y(n_865) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g852 ( .A(n_819), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g1370 ( .A1(n_825), .A2(n_1371), .B1(n_1372), .B2(n_1374), .Y(n_1370) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AND4x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_836), .C(n_837), .D(n_838), .Y(n_832) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_861), .B(n_878), .Y(n_841) );
OA21x2_ASAP7_75t_L g882 ( .A1(n_842), .A2(n_861), .B(n_878), .Y(n_882) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g879 ( .A(n_843), .Y(n_879) );
NOR2x1_ASAP7_75t_L g845 ( .A(n_846), .B(n_854), .Y(n_845) );
NAND4xp25_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .C(n_851), .D(n_853), .Y(n_846) );
BUFx3_ASAP7_75t_L g978 ( .A(n_852), .Y(n_978) );
NAND4xp25_ASAP7_75t_L g854 ( .A(n_855), .B(n_857), .C(n_858), .D(n_859), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_861), .B(n_879), .Y(n_878) );
OR2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_873), .Y(n_862) );
NAND4xp25_ASAP7_75t_L g863 ( .A(n_864), .B(n_866), .C(n_870), .D(n_872), .Y(n_863) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g898 ( .A(n_868), .Y(n_898) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_868), .Y(n_958) );
INVx2_ASAP7_75t_L g1071 ( .A(n_868), .Y(n_1071) );
INVx1_ASAP7_75t_L g1379 ( .A(n_868), .Y(n_1379) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g990 ( .A(n_869), .Y(n_990) );
INVx1_ASAP7_75t_L g1339 ( .A(n_869), .Y(n_1339) );
NAND4xp25_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .C(n_876), .D(n_877), .Y(n_873) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g1085 ( .A(n_883), .Y(n_1085) );
XNOR2x2_ASAP7_75t_L g883 ( .A(n_884), .B(n_970), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_935), .B1(n_936), .B2(n_969), .Y(n_886) );
INVx1_ASAP7_75t_L g969 ( .A(n_887), .Y(n_969) );
AO22x2_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_907), .B1(n_933), .B2(n_934), .Y(n_887) );
INVx1_ASAP7_75t_L g933 ( .A(n_888), .Y(n_933) );
XOR2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_906), .Y(n_888) );
NOR2x1_ASAP7_75t_L g889 ( .A(n_890), .B(n_896), .Y(n_889) );
NAND4xp25_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .C(n_894), .D(n_895), .Y(n_890) );
NAND3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .C(n_905), .Y(n_896) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx2_ASAP7_75t_L g934 ( .A(n_907), .Y(n_934) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_926), .Y(n_910) );
NOR3xp33_ASAP7_75t_SL g911 ( .A(n_912), .B(n_917), .C(n_922), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_944), .C(n_953), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_942), .Y(n_939) );
NOR2x1_ASAP7_75t_L g944 ( .A(n_945), .B(n_947), .Y(n_944) );
OAI22x1_ASAP7_75t_SL g947 ( .A1(n_948), .A2(n_949), .B1(n_950), .B2(n_952), .Y(n_947) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
NOR3xp33_ASAP7_75t_SL g953 ( .A(n_954), .B(n_959), .C(n_962), .Y(n_953) );
OAI22xp5_ASAP7_75t_SL g954 ( .A1(n_955), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_956), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1375) );
OAI21xp33_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_964), .B(n_967), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
XNOR2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_1040), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
XNOR2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_997), .Y(n_972) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_976), .B(n_991), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_977), .B(n_984), .C(n_985), .Y(n_976) );
INVx4_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g1335 ( .A1(n_987), .A2(n_1336), .B1(n_1337), .B2(n_1338), .Y(n_1335) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
NAND4xp25_ASAP7_75t_SL g991 ( .A(n_992), .B(n_993), .C(n_994), .D(n_995), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1016), .B1(n_1017), .B2(n_1039), .Y(n_997) );
INVx1_ASAP7_75t_L g1039 ( .A(n_998), .Y(n_1039) );
XNOR2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1000), .Y(n_998) );
NOR4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1004), .C(n_1007), .D(n_1010), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
NAND2xp5_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1013), .Y(n_1010) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1017), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1026), .Y(n_1018) );
NOR3xp33_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1022), .C(n_1023), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NOR3xp33_ASAP7_75t_L g1037 ( .A(n_1022), .B(n_1030), .C(n_1038), .Y(n_1037) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_1023), .B(n_1027), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1030), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1034), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B1(n_1062), .B2(n_1063), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
OA22x2_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1044), .B1(n_1045), .B2(n_1061), .Y(n_1042) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1043), .Y(n_1061) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NOR2x1_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1055), .Y(n_1047) );
NAND3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1052), .C(n_1054), .Y(n_1048) );
NAND4xp25_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1058), .C(n_1059), .D(n_1060), .Y(n_1055) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
XNOR2x1_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1075), .Y(n_1065) );
NAND4xp25_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1070), .C(n_1072), .D(n_1073), .Y(n_1066) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_1069), .Y(n_1068) );
NAND4xp25_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1079), .C(n_1080), .D(n_1081), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1330), .B1(n_1331), .B2(n_1355), .C(n_1359), .Y(n_1086) );
O2A1O1Ixp33_ASAP7_75t_SL g1087 ( .A1(n_1088), .A2(n_1211), .B(n_1235), .C(n_1301), .Y(n_1087) );
NAND5xp2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1177), .C(n_1192), .D(n_1201), .E(n_1206), .Y(n_1088) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1137), .B1(n_1142), .B2(n_1150), .C(n_1153), .Y(n_1089) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1107), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1092), .B(n_1240), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1092), .B(n_1255), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1093), .B(n_1120), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1093), .B(n_1139), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_1093), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_1093), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1093), .B(n_1181), .Y(n_1205) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_1093), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1093), .B(n_1120), .Y(n_1222) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1093), .B(n_1227), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1093), .B(n_1139), .Y(n_1273) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1101), .Y(n_1093) );
AND2x4_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1098), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_1096), .B(n_1105), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1096), .B(n_1098), .Y(n_1130) );
AND2x4_ASAP7_75t_L g1165 ( .A(n_1096), .B(n_1098), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_1096), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1098), .B(n_1100), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_1098), .B(n_1100), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1098), .B(n_1100), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1100), .B(n_1105), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1100), .B(n_1105), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_1100), .B(n_1105), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1118), .Y(n_1107) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1108), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1108), .B(n_1147), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1108), .B(n_1144), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1108), .B(n_1132), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1113), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_1109), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1109), .B(n_1113), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1112), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1113), .B(n_1149), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1113), .B(n_1149), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1113), .B(n_1144), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1113), .B(n_1203), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1113), .B(n_1133), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1117), .Y(n_1113) );
INVx3_ASAP7_75t_L g1128 ( .A(n_1115), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1118), .B(n_1169), .Y(n_1176) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1119), .B(n_1148), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1132), .Y(n_1119) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1120), .Y(n_1147) );
INVx3_ASAP7_75t_L g1181 ( .A(n_1120), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1120), .B(n_1186), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1120), .B(n_1148), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1120), .B(n_1273), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_1120), .Y(n_1277) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1120), .B(n_1139), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1127), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_1122), .A2(n_1125), .B1(n_1209), .B2(n_1210), .Y(n_1208) );
INVx3_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1129), .B1(n_1130), .B2(n_1131), .Y(n_1127) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1128), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1330 ( .A(n_1130), .Y(n_1330) );
OAI311xp33_ASAP7_75t_L g1153 ( .A1(n_1132), .A2(n_1154), .A3(n_1158), .B1(n_1167), .C1(n_1173), .Y(n_1153) );
A2O1A1Ixp33_ASAP7_75t_L g1167 ( .A1(n_1132), .A2(n_1168), .B(n_1169), .C(n_1170), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1132), .B(n_1149), .Y(n_1183) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_1132), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1132), .B(n_1157), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1132), .B(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1132), .B(n_1231), .Y(n_1230) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1132), .B(n_1149), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1132), .B(n_1200), .Y(n_1286) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1132), .B(n_1148), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1132), .B(n_1257), .Y(n_1310) );
INVx3_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1133), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1133), .B(n_1181), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1136), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1137), .B(n_1172), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1137), .B(n_1160), .Y(n_1228) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
CKINVDCx6p67_ASAP7_75t_R g1152 ( .A(n_1139), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1139), .B(n_1187), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1139), .B(n_1160), .Y(n_1227) );
OR2x6_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1146), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1144), .B(n_1169), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1144), .B(n_1149), .Y(n_1250) );
AOI211xp5_ASAP7_75t_L g1306 ( .A1(n_1144), .A2(n_1147), .B(n_1148), .C(n_1307), .Y(n_1306) );
AND3x1_ASAP7_75t_L g1323 ( .A(n_1144), .B(n_1198), .C(n_1200), .Y(n_1323) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1148), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1147), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1147), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1147), .B(n_1279), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1147), .B(n_1261), .Y(n_1319) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1148), .Y(n_1231) );
AOI21xp33_ASAP7_75t_L g1292 ( .A1(n_1150), .A2(n_1293), .B(n_1294), .Y(n_1292) );
CKINVDCx14_ASAP7_75t_R g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1201 ( .A(n_1152), .B(n_1202), .C(n_1204), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1152), .B(n_1160), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1152), .B(n_1219), .Y(n_1284) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1157), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1157), .B(n_1181), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1157), .B(n_1277), .Y(n_1325) );
INVx3_ASAP7_75t_L g1168 ( .A(n_1159), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1159), .B(n_1186), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1159), .B(n_1195), .Y(n_1194) );
INVx5_ASAP7_75t_L g1248 ( .A(n_1159), .Y(n_1248) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_1159), .A2(n_1300), .B1(n_1312), .B2(n_1315), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1159), .B(n_1273), .Y(n_1316) );
INVx3_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1160), .B(n_1198), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1160), .B(n_1219), .Y(n_1218) );
INVx3_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1161), .B(n_1289), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1161), .B(n_1175), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1166), .Y(n_1161) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1168), .B(n_1186), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1169), .B(n_1181), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1169), .B(n_1180), .Y(n_1258) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1169), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1169), .B(n_1203), .Y(n_1329) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OAI21xp33_ASAP7_75t_L g1312 ( .A1(n_1171), .A2(n_1270), .B(n_1313), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1176), .Y(n_1173) );
AOI222xp33_ASAP7_75t_L g1253 ( .A1(n_1174), .A2(n_1193), .B1(n_1225), .B2(n_1254), .C1(n_1255), .C2(n_1258), .Y(n_1253) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1176), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_1178), .A2(n_1184), .B1(n_1188), .B2(n_1190), .Y(n_1177) );
INVxp33_ASAP7_75t_SL g1178 ( .A(n_1179), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1182), .Y(n_1179) );
INVx1_ASAP7_75t_SL g1180 ( .A(n_1181), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1181), .B(n_1224), .Y(n_1300) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
OAI32xp33_ASAP7_75t_L g1326 ( .A1(n_1185), .A2(n_1205), .A3(n_1227), .B1(n_1327), .B2(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1187), .Y(n_1199) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
AOI222xp33_ASAP7_75t_L g1302 ( .A1(n_1190), .A2(n_1284), .B1(n_1303), .B2(n_1304), .C1(n_1306), .C2(n_1309), .Y(n_1302) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1196), .B1(n_1197), .B2(n_1200), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1290 ( .A(n_1195), .B(n_1241), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1197), .B(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
A2O1A1Ixp33_ASAP7_75t_L g1291 ( .A1(n_1202), .A2(n_1251), .B(n_1292), .C(n_1296), .Y(n_1291) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1202), .Y(n_1327) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1206), .Y(n_1267) );
A2O1A1Ixp33_ASAP7_75t_L g1211 ( .A1(n_1212), .A2(n_1213), .B(n_1217), .C(n_1220), .Y(n_1211) );
AOI21xp33_ASAP7_75t_L g1320 ( .A1(n_1212), .A2(n_1264), .B(n_1293), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1215), .Y(n_1213) );
O2A1O1Ixp33_ASAP7_75t_L g1324 ( .A1(n_1215), .A2(n_1254), .B(n_1325), .C(n_1326), .Y(n_1324) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AOI221xp5_ASAP7_75t_SL g1220 ( .A1(n_1221), .A2(n_1226), .B1(n_1228), .B2(n_1229), .C(n_1232), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1222), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1223), .B(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1246 ( .A(n_1224), .B(n_1247), .C(n_1248), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_1226), .A2(n_1269), .B1(n_1271), .B2(n_1274), .C(n_1280), .Y(n_1268) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1228), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1229), .B(n_1250), .Y(n_1275) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1231), .B(n_1242), .Y(n_1241) );
INVxp67_ASAP7_75t_SL g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1234), .Y(n_1244) );
NAND5xp2_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1268), .C(n_1282), .D(n_1291), .E(n_1297), .Y(n_1235) );
AOI211xp5_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1238), .B(n_1245), .C(n_1259), .Y(n_1236) );
OAI221xp5_ASAP7_75t_L g1259 ( .A1(n_1237), .A2(n_1260), .B1(n_1262), .B2(n_1265), .C(n_1267), .Y(n_1259) );
INVxp67_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1244), .Y(n_1240) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1249), .C(n_1253), .Y(n_1245) );
NOR2xp33_ASAP7_75t_L g1262 ( .A(n_1247), .B(n_1263), .Y(n_1262) );
CKINVDCx14_ASAP7_75t_R g1296 ( .A(n_1248), .Y(n_1296) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1248), .B(n_1299), .Y(n_1298) );
A2O1A1Ixp33_ASAP7_75t_L g1321 ( .A1(n_1248), .A2(n_1250), .B(n_1322), .C(n_1323), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1252), .B(n_1281), .Y(n_1280) );
INVx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVxp67_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
O2A1O1Ixp33_ASAP7_75t_L g1317 ( .A1(n_1266), .A2(n_1287), .B(n_1318), .C(n_1320), .Y(n_1317) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1273), .Y(n_1289) );
OAI21xp33_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1276), .B(n_1278), .Y(n_1274) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1278), .Y(n_1303) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1284), .B1(n_1285), .B2(n_1287), .C(n_1290), .Y(n_1282) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1289), .Y(n_1314) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1295), .B(n_1314), .Y(n_1313) );
INVxp67_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
NAND5xp2_ASAP7_75t_SL g1301 ( .A(n_1302), .B(n_1311), .C(n_1317), .D(n_1321), .E(n_1324), .Y(n_1301) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVxp67_ASAP7_75t_SL g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx2_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1348), .Y(n_1333) );
NOR3xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1340), .C(n_1345), .Y(n_1334) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_1341), .A2(n_1342), .B1(n_1343), .B2(n_1344), .Y(n_1340) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1352), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .Y(n_1352) );
CKINVDCx16_ASAP7_75t_R g1355 ( .A(n_1356), .Y(n_1355) );
BUFx2_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVxp67_ASAP7_75t_SL g1362 ( .A(n_1363), .Y(n_1362) );
INVxp67_ASAP7_75t_SL g1386 ( .A(n_1364), .Y(n_1386) );
AND2x4_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1380), .Y(n_1364) );
NOR3xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1370), .C(n_1375), .Y(n_1365) );
OAI21xp5_ASAP7_75t_L g1366 ( .A1(n_1367), .A2(n_1368), .B(n_1369), .Y(n_1366) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVxp67_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
AND4x1_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1382), .C(n_1383), .D(n_1384), .Y(n_1380) );
HB1xp67_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
endmodule