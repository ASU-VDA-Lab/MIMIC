module fake_jpeg_2213_n_405 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_405);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_66),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_53),
.Y(n_149)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_56),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_72),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_81),
.Y(n_128)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_35),
.B(n_41),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_26),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_32),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_68),
.B1(n_76),
.B2(n_78),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_109),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_150),
.C(n_8),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_71),
.B1(n_70),
.B2(n_64),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_134),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_32),
.B1(n_34),
.B2(n_14),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_124),
.B1(n_130),
.B2(n_144),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_51),
.A2(n_32),
.B1(n_60),
.B2(n_52),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_45),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_45),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_41),
.B1(n_29),
.B2(n_30),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_28),
.B1(n_23),
.B2(n_18),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_69),
.B1(n_58),
.B2(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_53),
.B(n_23),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_9),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_28),
.B1(n_18),
.B2(n_14),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_26),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_148),
.B1(n_89),
.B2(n_67),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_90),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_46),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_168),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_46),
.B(n_47),
.C(n_54),
.D(n_62),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_127),
.A3(n_120),
.B1(n_131),
.B2(n_111),
.Y(n_195)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_162),
.Y(n_196)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_114),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_97),
.B(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_167),
.B(n_172),
.Y(n_215)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_58),
.A3(n_94),
.B1(n_65),
.B2(n_84),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_77),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_110),
.B(n_7),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_147),
.B1(n_107),
.B2(n_98),
.Y(n_219)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_139),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_149),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_182),
.Y(n_197)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_11),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_100),
.B(n_11),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_188),
.Y(n_200)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_106),
.B(n_134),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_190),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_105),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_185),
.C(n_223),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_130),
.B1(n_133),
.B2(n_118),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_185),
.B1(n_156),
.B2(n_177),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_131),
.A3(n_127),
.B1(n_115),
.B2(n_111),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_218),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_144),
.B1(n_137),
.B2(n_133),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_219),
.B1(n_169),
.B2(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_99),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_222),
.Y(n_232)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_171),
.A2(n_189),
.A3(n_154),
.B1(n_165),
.B2(n_186),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_114),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_151),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_185),
.B1(n_158),
.B2(n_174),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_227),
.B1(n_250),
.B2(n_221),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_164),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_229),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_166),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_216),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_234),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_161),
.B(n_170),
.C(n_169),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_245),
.B(n_205),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_187),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_240),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_181),
.Y(n_239)
);

AOI32xp33_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_194),
.A3(n_206),
.B1(n_204),
.B2(n_200),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_161),
.B(n_160),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_178),
.B1(n_107),
.B2(n_98),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_219),
.B1(n_207),
.B2(n_193),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_157),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_198),
.B(n_151),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_145),
.B1(n_136),
.B2(n_143),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_258),
.B1(n_265),
.B2(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_236),
.A2(n_205),
.B1(n_204),
.B2(n_213),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_259),
.A2(n_231),
.B(n_227),
.Y(n_293)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_193),
.C(n_200),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_238),
.C(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_212),
.B1(n_223),
.B2(n_209),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_265),
.B1(n_251),
.B2(n_259),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_228),
.A2(n_232),
.B1(n_239),
.B2(n_246),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_228),
.B1(n_232),
.B2(n_250),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_226),
.B1(n_248),
.B2(n_252),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_283),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_240),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_247),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_272),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_266),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_288),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_229),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_290),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_258),
.B1(n_264),
.B2(n_253),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_256),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_223),
.B(n_237),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_294),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_237),
.B(n_233),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_252),
.B(n_241),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_269),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_264),
.C(n_270),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_301),
.C(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_299),
.A2(n_317),
.B1(n_287),
.B2(n_295),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_288),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_267),
.C(n_273),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_309),
.B(n_290),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_284),
.B(n_215),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_268),
.C(n_257),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_301),
.C(n_298),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_280),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_283),
.B1(n_285),
.B2(n_294),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_276),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_234),
.B1(n_241),
.B2(n_230),
.Y(n_317)
);

XOR2x2_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_291),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g351 ( 
.A(n_319),
.B(n_304),
.CI(n_310),
.CON(n_351),
.SN(n_351)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_336),
.B1(n_304),
.B2(n_310),
.Y(n_348)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_326),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_324),
.B(n_306),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_330),
.Y(n_346)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_287),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_329),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_312),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_332),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_277),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_293),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_309),
.B(n_306),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_276),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_333),
.Y(n_339)
);

OA22x2_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_317),
.B1(n_311),
.B2(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_335),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_305),
.A2(n_286),
.B1(n_281),
.B2(n_275),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_324),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_342),
.A2(n_344),
.B(n_322),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_311),
.B(n_315),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_315),
.B(n_312),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_345),
.A2(n_332),
.B(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_348),
.A2(n_329),
.B1(n_334),
.B2(n_275),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_305),
.C(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_351),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_353),
.Y(n_367)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_334),
.B(n_319),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_356),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_318),
.C(n_325),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_357),
.B(n_358),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_347),
.A2(n_327),
.B1(n_289),
.B2(n_196),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_209),
.B1(n_208),
.B2(n_199),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_348),
.C(n_337),
.Y(n_368)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_362),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_364),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_208),
.Y(n_364)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_346),
.C(n_349),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_369),
.B(n_373),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_360),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_375),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_349),
.C(n_345),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_347),
.C(n_344),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_338),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_376),
.A2(n_356),
.B(n_351),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_371),
.B(n_352),
.C(n_355),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_SL g392 ( 
.A(n_377),
.B(n_384),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_382),
.Y(n_387)
);

OA21x2_ASAP7_75t_SL g382 ( 
.A1(n_365),
.A2(n_351),
.B(n_199),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_136),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_385),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_168),
.C(n_162),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_148),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_380),
.B(n_372),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_386),
.B(n_388),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_374),
.Y(n_388)
);

AO221x1_ASAP7_75t_L g389 ( 
.A1(n_377),
.A2(n_367),
.B1(n_146),
.B2(n_175),
.C(n_145),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_147),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_384),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_159),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_381),
.C(n_367),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_393),
.A2(n_394),
.B(n_396),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_383),
.C(n_385),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_397),
.B(n_163),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_391),
.C(n_108),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_399),
.A2(n_400),
.B(n_398),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_401),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_398),
.A2(n_108),
.B(n_190),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_402),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_132),
.Y(n_405)
);


endmodule