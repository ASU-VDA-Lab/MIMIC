module fake_jpeg_2986_n_637 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_637);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_637;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_60),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_50),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_61),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_62),
.Y(n_189)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_63),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_75),
.B(n_81),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_8),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_83),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_85),
.Y(n_210)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_27),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_90),
.Y(n_212)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_47),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_101),
.Y(n_161)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_33),
.B(n_8),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_12),
.C(n_1),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_21),
.B(n_19),
.Y(n_160)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_109),
.Y(n_202)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_32),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_115),
.A2(n_51),
.B1(n_63),
.B2(n_127),
.Y(n_190)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_45),
.B(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_52),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_132),
.B(n_15),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_57),
.B1(n_56),
.B2(n_19),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_138),
.A2(n_166),
.B1(n_190),
.B2(n_37),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_143),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_59),
.A2(n_52),
.B1(n_56),
.B2(n_21),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_140),
.A2(n_34),
.B1(n_35),
.B2(n_120),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_65),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_142),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_61),
.B(n_23),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_156),
.B(n_162),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_160),
.B(n_15),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_45),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_78),
.B(n_41),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_165),
.B(n_181),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_66),
.A2(n_56),
.B1(n_21),
.B2(n_19),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_115),
.A2(n_117),
.B1(n_128),
.B2(n_67),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_177),
.A2(n_178),
.B1(n_102),
.B2(n_37),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_64),
.A2(n_56),
.B1(n_22),
.B2(n_23),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_49),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_90),
.B(n_49),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_183),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_68),
.B(n_51),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_188),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_60),
.B(n_55),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_70),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_55),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_201),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_76),
.B(n_54),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_83),
.B(n_54),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_80),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_96),
.B(n_41),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_111),
.B(n_35),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_217),
.B(n_219),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_90),
.B(n_53),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_125),
.B(n_53),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_224),
.B(n_7),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_225),
.B(n_240),
.Y(n_321)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_227),
.Y(n_347)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_229),
.Y(n_357)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_231),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_232),
.Y(n_356)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_233),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_234),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_189),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_263),
.Y(n_311)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_131),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_242),
.Y(n_362)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_245),
.Y(n_360)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_152),
.Y(n_247)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_247),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_248),
.A2(n_277),
.B1(n_173),
.B2(n_214),
.Y(n_331)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_146),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_161),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_252),
.B(n_253),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_161),
.B(n_34),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_138),
.A2(n_124),
.B1(n_122),
.B2(n_118),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_254),
.A2(n_269),
.B(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_259),
.B(n_278),
.Y(n_364)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_260),
.Y(n_343)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_189),
.Y(n_263)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_184),
.Y(n_267)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_267),
.Y(n_359)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_268),
.A2(n_296),
.B(n_297),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_133),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_270),
.B(n_275),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_271),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_154),
.A2(n_114),
.B1(n_113),
.B2(n_108),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_272),
.A2(n_276),
.B1(n_284),
.B2(n_289),
.Y(n_340)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_274),
.Y(n_319)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_137),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_155),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_140),
.A2(n_37),
.B1(n_0),
.B2(n_4),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_187),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_137),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_281),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_13),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_282),
.Y(n_339)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_134),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_175),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_283),
.B(n_290),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_154),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_163),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_287),
.Y(n_335)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_170),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_288),
.B(n_291),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_186),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_168),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_150),
.A2(n_37),
.B1(n_3),
.B2(n_5),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_295),
.B1(n_301),
.B2(n_302),
.Y(n_344)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_298),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_166),
.A2(n_15),
.B1(n_7),
.B2(n_12),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_183),
.B(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_222),
.B(n_145),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_174),
.B(n_7),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_303),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

NAND2x1_ASAP7_75t_SL g352 ( 
.A(n_300),
.B(n_232),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_210),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_167),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_149),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_134),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_190),
.A2(n_16),
.B(n_18),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_292),
.B1(n_254),
.B2(n_269),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_307),
.A2(n_353),
.B1(n_284),
.B2(n_263),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_190),
.B1(n_147),
.B2(n_141),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_312),
.A2(n_325),
.B1(n_329),
.B2(n_331),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_164),
.C(n_171),
.Y(n_320)
);

A2O1A1O1Ixp25_ASAP7_75t_L g403 ( 
.A1(n_320),
.A2(n_351),
.B(n_358),
.C(n_242),
.D(n_244),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_246),
.A2(n_171),
.B1(n_192),
.B2(n_172),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_250),
.A2(n_194),
.B1(n_169),
.B2(n_153),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_233),
.A2(n_159),
.B(n_133),
.C(n_151),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_337),
.A2(n_303),
.B(n_258),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_153),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_345),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_208),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_272),
.A2(n_208),
.B1(n_135),
.B2(n_200),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_348),
.A2(n_355),
.B1(n_305),
.B2(n_234),
.Y(n_404)
);

FAx1_ASAP7_75t_SL g351 ( 
.A(n_228),
.B(n_159),
.CI(n_151),
.CON(n_351),
.SN(n_351)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_352),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_236),
.A2(n_195),
.B1(n_214),
.B2(n_157),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_264),
.A2(n_135),
.B1(n_200),
.B2(n_157),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_237),
.A2(n_179),
.B(n_0),
.C(n_173),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_265),
.B(n_195),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_363),
.B(n_337),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_331),
.A2(n_243),
.B1(n_289),
.B2(n_277),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_368),
.A2(n_378),
.B1(n_404),
.B2(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

NAND2x1_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_227),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_384),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_371),
.A2(n_344),
.B1(n_361),
.B2(n_320),
.Y(n_425)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_373),
.B(n_400),
.Y(n_446)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_375),
.B(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_286),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_377),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_302),
.B1(n_273),
.B2(n_281),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_352),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_323),
.A2(n_288),
.B(n_300),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_386),
.B(n_403),
.Y(n_419)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_323),
.A2(n_238),
.B(n_301),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_383),
.A2(n_391),
.B(n_399),
.Y(n_433)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_385),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g386 ( 
.A1(n_363),
.A2(n_229),
.B(n_231),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_352),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_389),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_342),
.B(n_226),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_395),
.Y(n_423)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_351),
.A2(n_230),
.B(n_235),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_393),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_330),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_310),
.B(n_294),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_401),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_397),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_398),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_312),
.A2(n_262),
.B1(n_266),
.B2(n_279),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_274),
.B1(n_270),
.B2(n_257),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_402),
.A2(n_361),
.B1(n_334),
.B2(n_319),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_316),
.B(n_287),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_321),
.B(n_338),
.Y(n_427)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_408),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_358),
.A2(n_241),
.B(n_245),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_407),
.A2(n_335),
.B(n_334),
.Y(n_437)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_411),
.Y(n_440)
);

AOI32xp33_ASAP7_75t_L g410 ( 
.A1(n_351),
.A2(n_339),
.A3(n_310),
.B1(n_350),
.B2(n_316),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_335),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_364),
.B(n_196),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_412),
.A2(n_427),
.B(n_437),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_413),
.A2(n_434),
.B1(n_438),
.B2(n_447),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_378),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_422),
.A2(n_441),
.B1(n_367),
.B2(n_387),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_396),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_424),
.B(n_435),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_425),
.A2(n_380),
.B1(n_385),
.B2(n_405),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_366),
.A2(n_341),
.B1(n_319),
.B2(n_334),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_370),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_391),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_443),
.C(n_445),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_366),
.A2(n_341),
.B1(n_319),
.B2(n_329),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_369),
.A2(n_346),
.B1(n_332),
.B2(n_322),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_370),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_367),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_322),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_359),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_404),
.A2(n_282),
.B1(n_196),
.B2(n_218),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_392),
.Y(n_471)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_452),
.Y(n_517)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_450),
.Y(n_453)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_395),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_454),
.B(n_455),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_426),
.Y(n_455)
);

AO22x2_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_381),
.B1(n_407),
.B2(n_403),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_456),
.A2(n_415),
.B1(n_442),
.B2(n_435),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_410),
.Y(n_457)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_457),
.Y(n_501)
);

AOI322xp5_ASAP7_75t_L g458 ( 
.A1(n_446),
.A2(n_373),
.A3(n_383),
.B1(n_377),
.B2(n_411),
.C1(n_388),
.C2(n_381),
.Y(n_458)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_458),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_459),
.A2(n_469),
.B1(n_434),
.B2(n_414),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_460),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_429),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_462),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_409),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_421),
.Y(n_464)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_465),
.A2(n_479),
.B1(n_481),
.B2(n_415),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_429),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_466),
.A2(n_473),
.B1(n_476),
.B2(n_477),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_422),
.A2(n_406),
.B1(n_376),
.B2(n_382),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_443),
.Y(n_470)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

XNOR2x1_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_418),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_419),
.A2(n_346),
.B(n_400),
.C(n_389),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_472),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_384),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_359),
.C(n_333),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_484),
.C(n_437),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_445),
.B(n_326),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_480),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_417),
.B(n_374),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_413),
.A2(n_390),
.B1(n_408),
.B2(n_379),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_430),
.A2(n_335),
.B(n_326),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_419),
.A2(n_360),
.B1(n_324),
.B2(n_357),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_482),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_441),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_486),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_333),
.C(n_308),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_318),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_440),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_418),
.B(n_349),
.Y(n_486)
);

XOR2x2_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_427),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_457),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_485),
.B(n_431),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_491),
.B(n_500),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_495),
.B(n_478),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_497),
.A2(n_467),
.B1(n_466),
.B2(n_460),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_431),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_498),
.B(n_512),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g502 ( 
.A(n_463),
.B(n_433),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_502),
.B(n_507),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_503),
.A2(n_510),
.B1(n_511),
.B2(n_518),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_414),
.Y(n_504)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_504),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_480),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_416),
.C(n_439),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_509),
.C(n_520),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_452),
.B(n_416),
.C(n_437),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_483),
.A2(n_416),
.B1(n_440),
.B2(n_447),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_469),
.A2(n_433),
.B1(n_448),
.B2(n_428),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_448),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_455),
.B(n_432),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_507),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_465),
.A2(n_412),
.B1(n_420),
.B2(n_432),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_457),
.C(n_459),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_523),
.B(n_541),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_524),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_532),
.C(n_537),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_511),
.A2(n_468),
.B(n_456),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_527),
.A2(n_497),
.B(n_518),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_496),
.A2(n_468),
.B1(n_478),
.B2(n_467),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_528),
.B(n_544),
.Y(n_555)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_519),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_531),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_453),
.C(n_473),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_476),
.Y(n_533)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_517),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_499),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_481),
.C(n_464),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_506),
.B(n_490),
.C(n_502),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_540),
.C(n_517),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_477),
.C(n_486),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_456),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_548),
.Y(n_551)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_515),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_545),
.B(n_479),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_513),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_546),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_R g556 ( 
.A(n_547),
.B(n_516),
.C(n_501),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_491),
.B(n_509),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_552),
.B(n_560),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_554),
.B(n_556),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_521),
.B(n_514),
.C(n_494),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_568),
.C(n_570),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_529),
.B(n_503),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_563),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_526),
.B(n_508),
.Y(n_559)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_559),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_456),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_527),
.A2(n_489),
.B(n_472),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_562),
.A2(n_543),
.B(n_522),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_525),
.B(n_456),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_510),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_564),
.B(n_522),
.Y(n_583)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_565),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_482),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_521),
.B(n_537),
.C(n_548),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_549),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_574),
.Y(n_599)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_553),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_580),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_569),
.A2(n_524),
.B1(n_528),
.B2(n_547),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_577),
.A2(n_578),
.B1(n_564),
.B2(n_560),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g578 ( 
.A1(n_561),
.A2(n_533),
.B1(n_541),
.B2(n_538),
.C(n_539),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_538),
.C(n_540),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_581),
.C(n_573),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_555),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_547),
.C(n_543),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_586),
.Y(n_595)
);

XNOR2x1_ASAP7_75t_L g591 ( 
.A(n_583),
.B(n_551),
.Y(n_591)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_585),
.B(n_588),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_569),
.A2(n_362),
.B(n_482),
.Y(n_586)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_566),
.Y(n_588)
);

NOR2xp67_ASAP7_75t_SL g610 ( 
.A(n_589),
.B(n_598),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_584),
.A2(n_554),
.B(n_557),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_590),
.A2(n_600),
.B(n_362),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_583),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_572),
.A2(n_562),
.B1(n_487),
.B2(n_568),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_592),
.B(n_596),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_577),
.A2(n_563),
.B1(n_558),
.B2(n_551),
.Y(n_593)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_593),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_570),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_567),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_567),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_602),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_581),
.B(n_487),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_587),
.C(n_576),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_603),
.B(n_598),
.C(n_601),
.Y(n_607)
);

BUFx24_ASAP7_75t_SL g604 ( 
.A(n_596),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_614),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_589),
.A2(n_582),
.B(n_586),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_605),
.A2(n_606),
.B(n_608),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_611),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_602),
.A2(n_571),
.B(n_576),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_597),
.A2(n_574),
.B(n_324),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_609),
.A2(n_347),
.B(n_318),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_613),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_349),
.C(n_343),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_617),
.A2(n_618),
.B(n_622),
.Y(n_624)
);

O2A1O1Ixp33_ASAP7_75t_SL g619 ( 
.A1(n_615),
.A2(n_594),
.B(n_595),
.C(n_599),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_619),
.A2(n_616),
.B(n_623),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_595),
.Y(n_620)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_620),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_593),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g626 ( 
.A(n_621),
.Y(n_626)
);

O2A1O1Ixp33_ASAP7_75t_SL g627 ( 
.A1(n_620),
.A2(n_606),
.B(n_591),
.C(n_327),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_SL g629 ( 
.A1(n_627),
.A2(n_327),
.B(n_356),
.C(n_347),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_628),
.B(n_343),
.C(n_218),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_629),
.A2(n_631),
.B(n_356),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_626),
.B(n_327),
.Y(n_630)
);

OAI21x1_ASAP7_75t_SL g632 ( 
.A1(n_630),
.A2(n_625),
.B(n_624),
.Y(n_632)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_632),
.A2(n_633),
.B(n_327),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_634),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_360),
.B(n_0),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_636),
.B(n_0),
.Y(n_637)
);


endmodule