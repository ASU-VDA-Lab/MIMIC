module fake_jpeg_2766_n_469 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_50),
.Y(n_145)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_57),
.B(n_92),
.Y(n_129)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_88),
.Y(n_109)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_25),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_39),
.B1(n_32),
.B2(n_15),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_11),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_96),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_95),
.B(n_38),
.Y(n_135)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_98),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_23),
.B1(n_42),
.B2(n_44),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_105),
.A2(n_114),
.B1(n_117),
.B2(n_121),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_23),
.B1(n_42),
.B2(n_44),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_128),
.B1(n_133),
.B2(n_32),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_SL g127 ( 
.A(n_77),
.Y(n_127)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_19),
.B1(n_27),
.B2(n_39),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_62),
.A2(n_29),
.B1(n_24),
.B2(n_43),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_37),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_86),
.A2(n_44),
.B1(n_37),
.B2(n_31),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_37),
.B1(n_31),
.B2(n_85),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_167),
.Y(n_202)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g218 ( 
.A(n_158),
.B(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_160),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_29),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_169),
.Y(n_203)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_43),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_183),
.Y(n_222)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_40),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_101),
.A2(n_40),
.B1(n_36),
.B2(n_30),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_170),
.A2(n_187),
.B1(n_192),
.B2(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_30),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_185),
.Y(n_207)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_98),
.B1(n_48),
.B2(n_52),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_126),
.B1(n_70),
.B2(n_59),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_46),
.B1(n_74),
.B2(n_72),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_189),
.B1(n_154),
.B2(n_114),
.Y(n_209)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_118),
.B(n_37),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_31),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_99),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_190),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_99),
.B(n_37),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_197),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_102),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_75),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_142),
.B(n_112),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_176),
.B1(n_180),
.B2(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_221),
.B1(n_175),
.B2(n_131),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_110),
.C(n_119),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_231),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_150),
.B1(n_147),
.B2(n_138),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_166),
.B1(n_178),
.B2(n_187),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_53),
.B1(n_71),
.B2(n_56),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_158),
.B(n_119),
.C(n_120),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_240),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_167),
.B1(n_158),
.B2(n_171),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_248),
.B1(n_251),
.B2(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_188),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_247),
.B1(n_249),
.B2(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_185),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_258),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_162),
.B1(n_126),
.B2(n_120),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_156),
.B1(n_151),
.B2(n_179),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_207),
.B1(n_205),
.B2(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_205),
.A2(n_210),
.B1(n_199),
.B2(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_200),
.A2(n_151),
.B1(n_47),
.B2(n_131),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_192),
.B(n_187),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_204),
.B(n_227),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_173),
.B1(n_190),
.B2(n_103),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_200),
.B1(n_212),
.B2(n_229),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_226),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_200),
.A2(n_103),
.B1(n_157),
.B2(n_198),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_200),
.A2(n_184),
.B(n_172),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_206),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_267),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_263),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_238),
.B(n_222),
.CI(n_224),
.CON(n_267),
.SN(n_267)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_237),
.B1(n_259),
.B2(n_252),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_280),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_206),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_273),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_201),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_284),
.C(n_285),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_287),
.B(n_237),
.Y(n_296)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_239),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_255),
.B(n_247),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_212),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_225),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_229),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_164),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_220),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_280),
.C(n_285),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_279),
.B1(n_271),
.B2(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_299),
.B1(n_314),
.B2(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_297),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_296),
.A2(n_311),
.B(n_273),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_255),
.B(n_248),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_286),
.B(n_227),
.Y(n_337)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_254),
.B1(n_248),
.B2(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_304),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_233),
.B1(n_244),
.B2(n_250),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_277),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_306),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_269),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_276),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_315),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_245),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_284),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_258),
.B(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_241),
.B1(n_215),
.B2(n_219),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_318),
.A2(n_337),
.B(n_307),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_334),
.B1(n_336),
.B2(n_291),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_325),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_290),
.B(n_266),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_306),
.B(n_263),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_300),
.A2(n_265),
.B1(n_270),
.B2(n_266),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_331),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_294),
.A2(n_270),
.B1(n_276),
.B2(n_287),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_260),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_340),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_308),
.A2(n_267),
.B1(n_273),
.B2(n_274),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_292),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_295),
.A2(n_267),
.B1(n_273),
.B2(n_268),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_297),
.B(n_286),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_204),
.Y(n_339)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_220),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_232),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_335),
.C(n_332),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_217),
.B(n_181),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_351),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_357),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_292),
.C(n_288),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_360),
.C(n_353),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_352),
.B1(n_362),
.B2(n_342),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_289),
.B1(n_314),
.B2(n_299),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_288),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_355),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_296),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_321),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_358),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_311),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_365),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_323),
.A2(n_303),
.B1(n_305),
.B2(n_304),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_293),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_313),
.Y(n_366)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_331),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_354),
.A2(n_317),
.B1(n_330),
.B2(n_323),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_370),
.A2(n_375),
.B1(n_380),
.B2(n_389),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_371),
.B(n_348),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_355),
.B(n_318),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_387),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_327),
.B1(n_322),
.B2(n_316),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_333),
.C(n_322),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_361),
.C(n_217),
.Y(n_398)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_333),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_351),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_312),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_219),
.B1(n_232),
.B2(n_174),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_362),
.B1(n_359),
.B2(n_365),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_404),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_395),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_359),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_394),
.Y(n_412)
);

INVx11_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_396),
.A2(n_397),
.B1(n_399),
.B2(n_0),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_370),
.A2(n_345),
.B1(n_354),
.B2(n_344),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_400),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_373),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_143),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_144),
.Y(n_402)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_144),
.C(n_143),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_407),
.C(n_381),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_144),
.B1(n_177),
.B2(n_178),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_177),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_3),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_391),
.A2(n_372),
.B(n_376),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_414),
.B(n_416),
.Y(n_430)
);

AOI21xp33_ASAP7_75t_L g414 ( 
.A1(n_405),
.A2(n_387),
.B(n_382),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_388),
.C(n_141),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_417),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_390),
.A2(n_388),
.B(n_10),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_38),
.B(n_45),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_0),
.C(n_1),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_422),
.Y(n_429)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_421),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_408),
.A2(n_7),
.B(n_1),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_0),
.C(n_1),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_424),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_1),
.C(n_2),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_2),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_393),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_431),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_412),
.B(n_406),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_407),
.C(n_403),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_434),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_410),
.B(n_404),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_419),
.C(n_409),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_436),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_396),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_2),
.Y(n_437)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_3),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_439),
.B(n_423),
.Y(n_440)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_440),
.Y(n_451)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_430),
.A2(n_419),
.B(n_422),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_442),
.B(n_446),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_415),
.Y(n_442)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_426),
.B(n_418),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_445),
.B(n_450),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_417),
.B(n_425),
.Y(n_446)
);

INVx11_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_449),
.A2(n_433),
.B(n_428),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_453),
.A2(n_454),
.B(n_4),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_448),
.A2(n_429),
.B(n_4),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_4),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_4),
.Y(n_460)
);

A2O1A1O1Ixp25_ASAP7_75t_L g458 ( 
.A1(n_452),
.A2(n_442),
.B(n_446),
.C(n_450),
.D(n_447),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_462),
.B(n_456),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_460),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_5),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_5),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_463),
.A2(n_5),
.B(n_465),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_464),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_468),
.B(n_5),
.Y(n_469)
);


endmodule