module fake_jpeg_825_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_16),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_12),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_63),
.B(n_55),
.C(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_84),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_63),
.B(n_61),
.C(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_78),
.B1(n_76),
.B2(n_59),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_107),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_111),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_112),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_70),
.A3(n_54),
.B1(n_49),
.B2(n_52),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_2),
.B(n_5),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_60),
.B1(n_70),
.B2(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_85),
.B1(n_69),
.B2(n_67),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_0),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_52),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_134),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_67),
.B(n_90),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_129),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_69),
.B1(n_20),
.B2(n_21),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_1),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_69),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_133),
.B1(n_9),
.B2(n_11),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_23),
.C(n_42),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_25),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_2),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_120),
.B1(n_115),
.B2(n_130),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_104),
.B1(n_111),
.B2(n_24),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_6),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_7),
.B(n_8),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_14),
.B(n_17),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_7),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_8),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_155),
.B1(n_18),
.B2(n_30),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_29),
.B1(n_41),
.B2(n_40),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_131),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_164),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_28),
.C(n_35),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_166),
.C(n_137),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_18),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_19),
.C(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_150),
.B1(n_154),
.B2(n_156),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_145),
.B1(n_149),
.B2(n_143),
.Y(n_176)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_150),
.C(n_155),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_171),
.C(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_159),
.B1(n_165),
.B2(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_184),
.C(n_175),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_179),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_170),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_169),
.Y(n_186)
);

OAI31xp33_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_177),
.A3(n_176),
.B(n_182),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_172),
.A3(n_166),
.B1(n_174),
.B2(n_160),
.C1(n_33),
.C2(n_32),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_189),
.C(n_47),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_192),
.Y(n_193)
);


endmodule