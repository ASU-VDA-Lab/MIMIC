module fake_netlist_6_2683_n_1974 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1974);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1974;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx8_ASAP7_75t_SL g197 ( 
.A(n_120),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_54),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_82),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_52),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_80),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_78),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_93),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_149),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_9),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_163),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_12),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_164),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_61),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_27),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_91),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_3),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_51),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_34),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_20),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_41),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_50),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_190),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_61),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_99),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_70),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_139),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_166),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_70),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_178),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_137),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_79),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_55),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_63),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_106),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_41),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_113),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_21),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_51),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_140),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_58),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_156),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_83),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_72),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_6),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_60),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_123),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_87),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_132),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_42),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_67),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_194),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_135),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_38),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_42),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_31),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_102),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_124),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_148),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_32),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_30),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_75),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_103),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_90),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_171),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_101),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_71),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_43),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_94),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_57),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_44),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_153),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_92),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_186),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_188),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_174),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_125),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_12),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_84),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_131),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_56),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_65),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_175),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_119),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_129),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_68),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_168),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_169),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_187),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_114),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_11),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_45),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_57),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_7),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_17),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_115),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_179),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_29),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_127),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_130),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_26),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_118),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_2),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_63),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_145),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_1),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_152),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_67),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_39),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_47),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_77),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_107),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_31),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_55),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_98),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_0),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_136),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_88),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_111),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_97),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_22),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_7),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_65),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_96),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_181),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_16),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_39),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_142),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_134),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_29),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_122),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_3),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_21),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_59),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_112),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_50),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_58),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_100),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_133),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_159),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_53),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_56),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_72),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_138),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_105),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_47),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_121),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_89),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_216),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_197),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_235),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_236),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_239),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_240),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_252),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_298),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_256),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_198),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_265),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_258),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_230),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_224),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_259),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_350),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_261),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_327),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_264),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_303),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_266),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_246),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_375),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_359),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_246),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_275),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_237),
.B(n_5),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_290),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_286),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_288),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_290),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_290),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_209),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_290),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_301),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_208),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_308),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_290),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_306),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_307),
.B(n_234),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_388),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_311),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_202),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_315),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_316),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_317),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_322),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_326),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_331),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_388),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_332),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_260),
.B(n_5),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_260),
.B(n_6),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_334),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_293),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_340),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_234),
.B(n_8),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_214),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_218),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_347),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_293),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_220),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_339),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_353),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_339),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_225),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_279),
.B(n_8),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_227),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_244),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_241),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_279),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_243),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_245),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_248),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_247),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_220),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_318),
.B(n_9),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_250),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_318),
.B(n_10),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_263),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_270),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_272),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_273),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_202),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_465),
.B(n_298),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_406),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_465),
.B(n_215),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_461),
.B(n_204),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_444),
.B(n_215),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_448),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_451),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_400),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_408),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_452),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_463),
.B(n_470),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_395),
.A2(n_324),
.B1(n_289),
.B2(n_367),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_471),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_403),
.A2(n_282),
.B(n_281),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_242),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_405),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_410),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_410),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_412),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_242),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_422),
.A2(n_297),
.B(n_291),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_409),
.A2(n_254),
.B1(n_285),
.B2(n_368),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_424),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_424),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_425),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_425),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_414),
.B(n_368),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_419),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_404),
.B(n_291),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g559 ( 
.A(n_450),
.B(n_262),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_480),
.B(n_204),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_432),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_428),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_428),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_430),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

AO22x1_ASAP7_75t_L g568 ( 
.A1(n_490),
.A2(n_232),
.B1(n_222),
.B2(n_392),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_468),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

CKINVDCx8_ASAP7_75t_R g571 ( 
.A(n_416),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_479),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_485),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_536),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_509),
.B(n_559),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_413),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_539),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_539),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_397),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_543),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_548),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_398),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_508),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_542),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_558),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_297),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_503),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_SL g599 ( 
.A1(n_554),
.A2(n_497),
.B1(n_454),
.B2(n_433),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_562),
.B(n_541),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_508),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_556),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_522),
.B(n_446),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_503),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_562),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_522),
.B(n_481),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_531),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_509),
.B(n_321),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_549),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_559),
.B(n_399),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_509),
.B(n_401),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_513),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_404),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_509),
.B(n_321),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_565),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_565),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_556),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_566),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_503),
.B(n_325),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_504),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_531),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_566),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_522),
.B(n_435),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_531),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_567),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_540),
.B(n_325),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_531),
.A2(n_492),
.B1(n_437),
.B2(n_466),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_558),
.B(n_402),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_504),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_549),
.B(n_407),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_558),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_549),
.B(n_411),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_520),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_526),
.B(n_198),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_549),
.B(n_415),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_549),
.Y(n_649)
);

CKINVDCx11_ASAP7_75t_R g650 ( 
.A(n_571),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

NOR2x1p5_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_396),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_504),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_528),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_528),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_549),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_541),
.B(n_511),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_511),
.B(n_417),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_568),
.B(n_420),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_533),
.Y(n_660)
);

AND2x6_ASAP7_75t_L g661 ( 
.A(n_540),
.B(n_381),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_532),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_557),
.B(n_572),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_532),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_568),
.B(n_429),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_528),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_533),
.B(n_436),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_532),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_532),
.Y(n_669)
);

BUFx4f_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_540),
.B(n_381),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_528),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_571),
.B(n_421),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_564),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_540),
.B(n_198),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_564),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_540),
.B(n_198),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_557),
.A2(n_475),
.B1(n_489),
.B2(n_443),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_535),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_530),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_512),
.B(n_198),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_564),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_533),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_535),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_535),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_R g687 ( 
.A(n_571),
.B(n_439),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_572),
.B(n_440),
.Y(n_688)
);

BUFx8_ASAP7_75t_SL g689 ( 
.A(n_527),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_512),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_512),
.B(n_199),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_504),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_527),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_573),
.B(n_472),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_504),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_554),
.B(n_445),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_551),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_512),
.B(n_199),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_L g699 ( 
.A1(n_573),
.A2(n_201),
.B1(n_295),
.B2(n_354),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_551),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_574),
.B(n_453),
.C(n_449),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_546),
.B(n_283),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_574),
.B(n_456),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_457),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_564),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_459),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_576),
.B(n_460),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_537),
.B(n_464),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_512),
.A2(n_362),
.B1(n_284),
.B2(n_310),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_534),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_537),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_537),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_577),
.B(n_474),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_577),
.B(n_474),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_546),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_538),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_SL g718 ( 
.A(n_534),
.B(n_447),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_504),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_534),
.B(n_199),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_530),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_534),
.B(n_477),
.C(n_469),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_498),
.B(n_455),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_538),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_505),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_538),
.B(n_484),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_516),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_600),
.A2(n_516),
.B1(n_534),
.B2(n_552),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_584),
.B(n_542),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_589),
.B(n_542),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_R g732 ( 
.A(n_687),
.B(n_462),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_628),
.B(n_542),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_598),
.B(n_467),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_628),
.B(n_670),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_714),
.Y(n_736)
);

AO221x1_ASAP7_75t_L g737 ( 
.A1(n_699),
.A2(n_199),
.B1(n_287),
.B2(n_371),
.C(n_376),
.Y(n_737)
);

AND2x6_ASAP7_75t_SL g738 ( 
.A(n_702),
.B(n_323),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_600),
.A2(n_516),
.B1(n_553),
.B2(n_552),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_714),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_610),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_657),
.A2(n_598),
.B1(n_607),
.B2(n_659),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_628),
.B(n_670),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_715),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_715),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_610),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_633),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_L g748 ( 
.A(n_657),
.B(n_473),
.C(n_253),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_670),
.B(n_542),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_606),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_618),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_658),
.B(n_484),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_663),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_663),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_607),
.B(n_545),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_SL g756 ( 
.A(n_673),
.B(n_202),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_633),
.B(n_545),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_694),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_637),
.A2(n_217),
.B1(n_211),
.B2(n_200),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_618),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_578),
.B(n_580),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_582),
.B(n_545),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_658),
.B(n_545),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_583),
.B(n_545),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_585),
.B(n_545),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_694),
.B(n_579),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_587),
.B(n_588),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_701),
.B(n_498),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_650),
.Y(n_769)
);

AND2x6_ASAP7_75t_SL g770 ( 
.A(n_702),
.B(n_329),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_704),
.B(n_545),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_694),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_688),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_642),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_703),
.B(n_206),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_597),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_545),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_706),
.B(n_616),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_579),
.A2(n_366),
.B1(n_231),
.B2(n_229),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_596),
.B(n_214),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_586),
.Y(n_781)
);

NOR2x1p5_ASAP7_75t_L g782 ( 
.A(n_660),
.B(n_222),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_547),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_590),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_708),
.B(n_547),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_608),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_688),
.B(n_206),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_621),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_547),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_590),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_630),
.B(n_547),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_596),
.B(n_214),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_634),
.B(n_547),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_596),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_635),
.B(n_547),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_591),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_641),
.B(n_547),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_696),
.B(n_486),
.C(n_485),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_690),
.B(n_547),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_596),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_707),
.B(n_575),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_595),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_591),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_644),
.B(n_550),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_707),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_690),
.B(n_550),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_693),
.A2(n_199),
.B1(n_287),
.B2(n_371),
.C(n_383),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_722),
.B(n_203),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_648),
.B(n_550),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_647),
.A2(n_563),
.B(n_561),
.C(n_553),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_639),
.B(n_550),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_602),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_681),
.A2(n_516),
.B(n_552),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_601),
.B(n_207),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_662),
.B(n_550),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_664),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_668),
.B(n_550),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_601),
.B(n_207),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_602),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_690),
.B(n_710),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_669),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_674),
.B(n_550),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_710),
.B(n_550),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_677),
.B(n_552),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_710),
.B(n_287),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_683),
.B(n_553),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_667),
.B(n_486),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_603),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_659),
.A2(n_304),
.B1(n_341),
.B2(n_333),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_603),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_647),
.A2(n_553),
.B(n_563),
.C(n_561),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_705),
.B(n_561),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_721),
.B(n_561),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_726),
.B(n_563),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_665),
.A2(n_328),
.B1(n_319),
.B2(n_343),
.Y(n_836)
);

BUFx5_ASAP7_75t_L g837 ( 
.A(n_596),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_619),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_619),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_711),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_649),
.B(n_563),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_606),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_665),
.B(n_287),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_713),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_625),
.B(n_205),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_723),
.B(n_287),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_605),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_717),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_724),
.Y(n_849)
);

NOR2x1_ASAP7_75t_L g850 ( 
.A(n_652),
.B(n_219),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_605),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_649),
.B(n_530),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_656),
.B(n_530),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_684),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_613),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_614),
.A2(n_679),
.B1(n_581),
.B2(n_656),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_636),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_613),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_625),
.A2(n_544),
.B1(n_280),
.B2(n_226),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_606),
.B(n_487),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_581),
.B(n_487),
.Y(n_861)
);

AO221x1_ASAP7_75t_L g862 ( 
.A1(n_592),
.A2(n_371),
.B1(n_335),
.B2(n_337),
.C(n_345),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_625),
.B(n_530),
.Y(n_863)
);

AOI221xp5_ASAP7_75t_L g864 ( 
.A1(n_599),
.A2(n_360),
.B1(n_392),
.B2(n_389),
.C(n_294),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_606),
.B(n_575),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_594),
.B(n_210),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_625),
.B(n_530),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_636),
.A2(n_524),
.B(n_518),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_625),
.A2(n_544),
.B1(n_228),
.B2(n_296),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_210),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_609),
.B(n_212),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_617),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_609),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_SL g874 ( 
.A(n_660),
.B(n_269),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_612),
.B(n_371),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_612),
.B(n_371),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_625),
.B(n_530),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_596),
.B(n_530),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_611),
.B(n_524),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_626),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_612),
.B(n_214),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_611),
.B(n_524),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_626),
.B(n_214),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_617),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_629),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_629),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_638),
.B(n_214),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_638),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_631),
.A2(n_302),
.B1(n_344),
.B2(n_351),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_645),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_609),
.B(n_491),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_645),
.B(n_214),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_654),
.B(n_214),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_611),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_675),
.A2(n_524),
.B(n_518),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_611),
.B(n_524),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_611),
.B(n_500),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_778),
.B(n_611),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_757),
.A2(n_655),
.B(n_654),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_797),
.A2(n_651),
.B(n_632),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_773),
.B(n_609),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_766),
.A2(n_631),
.B1(n_671),
.B2(n_661),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_828),
.B(n_661),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_804),
.A2(n_651),
.B(n_632),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_801),
.B(n_631),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_759),
.A2(n_675),
.B(n_678),
.C(n_720),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_885),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_809),
.A2(n_651),
.B(n_632),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_775),
.A2(n_702),
.B(n_631),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_801),
.B(n_661),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_734),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_733),
.A2(n_653),
.B(n_640),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_861),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_787),
.A2(n_544),
.B(n_678),
.C(n_314),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_751),
.B(n_760),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_751),
.B(n_760),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_802),
.B(n_661),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_733),
.A2(n_653),
.B(n_640),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_SL g919 ( 
.A(n_854),
.B(n_604),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_774),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_773),
.B(n_805),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_805),
.B(n_622),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_776),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_741),
.B(n_661),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_860),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_815),
.B(n_650),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_837),
.B(n_640),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_742),
.B(n_702),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_891),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_843),
.A2(n_698),
.B(n_682),
.C(n_720),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_741),
.B(n_746),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_837),
.B(n_640),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_746),
.B(n_661),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_808),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_747),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_819),
.A2(n_294),
.B(n_232),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_747),
.B(n_671),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_894),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_766),
.B(n_671),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_766),
.B(n_671),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_786),
.B(n_716),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_885),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_894),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_749),
.A2(n_653),
.B(n_640),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_749),
.A2(n_692),
.B(n_653),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_846),
.A2(n_843),
.B(n_731),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_865),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_730),
.A2(n_692),
.B(n_653),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_SL g949 ( 
.A(n_756),
.B(n_689),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_753),
.B(n_491),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_886),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_754),
.B(n_493),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_811),
.A2(n_725),
.B(n_692),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_837),
.B(n_692),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_837),
.B(n_692),
.Y(n_955)
);

BUFx8_ASAP7_75t_SL g956 ( 
.A(n_769),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_757),
.A2(n_725),
.B(n_593),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_L g958 ( 
.A1(n_752),
.A2(n_372),
.B(n_360),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_788),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_736),
.B(n_671),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_894),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_735),
.A2(n_725),
.B(n_593),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_886),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_735),
.A2(n_725),
.B(n_593),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_763),
.A2(n_728),
.B(n_691),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_738),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_856),
.B(n_655),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_743),
.A2(n_725),
.B(n_593),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_SL g969 ( 
.A(n_864),
.B(n_373),
.C(n_372),
.Y(n_969)
);

BUFx4f_ASAP7_75t_L g970 ( 
.A(n_842),
.Y(n_970)
);

BUFx12f_ASAP7_75t_L g971 ( 
.A(n_770),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_729),
.A2(n_672),
.B(n_666),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_838),
.A2(n_292),
.B(n_271),
.C(n_357),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_748),
.B(n_213),
.C(n_212),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_890),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_740),
.B(n_744),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_745),
.B(n_671),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_839),
.A2(n_709),
.B1(n_394),
.B2(n_365),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_837),
.B(n_592),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_870),
.A2(n_364),
.B(n_363),
.C(n_233),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_743),
.A2(n_593),
.B(n_592),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_863),
.A2(n_643),
.B(n_627),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_837),
.B(n_627),
.Y(n_983)
);

AOI33xp33_ASAP7_75t_L g984 ( 
.A1(n_808),
.A2(n_496),
.A3(n_495),
.B1(n_494),
.B2(n_493),
.B3(n_342),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_794),
.A2(n_255),
.B1(n_251),
.B2(n_238),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_763),
.B(n_666),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_761),
.B(n_672),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_739),
.A2(n_680),
.B(n_676),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_867),
.A2(n_643),
.B(n_627),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_782),
.B(n_643),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_767),
.B(n_676),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_865),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_814),
.A2(n_685),
.B(n_680),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_877),
.A2(n_719),
.B(n_695),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_890),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_758),
.B(n_685),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_785),
.A2(n_719),
.B(n_695),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_866),
.B(n_494),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_834),
.A2(n_697),
.B(n_686),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_737),
.A2(n_369),
.B1(n_352),
.B2(n_348),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_772),
.B(n_686),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_894),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_871),
.B(n_697),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_835),
.B(n_700),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_808),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_874),
.A2(n_779),
.B(n_798),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_812),
.B(n_700),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_817),
.B(n_712),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_830),
.B(n_257),
.C(n_249),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_836),
.B(n_221),
.C(n_213),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_794),
.A2(n_623),
.B1(n_682),
.B2(n_691),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_837),
.B(n_800),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_822),
.B(n_712),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_785),
.A2(n_771),
.B(n_852),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_846),
.B(n_727),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_878),
.A2(n_719),
.B(n_695),
.Y(n_1017)
);

AO21x1_ASAP7_75t_L g1018 ( 
.A1(n_771),
.A2(n_826),
.B(n_881),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_853),
.A2(n_698),
.B(n_727),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_873),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_755),
.A2(n_514),
.B(n_500),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_732),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_768),
.B(n_495),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_799),
.A2(n_518),
.B(n_505),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_873),
.B(n_496),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_755),
.A2(n_501),
.B(n_502),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_800),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_845),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_840),
.B(n_623),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_889),
.B(n_844),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_848),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_849),
.B(n_623),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_873),
.B(n_623),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_781),
.B(n_501),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_845),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_799),
.A2(n_518),
.B(n_505),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_781),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_784),
.B(n_502),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_769),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_784),
.B(n_506),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_806),
.A2(n_518),
.B(n_505),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_850),
.B(n_476),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_806),
.A2(n_518),
.B(n_505),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_859),
.A2(n_869),
.B1(n_821),
.B2(n_824),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_790),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_824),
.A2(n_518),
.B(n_505),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_790),
.B(n_506),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_821),
.B(n_845),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_826),
.B(n_476),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_750),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_796),
.B(n_803),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_762),
.A2(n_764),
.B(n_765),
.C(n_777),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_796),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_825),
.A2(n_521),
.B(n_515),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_883),
.A2(n_517),
.B(n_507),
.C(n_529),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_L g1056 ( 
.A(n_880),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_827),
.A2(n_521),
.B(n_515),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_750),
.B(n_267),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_783),
.A2(n_229),
.B(n_231),
.C(n_223),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_881),
.A2(n_519),
.B(n_507),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_833),
.A2(n_525),
.B(n_514),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_883),
.A2(n_892),
.B(n_887),
.C(n_893),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_803),
.B(n_510),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_750),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_813),
.B(n_510),
.Y(n_1065)
);

NAND2x1_ASAP7_75t_L g1066 ( 
.A(n_813),
.B(n_820),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_879),
.A2(n_505),
.B(n_518),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_820),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_882),
.A2(n_505),
.B(n_499),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_896),
.B(n_221),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_829),
.B(n_517),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_841),
.A2(n_499),
.B(n_523),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_829),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_887),
.A2(n_519),
.B(n_529),
.C(n_525),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_897),
.B(n_689),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_807),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_875),
.A2(n_523),
.B(n_499),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_789),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_831),
.B(n_575),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_831),
.B(n_223),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_875),
.A2(n_523),
.B(n_499),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_876),
.A2(n_792),
.B(n_780),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_847),
.B(n_358),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_892),
.A2(n_523),
.B(n_499),
.C(n_478),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_847),
.B(n_358),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_791),
.A2(n_478),
.B(n_523),
.Y(n_1086)
);

OR2x2_ASAP7_75t_SL g1087 ( 
.A(n_793),
.B(n_269),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_1002),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1082),
.A2(n_780),
.B(n_792),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_998),
.B(n_862),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_911),
.B(n_795),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_SL g1092 ( 
.A1(n_1070),
.A2(n_893),
.B(n_876),
.C(n_888),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1062),
.A2(n_1015),
.B(n_914),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_913),
.B(n_816),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_947),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1002),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_922),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_947),
.Y(n_1098)
);

OAI21xp33_ASAP7_75t_L g1099 ( 
.A1(n_936),
.A2(n_373),
.B(n_378),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_928),
.A2(n_382),
.B1(n_380),
.B2(n_379),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1020),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_928),
.A2(n_810),
.B(n_832),
.C(n_823),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_992),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_951),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_898),
.A2(n_818),
.B(n_868),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_925),
.B(n_851),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_992),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_923),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_913),
.A2(n_851),
.B1(n_884),
.B2(n_872),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_905),
.B(n_268),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_929),
.B(n_274),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1007),
.A2(n_895),
.B(n_884),
.C(n_872),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_909),
.B(n_380),
.C(n_378),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_911),
.B(n_855),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_976),
.A2(n_858),
.B1(n_855),
.B2(n_379),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_949),
.B(n_269),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_925),
.B(n_858),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_959),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1006),
.B(n_361),
.Y(n_1119)
);

CKINVDCx14_ASAP7_75t_R g1120 ( 
.A(n_1039),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1006),
.B(n_361),
.Y(n_1121)
);

AOI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1076),
.A2(n_366),
.B1(n_393),
.B2(n_391),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_910),
.A2(n_385),
.B(n_393),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_903),
.A2(n_385),
.B(n_391),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1003),
.B(n_569),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_900),
.A2(n_390),
.B(n_386),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_904),
.A2(n_390),
.B(n_386),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1003),
.B(n_569),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_951),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_934),
.B(n_370),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_921),
.B(n_276),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_908),
.A2(n_384),
.B(n_377),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_939),
.A2(n_384),
.B(n_377),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_929),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1005),
.A2(n_382),
.B1(n_389),
.B2(n_387),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_963),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_963),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_906),
.A2(n_930),
.B(n_967),
.C(n_901),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_L g1139 ( 
.A(n_969),
.B(n_320),
.C(n_278),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_967),
.A2(n_370),
.B(n_374),
.C(n_277),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_921),
.B(n_374),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_SL g1142 ( 
.A1(n_1018),
.A2(n_196),
.B(n_195),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1044),
.A2(n_387),
.B1(n_330),
.B2(n_356),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_966),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_919),
.B(n_349),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_987),
.B(n_569),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_974),
.A2(n_158),
.B(n_76),
.C(n_81),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_970),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_940),
.A2(n_569),
.B(n_184),
.Y(n_1150)
);

INVx3_ASAP7_75t_SL g1151 ( 
.A(n_1022),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_927),
.A2(n_569),
.B(n_172),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_SL g1153 ( 
.A(n_956),
.B(n_299),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_SL g1154 ( 
.A(n_1050),
.B(n_313),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_991),
.B(n_569),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_935),
.B(n_569),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_995),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_938),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1078),
.B(n_569),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_958),
.A2(n_346),
.B(n_338),
.Y(n_1160)
);

BUFx8_ASAP7_75t_L g1161 ( 
.A(n_971),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_990),
.B(n_154),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_927),
.A2(n_128),
.B(n_85),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_941),
.B(n_336),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_901),
.B(n_1056),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1062),
.A2(n_312),
.B(n_309),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_935),
.B(n_305),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_926),
.B(n_300),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1056),
.B(n_147),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_915),
.B(n_916),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1075),
.B(n_116),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_995),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1027),
.B(n_931),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1025),
.B(n_10),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1027),
.B(n_110),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1004),
.B(n_74),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_907),
.B(n_11),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_970),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1045),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_950),
.B(n_13),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_950),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_942),
.B(n_14),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_975),
.B(n_16),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_941),
.B(n_1058),
.C(n_1010),
.Y(n_1184)
);

OAI21xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1013),
.A2(n_17),
.B(n_18),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_974),
.B(n_18),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_997),
.A2(n_19),
.B(n_20),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_R g1188 ( 
.A(n_1050),
.B(n_73),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_932),
.A2(n_73),
.B(n_23),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_952),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_920),
.B(n_19),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_952),
.B(n_1023),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1031),
.B(n_23),
.Y(n_1193)
);

AO32x1_ASAP7_75t_L g1194 ( 
.A1(n_985),
.A2(n_24),
.A3(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1030),
.A2(n_24),
.B(n_30),
.C(n_33),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_938),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_938),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_954),
.A2(n_71),
.B(n_34),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_954),
.A2(n_69),
.B(n_36),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1049),
.B(n_984),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_938),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1011),
.B(n_33),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1042),
.B(n_36),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_SL g1204 ( 
.A(n_1011),
.B(n_69),
.C(n_38),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1023),
.B(n_1058),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_955),
.A2(n_68),
.B(n_40),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_943),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_955),
.A2(n_37),
.B(n_40),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1052),
.A2(n_37),
.B(n_45),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1053),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1064),
.B(n_48),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1023),
.B(n_48),
.Y(n_1212)
);

BUFx4f_ASAP7_75t_L g1213 ( 
.A(n_1028),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_924),
.A2(n_49),
.B(n_52),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1070),
.A2(n_66),
.B1(n_53),
.B2(n_59),
.Y(n_1215)
);

O2A1O1Ixp5_ASAP7_75t_L g1216 ( 
.A1(n_946),
.A2(n_49),
.B(n_60),
.C(n_62),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_SL g1217 ( 
.A(n_980),
.B(n_62),
.C(n_64),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_902),
.A2(n_64),
.B(n_66),
.C(n_960),
.Y(n_1218)
);

AO32x1_ASAP7_75t_L g1219 ( 
.A1(n_978),
.A2(n_1012),
.A3(n_1068),
.B1(n_1073),
.B2(n_1000),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_943),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1042),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1064),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_943),
.B(n_961),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_SL g1224 ( 
.A1(n_1054),
.A2(n_1057),
.B(n_1061),
.C(n_993),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_996),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_933),
.A2(n_937),
.B(n_948),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1000),
.A2(n_943),
.B1(n_961),
.B2(n_1048),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1013),
.A2(n_953),
.B(n_979),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_979),
.A2(n_983),
.B(n_912),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_977),
.A2(n_1016),
.B(n_917),
.C(n_1059),
.Y(n_1231)
);

NAND2xp33_ASAP7_75t_R g1232 ( 
.A(n_1033),
.B(n_986),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1087),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_961),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_961),
.B(n_1051),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1001),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1016),
.A2(n_1033),
.B(n_999),
.C(n_972),
.Y(n_1237)
);

AO22x1_ASAP7_75t_L g1238 ( 
.A1(n_1028),
.A2(n_1035),
.B1(n_1085),
.B2(n_1029),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1239)
);

OA22x2_ASAP7_75t_L g1240 ( 
.A1(n_899),
.A2(n_983),
.B1(n_988),
.B2(n_1014),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1028),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_918),
.A2(n_944),
.B(n_945),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1035),
.B(n_1048),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1034),
.B(n_1047),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1038),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_982),
.A2(n_994),
.B(n_989),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1226),
.A2(n_965),
.B(n_1021),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1213),
.B(n_1035),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1138),
.A2(n_1019),
.B(n_1074),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1164),
.B(n_1032),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1134),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1089),
.A2(n_1237),
.B(n_1246),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1242),
.A2(n_1026),
.B(n_981),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1209),
.A2(n_973),
.B(n_1066),
.C(n_1065),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1228),
.A2(n_1067),
.B(n_962),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1151),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1146),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1102),
.A2(n_1060),
.A3(n_964),
.B(n_968),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1213),
.B(n_1088),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1139),
.A2(n_1071),
.B1(n_1040),
.B2(n_1063),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1093),
.A2(n_1069),
.B(n_1079),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1149),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1093),
.A2(n_957),
.B(n_1024),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1184),
.B(n_1131),
.C(n_1116),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1101),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1202),
.A2(n_1055),
.B(n_1074),
.C(n_1084),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1244),
.A2(n_1036),
.B(n_1041),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1230),
.A2(n_1105),
.B(n_1240),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1231),
.A2(n_1072),
.A3(n_1046),
.B(n_1043),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1118),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1209),
.A2(n_1086),
.B(n_1084),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1244),
.A2(n_1077),
.B(n_1081),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1218),
.A2(n_1227),
.A3(n_1112),
.B(n_1125),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1224),
.A2(n_1092),
.B(n_1240),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1176),
.A2(n_1128),
.B(n_1125),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1176),
.A2(n_1239),
.B(n_1128),
.Y(n_1277)
);

O2A1O1Ixp5_ASAP7_75t_L g1278 ( 
.A1(n_1238),
.A2(n_1165),
.B(n_1166),
.C(n_1216),
.Y(n_1278)
);

NAND3x1_ASAP7_75t_L g1279 ( 
.A(n_1205),
.B(n_1212),
.C(n_1215),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1239),
.A2(n_1227),
.B(n_1155),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1192),
.B(n_1181),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1147),
.A2(n_1155),
.A3(n_1115),
.B(n_1195),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1158),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1159),
.A2(n_1219),
.B(n_1173),
.Y(n_1284)
);

NAND3x1_ASAP7_75t_L g1285 ( 
.A(n_1180),
.B(n_1168),
.C(n_1203),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1219),
.A2(n_1173),
.B(n_1229),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1219),
.A2(n_1245),
.B(n_1235),
.Y(n_1287)
);

CKINVDCx8_ASAP7_75t_R g1288 ( 
.A(n_1178),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1095),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1113),
.A2(n_1140),
.B(n_1090),
.C(n_1166),
.Y(n_1290)
);

AO21x1_ASAP7_75t_L g1291 ( 
.A1(n_1189),
.A2(n_1206),
.B(n_1198),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1222),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1143),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1199),
.A2(n_1208),
.B(n_1214),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1200),
.A2(n_1185),
.B(n_1160),
.C(n_1099),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1243),
.A2(n_1235),
.B(n_1091),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1175),
.A2(n_1150),
.B(n_1156),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1098),
.B(n_1103),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1186),
.A2(n_1204),
.B(n_1144),
.C(n_1217),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1221),
.B(n_1107),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1179),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1175),
.A2(n_1114),
.B(n_1170),
.Y(n_1303)
);

AOI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1144),
.A2(n_1100),
.B1(n_1135),
.B2(n_1233),
.C(n_1115),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1187),
.A2(n_1152),
.B(n_1109),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1211),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1109),
.A2(n_1142),
.B(n_1183),
.Y(n_1307)
);

OAI22x1_ASAP7_75t_L g1308 ( 
.A1(n_1122),
.A2(n_1211),
.B1(n_1174),
.B2(n_1162),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1094),
.A2(n_1124),
.B(n_1193),
.C(n_1191),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_SL g1310 ( 
.A(n_1154),
.B(n_1153),
.C(n_1121),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1190),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1141),
.B(n_1119),
.C(n_1130),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1148),
.A2(n_1171),
.B(n_1135),
.C(n_1167),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1177),
.A2(n_1182),
.B(n_1163),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1126),
.A2(n_1132),
.A3(n_1127),
.B(n_1123),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1169),
.A2(n_1223),
.B(n_1167),
.C(n_1241),
.Y(n_1316)
);

AOI221x1_ASAP7_75t_L g1317 ( 
.A1(n_1133),
.A2(n_1162),
.B1(n_1194),
.B2(n_1106),
.C(n_1117),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1210),
.A2(n_1129),
.B(n_1157),
.C(n_1104),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_SL g1319 ( 
.A(n_1158),
.B(n_1234),
.Y(n_1319)
);

AOI31xp67_ASAP7_75t_L g1320 ( 
.A1(n_1136),
.A2(n_1172),
.A3(n_1137),
.B(n_1106),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1088),
.A2(n_1096),
.B(n_1232),
.C(n_1194),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1196),
.B(n_1220),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1120),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1194),
.A2(n_1220),
.B(n_1207),
.C(n_1196),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1188),
.B(n_1207),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1158),
.A2(n_1234),
.A3(n_1197),
.B(n_1201),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1197),
.A2(n_1201),
.B(n_1145),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1197),
.A2(n_1201),
.B(n_1145),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1161),
.A2(n_928),
.B1(n_1144),
.B2(n_1164),
.C(n_864),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1161),
.B(n_1225),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1164),
.A2(n_778),
.B(n_1007),
.C(n_775),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1138),
.A2(n_1224),
.B(n_1102),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1108),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1209),
.A2(n_778),
.B1(n_928),
.B2(n_1138),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1134),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1108),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1108),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_SL g1339 ( 
.A(n_1178),
.B(n_1022),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1178),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1138),
.A2(n_946),
.A3(n_1018),
.B(n_967),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_1134),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1108),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1093),
.A2(n_1138),
.B(n_1209),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1202),
.A2(n_775),
.B(n_1164),
.C(n_1186),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_804),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1138),
.A2(n_946),
.A3(n_1018),
.B(n_967),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1138),
.A2(n_946),
.A3(n_1018),
.B(n_967),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_L g1353 ( 
.A(n_1164),
.B(n_775),
.C(n_778),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1134),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1142),
.A2(n_1209),
.B(n_1198),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1178),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1097),
.B(n_911),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1164),
.A2(n_778),
.B(n_1007),
.C(n_775),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1134),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1149),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1093),
.A2(n_1138),
.B(n_1246),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1366)
);

AO21x1_ASAP7_75t_L g1367 ( 
.A1(n_1209),
.A2(n_846),
.B(n_1227),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1138),
.A2(n_946),
.A3(n_1018),
.B(n_967),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1108),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1134),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1164),
.A2(n_716),
.B1(n_556),
.B2(n_928),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1108),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1164),
.B(n_395),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_SL g1379 ( 
.A1(n_1138),
.A2(n_1209),
.B(n_1218),
.C(n_1169),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1138),
.A2(n_946),
.A3(n_1018),
.B(n_967),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1178),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1134),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1238),
.A2(n_1128),
.B(n_1125),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1110),
.B(n_828),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_1138),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1138),
.A2(n_1224),
.B(n_1102),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1164),
.B(n_395),
.Y(n_1387)
);

BUFx12f_ASAP7_75t_L g1388 ( 
.A(n_1145),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1389)
);

BUFx8_ASAP7_75t_SL g1390 ( 
.A(n_1178),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1089),
.A2(n_1082),
.B(n_804),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1108),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1134),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1108),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1164),
.B(n_775),
.C(n_778),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1134),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1093),
.A2(n_1138),
.B(n_1209),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1226),
.A2(n_1017),
.B(n_1242),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1088),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1134),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1213),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1225),
.B(n_1236),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1340),
.Y(n_1403)
);

CKINVDCx6p67_ASAP7_75t_R g1404 ( 
.A(n_1388),
.Y(n_1404)
);

INVx8_ASAP7_75t_L g1405 ( 
.A(n_1390),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1335),
.A2(n_1395),
.B1(n_1353),
.B2(n_1329),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1271),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1337),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1401),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1358),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1393),
.Y(n_1412)
);

INVx8_ASAP7_75t_L g1413 ( 
.A(n_1281),
.Y(n_1413)
);

INVx8_ASAP7_75t_L g1414 ( 
.A(n_1281),
.Y(n_1414)
);

BUFx4_ASAP7_75t_R g1415 ( 
.A(n_1257),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1375),
.A2(n_1387),
.B1(n_1378),
.B2(n_1264),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1329),
.A2(n_1335),
.B1(n_1304),
.B2(n_1384),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1381),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1304),
.A2(n_1250),
.B1(n_1301),
.B2(n_1310),
.Y(n_1419)
);

INVx8_ASAP7_75t_L g1420 ( 
.A(n_1300),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1279),
.A2(n_1285),
.B1(n_1312),
.B2(n_1362),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1283),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1306),
.B(n_1300),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1367),
.A2(n_1397),
.B1(n_1345),
.B2(n_1257),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1346),
.A2(n_1299),
.B(n_1331),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1256),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1325),
.A2(n_1330),
.B1(n_1402),
.B2(n_1266),
.Y(n_1428)
);

BUFx4f_ASAP7_75t_SL g1429 ( 
.A(n_1262),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1265),
.Y(n_1430)
);

OAI22x1_ASAP7_75t_SL g1431 ( 
.A1(n_1364),
.A2(n_1382),
.B1(n_1400),
.B2(n_1394),
.Y(n_1431)
);

BUFx10_ASAP7_75t_L g1432 ( 
.A(n_1251),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1283),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1248),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1334),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1266),
.A2(n_1348),
.B1(n_1366),
.B2(n_1347),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1325),
.A2(n_1330),
.B1(n_1355),
.B2(n_1348),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1347),
.A2(n_1402),
.B1(n_1366),
.B2(n_1355),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1345),
.A2(n_1397),
.B1(n_1333),
.B2(n_1386),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1338),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1259),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1371),
.A2(n_1308),
.B1(n_1288),
.B2(n_1292),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1328),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1371),
.A2(n_1386),
.B(n_1333),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1344),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1323),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1400),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1298),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1248),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1311),
.A2(n_1360),
.B1(n_1372),
.B2(n_1396),
.Y(n_1450)
);

INVx11_ASAP7_75t_L g1451 ( 
.A(n_1339),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1392),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1290),
.A2(n_1379),
.B1(n_1342),
.B2(n_1291),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1289),
.A2(n_1302),
.B1(n_1293),
.B2(n_1295),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1277),
.B(n_1280),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1309),
.A2(n_1294),
.B1(n_1260),
.B2(n_1356),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1280),
.A2(n_1277),
.B1(n_1376),
.B2(n_1332),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1357),
.A2(n_1365),
.B1(n_1336),
.B2(n_1249),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1319),
.Y(n_1459)
);

INVx8_ASAP7_75t_L g1460 ( 
.A(n_1399),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1296),
.B(n_1341),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1327),
.Y(n_1462)
);

BUFx8_ASAP7_75t_L g1463 ( 
.A(n_1327),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1326),
.Y(n_1464)
);

BUFx4f_ASAP7_75t_SL g1465 ( 
.A(n_1399),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1316),
.Y(n_1466)
);

AOI22x1_ASAP7_75t_SL g1467 ( 
.A1(n_1313),
.A2(n_1278),
.B1(n_1322),
.B2(n_1317),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1365),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1320),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1303),
.A2(n_1343),
.B1(n_1359),
.B2(n_1332),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1303),
.A2(n_1376),
.B1(n_1359),
.B2(n_1370),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1322),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1326),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1343),
.A2(n_1370),
.B1(n_1385),
.B2(n_1249),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1318),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1286),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1341),
.Y(n_1477)
);

INVx2_ASAP7_75t_R g1478 ( 
.A(n_1324),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1385),
.A2(n_1286),
.B1(n_1307),
.B2(n_1252),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1351),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1276),
.A2(n_1287),
.B1(n_1383),
.B2(n_1297),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1275),
.Y(n_1482)
);

CKINVDCx14_ASAP7_75t_R g1483 ( 
.A(n_1321),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1252),
.A2(n_1275),
.B1(n_1314),
.B2(n_1276),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1263),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1351),
.Y(n_1486)
);

CKINVDCx6p67_ASAP7_75t_R g1487 ( 
.A(n_1254),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1351),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1287),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1284),
.A2(n_1261),
.B1(n_1267),
.B2(n_1263),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1297),
.A2(n_1273),
.B1(n_1261),
.B2(n_1269),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1273),
.A2(n_1272),
.B1(n_1284),
.B2(n_1268),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1272),
.A2(n_1268),
.B1(n_1305),
.B2(n_1391),
.Y(n_1493)
);

CKINVDCx10_ASAP7_75t_R g1494 ( 
.A(n_1282),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1349),
.A2(n_1274),
.B1(n_1380),
.B2(n_1368),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1247),
.A2(n_1255),
.B1(n_1253),
.B2(n_1389),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1350),
.A2(n_1354),
.B1(n_1374),
.B2(n_1373),
.Y(n_1497)
);

OAI22x1_ASAP7_75t_SL g1498 ( 
.A1(n_1282),
.A2(n_1352),
.B1(n_1380),
.B2(n_1368),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1361),
.A2(n_1398),
.B1(n_1380),
.B2(n_1352),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1274),
.A2(n_1282),
.B1(n_1315),
.B2(n_1258),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1274),
.A2(n_1258),
.B1(n_1315),
.B2(n_1270),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1315),
.A2(n_1258),
.B1(n_1270),
.B2(n_1378),
.Y(n_1502)
);

BUFx2_ASAP7_75t_SL g1503 ( 
.A(n_1288),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1375),
.A2(n_756),
.B1(n_1395),
.B2(n_1353),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1335),
.A2(n_1395),
.B1(n_1353),
.B2(n_1329),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1256),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1335),
.A2(n_1395),
.B1(n_1353),
.B2(n_1329),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1353),
.A2(n_756),
.B1(n_1395),
.B2(n_874),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1340),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1353),
.A2(n_1395),
.B1(n_1329),
.B2(n_1264),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1375),
.A2(n_756),
.B1(n_1395),
.B2(n_1353),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1388),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1375),
.A2(n_1335),
.B1(n_756),
.B2(n_874),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1353),
.A2(n_1395),
.B1(n_1329),
.B2(n_1264),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1353),
.A2(n_1395),
.B1(n_1329),
.B2(n_1264),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1271),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1340),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1271),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1335),
.A2(n_756),
.B1(n_874),
.B2(n_1116),
.Y(n_1519)
);

BUFx12f_ASAP7_75t_L g1520 ( 
.A(n_1256),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1335),
.B(n_1266),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1353),
.A2(n_1395),
.B1(n_1329),
.B2(n_1264),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1340),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1340),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1378),
.A2(n_716),
.B1(n_1387),
.B2(n_599),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1340),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1340),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1363),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1335),
.B(n_1266),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_1256),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1401),
.Y(n_1531)
);

CKINVDCx11_ASAP7_75t_R g1532 ( 
.A(n_1388),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1335),
.A2(n_1362),
.B(n_1331),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1353),
.A2(n_756),
.B1(n_1395),
.B2(n_874),
.Y(n_1534)
);

CKINVDCx12_ASAP7_75t_R g1535 ( 
.A(n_1301),
.Y(n_1535)
);

INVx3_ASAP7_75t_SL g1536 ( 
.A(n_1262),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1375),
.A2(n_756),
.B1(n_1395),
.B2(n_1353),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1375),
.A2(n_1335),
.B1(n_756),
.B2(n_874),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1378),
.A2(n_1387),
.B1(n_1395),
.B2(n_1353),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1353),
.A2(n_1395),
.B1(n_1329),
.B2(n_1264),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1477),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1473),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1486),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1488),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1438),
.B(n_1428),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1512),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1457),
.A2(n_1455),
.B(n_1474),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1464),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1436),
.B(n_1510),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1448),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1469),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1435),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1445),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1461),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1497),
.A2(n_1496),
.B(n_1493),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1468),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1443),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.B(n_1502),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1481),
.A2(n_1490),
.B(n_1455),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1440),
.B(n_1452),
.Y(n_1562)
);

OA21x2_ASAP7_75t_L g1563 ( 
.A1(n_1479),
.A2(n_1492),
.B(n_1491),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1539),
.B(n_1525),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1461),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1458),
.B(n_1439),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1498),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1409),
.B(n_1422),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1495),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1516),
.B(n_1518),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1473),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1439),
.B(n_1476),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1495),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1473),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1406),
.A2(n_1505),
.B1(n_1507),
.B2(n_1513),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1436),
.B(n_1514),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1444),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1515),
.B(n_1522),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1501),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1406),
.A2(n_1505),
.B(n_1507),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_SL g1581 ( 
.A(n_1503),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1407),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1489),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1408),
.Y(n_1584)
);

AOI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1475),
.A2(n_1490),
.B(n_1501),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1447),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1528),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1454),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1419),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1425),
.B(n_1521),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1454),
.Y(n_1591)
);

AO31x2_ASAP7_75t_L g1592 ( 
.A1(n_1457),
.A2(n_1529),
.A3(n_1500),
.B(n_1478),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1485),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1453),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1456),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1470),
.A2(n_1471),
.B(n_1499),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1417),
.B(n_1426),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1472),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1426),
.A2(n_1421),
.B(n_1487),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1462),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1467),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1483),
.A2(n_1494),
.B(n_1482),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1513),
.A2(n_1538),
.B1(n_1416),
.B2(n_1537),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1508),
.A2(n_1534),
.B1(n_1519),
.B2(n_1538),
.C(n_1504),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1450),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1511),
.B(n_1424),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1432),
.Y(n_1608)
);

AOI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1466),
.A2(n_1437),
.B(n_1442),
.Y(n_1609)
);

CKINVDCx6p67_ASAP7_75t_R g1610 ( 
.A(n_1405),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1412),
.A2(n_1431),
.B(n_1527),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1463),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1535),
.A2(n_1414),
.B1(n_1413),
.B2(n_1530),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1463),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1459),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1460),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1420),
.B(n_1411),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1459),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1459),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1451),
.A2(n_1434),
.B(n_1465),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1432),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1420),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1423),
.Y(n_1625)
);

AOI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1509),
.A2(n_1524),
.B(n_1415),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1403),
.B(n_1526),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1449),
.A2(n_1423),
.B(n_1433),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1531),
.A2(n_1433),
.B(n_1410),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1433),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1536),
.A2(n_1429),
.B1(n_1418),
.B2(n_1517),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1531),
.A2(n_1410),
.B(n_1523),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1517),
.B(n_1523),
.Y(n_1633)
);

INVx5_ASAP7_75t_L g1634 ( 
.A(n_1517),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1446),
.B(n_1404),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1405),
.B(n_1506),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1405),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1427),
.A2(n_1520),
.B(n_1532),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1430),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1447),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1580),
.A2(n_1546),
.B(n_1575),
.C(n_1604),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1605),
.A2(n_1548),
.B(n_1564),
.C(n_1598),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_R g1643 ( 
.A(n_1603),
.B(n_1616),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1558),
.B(n_1583),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1558),
.B(n_1583),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1557),
.A2(n_1585),
.B(n_1597),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1547),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1561),
.A2(n_1563),
.B(n_1550),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1578),
.A2(n_1589),
.B1(n_1576),
.B2(n_1596),
.C(n_1560),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1632),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1598),
.A2(n_1600),
.B(n_1560),
.C(n_1595),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1607),
.B(n_1572),
.Y(n_1654)
);

AOI211xp5_ASAP7_75t_L g1655 ( 
.A1(n_1602),
.A2(n_1600),
.B(n_1567),
.C(n_1606),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1561),
.A2(n_1563),
.B(n_1597),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1577),
.B(n_1574),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1577),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1595),
.A2(n_1566),
.B(n_1594),
.C(n_1588),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1562),
.B(n_1587),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1591),
.A2(n_1566),
.B1(n_1590),
.B2(n_1573),
.C(n_1569),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1541),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1609),
.A2(n_1603),
.B(n_1602),
.C(n_1611),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1547),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1590),
.A2(n_1569),
.B1(n_1573),
.B2(n_1579),
.C(n_1608),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1541),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1555),
.B(n_1565),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1611),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1603),
.A2(n_1601),
.B1(n_1561),
.B2(n_1611),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1579),
.A2(n_1568),
.B1(n_1570),
.B2(n_1594),
.C(n_1631),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1603),
.A2(n_1581),
.B1(n_1601),
.B2(n_1613),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1543),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1570),
.B(n_1611),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1593),
.B(n_1601),
.C(n_1584),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1552),
.A2(n_1542),
.B(n_1571),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1601),
.A2(n_1613),
.B1(n_1615),
.B2(n_1626),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1544),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1601),
.A2(n_1616),
.B1(n_1640),
.B2(n_1586),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1616),
.A2(n_1622),
.B(n_1629),
.C(n_1617),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1639),
.A2(n_1623),
.B1(n_1627),
.B2(n_1619),
.C(n_1633),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1623),
.A2(n_1620),
.B1(n_1619),
.B2(n_1640),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1617),
.A2(n_1592),
.B(n_1621),
.C(n_1634),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1563),
.A2(n_1628),
.B(n_1542),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_SL g1687 ( 
.A1(n_1621),
.A2(n_1637),
.B(n_1618),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1658),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1667),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1674),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1685),
.B(n_1563),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1669),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1679),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1641),
.A2(n_1586),
.B(n_1635),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1654),
.B(n_1549),
.Y(n_1696)
);

OR2x6_ASAP7_75t_SL g1697 ( 
.A(n_1678),
.B(n_1636),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1650),
.A2(n_1635),
.B1(n_1610),
.B2(n_1637),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1663),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1559),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1652),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1648),
.B(n_1559),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1641),
.A2(n_1610),
.B1(n_1614),
.B2(n_1612),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1687),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1661),
.B(n_1649),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1664),
.A2(n_1638),
.B1(n_1574),
.B2(n_1599),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1668),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1642),
.B(n_1680),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1684),
.B(n_1574),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1684),
.B(n_1559),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1657),
.B(n_1556),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1642),
.A2(n_1638),
.B1(n_1599),
.B2(n_1624),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1714),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1691),
.B(n_1656),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1699),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1688),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1702),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1711),
.Y(n_1721)
);

AO21x2_ASAP7_75t_L g1722 ( 
.A1(n_1702),
.A2(n_1646),
.B(n_1686),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1699),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1711),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1675),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1694),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1704),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1704),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1715),
.B(n_1692),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1689),
.Y(n_1730)
);

AND2x2_ASAP7_75t_SL g1731 ( 
.A(n_1710),
.B(n_1662),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1692),
.B(n_1670),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1710),
.B(n_1670),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1709),
.B(n_1682),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1694),
.Y(n_1735)
);

NOR2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1705),
.B(n_1647),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1705),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1666),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1693),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1694),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1695),
.B(n_1683),
.Y(n_1741)
);

INVx5_ASAP7_75t_L g1742 ( 
.A(n_1694),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1695),
.A2(n_1644),
.B1(n_1645),
.B2(n_1671),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1713),
.A2(n_1660),
.B(n_1655),
.C(n_1653),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1734),
.A2(n_1713),
.B1(n_1703),
.B2(n_1698),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1721),
.B(n_1690),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1718),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1721),
.B(n_1696),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1718),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1718),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1721),
.B(n_1696),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1723),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1738),
.B(n_1708),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1724),
.B(n_1706),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1742),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1723),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1716),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1706),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1730),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1716),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1701),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1744),
.B(n_1707),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1725),
.B(n_1672),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1742),
.B(n_1726),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1723),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1727),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1730),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1742),
.B(n_1694),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1733),
.B(n_1701),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1734),
.B(n_1697),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1727),
.Y(n_1772)
);

NOR2x1_ASAP7_75t_SL g1773 ( 
.A(n_1742),
.B(n_1694),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1727),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1742),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1725),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1741),
.B(n_1697),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1717),
.B(n_1693),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1728),
.Y(n_1781)
);

INVx3_ASAP7_75t_SL g1782 ( 
.A(n_1762),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1747),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1747),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1771),
.B(n_1731),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1749),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_1731),
.Y(n_1788)
);

AND2x4_ASAP7_75t_SL g1789 ( 
.A(n_1754),
.B(n_1712),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1750),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1750),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1770),
.B(n_1733),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1753),
.B(n_1720),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1754),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1770),
.B(n_1732),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1776),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_L g1797 ( 
.A(n_1776),
.B(n_1725),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1752),
.Y(n_1798)
);

INVx2_ASAP7_75t_SL g1799 ( 
.A(n_1765),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1761),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1753),
.B(n_1720),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1731),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1752),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1770),
.B(n_1732),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1776),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1761),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1773),
.B(n_1736),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1756),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1761),
.B(n_1732),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1777),
.B(n_1731),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1756),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1766),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1778),
.B(n_1731),
.Y(n_1814)
);

INVx2_ASAP7_75t_SL g1815 ( 
.A(n_1765),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1746),
.B(n_1732),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1746),
.B(n_1737),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1778),
.B(n_1720),
.Y(n_1819)
);

NOR2x1p5_ASAP7_75t_SL g1820 ( 
.A(n_1757),
.B(n_1760),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1767),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1767),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1772),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1755),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1780),
.B(n_1741),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1780),
.B(n_1729),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1782),
.B(n_1780),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1807),
.B(n_1754),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1782),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1796),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1794),
.B(n_1779),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1787),
.Y(n_1833)
);

NAND4xp75_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1762),
.C(n_1775),
.D(n_1763),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1787),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1810),
.B(n_1748),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1786),
.A2(n_1763),
.B(n_1745),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1807),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1807),
.B(n_1758),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1796),
.Y(n_1840)
);

INVxp67_ASAP7_75t_SL g1841 ( 
.A(n_1797),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1792),
.B(n_1758),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1817),
.B(n_1759),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1788),
.A2(n_1745),
.B(n_1744),
.C(n_1743),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1790),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1792),
.B(n_1758),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1825),
.B(n_1748),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1805),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1814),
.B(n_1743),
.C(n_1707),
.Y(n_1850)
);

AND2x4_ASAP7_75t_SL g1851 ( 
.A(n_1818),
.B(n_1765),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1795),
.B(n_1765),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1795),
.B(n_1748),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1804),
.B(n_1751),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1804),
.B(n_1759),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1819),
.B(n_1647),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1793),
.B(n_1779),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1818),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1751),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1790),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1827),
.B(n_1665),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1791),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1800),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1800),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1799),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1830),
.B(n_1665),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1840),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1849),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1830),
.B(n_1816),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1837),
.A2(n_1809),
.B1(n_1816),
.B2(n_1773),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1833),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1833),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1845),
.B(n_1789),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1835),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1865),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1865),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1851),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1828),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1835),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1846),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_L g1881 ( 
.A(n_1829),
.B(n_1799),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1834),
.A2(n_1703),
.B1(n_1736),
.B2(n_1643),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1855),
.B(n_1859),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1851),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1837),
.B(n_1806),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1806),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1834),
.A2(n_1736),
.B1(n_1643),
.B2(n_1789),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1851),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1836),
.B(n_1793),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1861),
.B(n_1751),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1846),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1850),
.A2(n_1698),
.B1(n_1722),
.B2(n_1801),
.Y(n_1892)
);

XNOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1878),
.B(n_1869),
.Y(n_1893)
);

AOI21xp33_ASAP7_75t_L g1894 ( 
.A1(n_1885),
.A2(n_1841),
.B(n_1850),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1869),
.B(n_1856),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1875),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1892),
.A2(n_1844),
.B1(n_1842),
.B2(n_1831),
.C(n_1855),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1866),
.B(n_1843),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1866),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1875),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1883),
.B(n_1848),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1876),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1892),
.A2(n_1838),
.B1(n_1844),
.B2(n_1854),
.C(n_1853),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1884),
.B(n_1829),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1877),
.B(n_1831),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1876),
.Y(n_1906)
);

XOR2x2_ASAP7_75t_L g1907 ( 
.A(n_1873),
.B(n_1839),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1877),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1871),
.Y(n_1909)
);

AOI222xp33_ASAP7_75t_L g1910 ( 
.A1(n_1873),
.A2(n_1831),
.B1(n_1842),
.B2(n_1820),
.C1(n_1860),
.C2(n_1862),
.Y(n_1910)
);

AOI31xp33_ASAP7_75t_L g1911 ( 
.A1(n_1870),
.A2(n_1842),
.A3(n_1680),
.B(n_1839),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1872),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1867),
.B(n_1843),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1899),
.B(n_1868),
.Y(n_1914)
);

OAI211xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1894),
.A2(n_1887),
.B(n_1888),
.C(n_1883),
.Y(n_1915)
);

AOI21xp33_ASAP7_75t_L g1916 ( 
.A1(n_1910),
.A2(n_1838),
.B(n_1877),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1903),
.A2(n_1882),
.B1(n_1881),
.B2(n_1838),
.Y(n_1917)
);

AOI21xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1893),
.A2(n_1838),
.B(n_1886),
.Y(n_1918)
);

OAI21xp33_ASAP7_75t_L g1919 ( 
.A1(n_1894),
.A2(n_1890),
.B(n_1889),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1904),
.B(n_1847),
.Y(n_1920)
);

NOR2x1_ASAP7_75t_SL g1921 ( 
.A(n_1908),
.B(n_1838),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1910),
.A2(n_1847),
.B1(n_1852),
.B2(n_1769),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1898),
.B(n_1874),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1911),
.A2(n_1880),
.B(n_1879),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1911),
.A2(n_1891),
.B(n_1864),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1924),
.B(n_1896),
.Y(n_1926)
);

NOR3xp33_ASAP7_75t_L g1927 ( 
.A(n_1915),
.B(n_1918),
.C(n_1914),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1925),
.B(n_1900),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1919),
.B(n_1902),
.Y(n_1929)
);

AND4x1_ASAP7_75t_L g1930 ( 
.A(n_1917),
.B(n_1906),
.C(n_1897),
.D(n_1922),
.Y(n_1930)
);

NAND4xp25_ASAP7_75t_L g1931 ( 
.A(n_1916),
.B(n_1895),
.C(n_1913),
.D(n_1901),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1923),
.B(n_1912),
.C(n_1909),
.Y(n_1932)
);

OR3x1_ASAP7_75t_L g1933 ( 
.A(n_1921),
.B(n_1907),
.C(n_1862),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1920),
.Y(n_1934)
);

NAND4xp25_ASAP7_75t_L g1935 ( 
.A(n_1917),
.B(n_1852),
.C(n_1864),
.D(n_1863),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1915),
.B(n_1864),
.C(n_1863),
.Y(n_1936)
);

OAI21xp33_ASAP7_75t_L g1937 ( 
.A1(n_1931),
.A2(n_1905),
.B(n_1863),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1927),
.A2(n_1905),
.B1(n_1755),
.B2(n_1775),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1933),
.A2(n_1860),
.B1(n_1824),
.B2(n_1815),
.C(n_1857),
.Y(n_1939)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1940 ( 
.A1(n_1926),
.A2(n_1791),
.B(n_1798),
.C(n_1826),
.D(n_1803),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1929),
.B(n_1815),
.C(n_1824),
.Y(n_1941)
);

O2A1O1Ixp5_ASAP7_75t_SL g1942 ( 
.A1(n_1928),
.A2(n_1798),
.B(n_1803),
.C(n_1826),
.Y(n_1942)
);

NAND4xp75_ASAP7_75t_L g1943 ( 
.A(n_1934),
.B(n_1820),
.C(n_1775),
.D(n_1726),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1938),
.A2(n_1930),
.B(n_1935),
.Y(n_1944)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1945 ( 
.A1(n_1937),
.A2(n_1936),
.B(n_1932),
.C(n_1821),
.D(n_1822),
.Y(n_1945)
);

OAI211xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1939),
.A2(n_1941),
.B(n_1940),
.C(n_1942),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1943),
.A2(n_1755),
.B1(n_1769),
.B2(n_1765),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_SL g1948 ( 
.A(n_1938),
.B(n_1832),
.C(n_1857),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1937),
.A2(n_1801),
.B(n_1832),
.Y(n_1949)
);

NOR2x1_ASAP7_75t_L g1950 ( 
.A(n_1937),
.B(n_1755),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1937),
.A2(n_1755),
.B1(n_1822),
.B2(n_1821),
.C(n_1823),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1950),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1948),
.A2(n_1769),
.B1(n_1737),
.B2(n_1823),
.Y(n_1953)
);

NOR2x1_ASAP7_75t_L g1954 ( 
.A(n_1946),
.B(n_1783),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1945),
.Y(n_1955)
);

INVxp33_ASAP7_75t_L g1956 ( 
.A(n_1944),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1949),
.Y(n_1957)
);

NOR2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1957),
.B(n_1951),
.Y(n_1958)
);

XNOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1956),
.B(n_1947),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1954),
.A2(n_1785),
.B(n_1784),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1955),
.A2(n_1737),
.B1(n_1812),
.B2(n_1811),
.C(n_1808),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1959),
.A2(n_1952),
.B(n_1953),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1958),
.B1(n_1961),
.B2(n_1960),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1963),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1963),
.Y(n_1965)
);

AOI22x1_ASAP7_75t_L g1966 ( 
.A1(n_1964),
.A2(n_1965),
.B1(n_1813),
.B2(n_1768),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1964),
.B(n_1769),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1967),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1966),
.A2(n_1768),
.B(n_1769),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1968),
.A2(n_1719),
.B1(n_1739),
.B2(n_1781),
.C(n_1774),
.Y(n_1970)
);

AO21x2_ASAP7_75t_L g1971 ( 
.A1(n_1970),
.A2(n_1969),
.B(n_1764),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1971),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1726),
.B1(n_1740),
.B2(n_1735),
.Y(n_1973)
);

AOI211xp5_ASAP7_75t_L g1974 ( 
.A1(n_1973),
.A2(n_1681),
.B(n_1630),
.C(n_1625),
.Y(n_1974)
);


endmodule