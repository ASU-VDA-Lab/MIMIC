module fake_aes_2060_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_0), .B(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_1), .B(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_7), .B(n_4), .Y(n_8) );
OAI21xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_4), .B(n_5), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_6), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_8), .B(n_5), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_11), .B(n_9), .Y(n_12) );
NAND3xp33_ASAP7_75t_SL g13 ( .A(n_10), .B(n_9), .C(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AOI221xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_1), .B1(n_2), .B2(n_10), .C(n_12), .Y(n_15) );
XOR2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_2), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_16), .B(n_15), .Y(n_17) );
endmodule