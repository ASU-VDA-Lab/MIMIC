module fake_jpeg_3534_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

AND2x6_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_3),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_24)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_21),
.B(n_23),
.Y(n_28)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_0),
.C(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx12_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_21),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_23),
.CON(n_31),
.SN(n_31)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_29),
.B(n_16),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_16),
.B(n_17),
.C(n_13),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_26),
.C(n_27),
.Y(n_35)
);

OAI21x1_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_35),
.B(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_32),
.C(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_11),
.A3(n_7),
.B1(n_13),
.B2(n_22),
.C1(n_20),
.C2(n_14),
.Y(n_41)
);

AOI211xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B(n_14),
.C(n_20),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_7),
.B(n_18),
.Y(n_42)
);


endmodule