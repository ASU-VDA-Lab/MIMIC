module real_aes_13399_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_905;
wire n_357;
wire n_386;
wire n_287;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OA21x2_ASAP7_75t_L g154 ( .A1(n_0), .A2(n_51), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g290 ( .A(n_0), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_1), .A2(n_901), .B1(n_907), .B2(n_908), .Y(n_900) );
INVx1_ASAP7_75t_L g907 ( .A(n_1), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_2), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g214 ( .A(n_3), .B(n_206), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_4), .B(n_204), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_5), .A2(n_99), .B1(n_238), .B2(n_264), .C(n_286), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_6), .B(n_191), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_7), .B(n_555), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_8), .B(n_159), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_9), .B(n_195), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_10), .Y(n_548) );
BUFx3_ASAP7_75t_L g161 ( .A(n_11), .Y(n_161) );
INVx1_ASAP7_75t_L g172 ( .A(n_11), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_12), .B(n_174), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_13), .A2(n_207), .B(n_573), .C(n_574), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_14), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_15), .A2(n_142), .B1(n_535), .B2(n_536), .Y(n_141) );
INVx1_ASAP7_75t_L g536 ( .A(n_15), .Y(n_536) );
OAI22x1_ASAP7_75t_SL g903 ( .A1(n_15), .A2(n_101), .B1(n_536), .B2(n_904), .Y(n_903) );
BUFx10_ASAP7_75t_L g126 ( .A(n_16), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_17), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_18), .B(n_309), .Y(n_625) );
INVx1_ASAP7_75t_L g912 ( .A(n_19), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_20), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_21), .B(n_182), .Y(n_272) );
OAI21xp33_ASAP7_75t_L g385 ( .A1(n_21), .A2(n_68), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_22), .B(n_307), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_23), .A2(n_564), .B(n_565), .C(n_567), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_24), .B(n_614), .Y(n_664) );
O2A1O1Ixp5_ASAP7_75t_L g317 ( .A1(n_25), .A2(n_208), .B(n_243), .C(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g606 ( .A(n_26), .B(n_191), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_27), .B(n_182), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_28), .A2(n_78), .B1(n_159), .B2(n_163), .Y(n_557) );
INVx1_ASAP7_75t_L g180 ( .A(n_29), .Y(n_180) );
INVx1_ASAP7_75t_L g587 ( .A(n_30), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_31), .B(n_164), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_32), .B(n_163), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_33), .B(n_182), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_34), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g116 ( .A(n_35), .Y(n_116) );
AND3x2_ASAP7_75t_L g888 ( .A(n_35), .B(n_108), .C(n_123), .Y(n_888) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_36), .B(n_238), .Y(n_663) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_37), .A2(n_46), .B1(n_132), .B2(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_37), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_38), .B(n_182), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_39), .B(n_243), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_40), .B(n_174), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_41), .Y(n_575) );
AND2x4_ASAP7_75t_L g179 ( .A(n_42), .B(n_180), .Y(n_179) );
NAND2x1_ASAP7_75t_L g205 ( .A(n_43), .B(n_206), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_44), .Y(n_282) );
INVx1_ASAP7_75t_L g200 ( .A(n_45), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_46), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_47), .Y(n_301) );
AND2x2_ASAP7_75t_L g213 ( .A(n_48), .B(n_170), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_49), .B(n_163), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_50), .A2(n_92), .B1(n_163), .B2(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g291 ( .A(n_51), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_52), .B(n_191), .Y(n_311) );
INVx1_ASAP7_75t_L g155 ( .A(n_53), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_54), .B(n_170), .Y(n_220) );
AOI21xp33_ASAP7_75t_L g883 ( .A1(n_55), .A2(n_884), .B(n_889), .Y(n_883) );
AND2x4_ASAP7_75t_L g113 ( .A(n_56), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_57), .B(n_182), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_58), .B(n_204), .Y(n_203) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_59), .B(n_80), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_60), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g669 ( .A(n_61), .B(n_183), .Y(n_669) );
INVx1_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_63), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_64), .B(n_614), .Y(n_613) );
NAND2x1_ASAP7_75t_L g636 ( .A(n_65), .B(n_573), .Y(n_636) );
AND2x2_ASAP7_75t_L g218 ( .A(n_66), .B(n_191), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_67), .B(n_174), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_68), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_69), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_70), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_71), .B(n_163), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_72), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_73), .B(n_298), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_74), .B(n_624), .Y(n_623) );
AND3x2_ASAP7_75t_L g107 ( .A(n_75), .B(n_108), .C(n_110), .Y(n_107) );
INVx2_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_76), .B(n_235), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_77), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_79), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_81), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_82), .B(n_238), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_83), .B(n_183), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_84), .B(n_170), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_85), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_86), .B(n_309), .Y(n_633) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_87), .B(n_281), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_88), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_89), .B(n_170), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_90), .B(n_237), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_91), .B(n_259), .Y(n_258) );
AOI22x1_ASAP7_75t_L g901 ( .A1(n_93), .A2(n_902), .B1(n_905), .B2(n_906), .Y(n_901) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_93), .Y(n_906) );
INVx1_ASAP7_75t_L g167 ( .A(n_94), .Y(n_167) );
BUFx3_ASAP7_75t_L g177 ( .A(n_94), .Y(n_177) );
INVx1_ASAP7_75t_L g209 ( .A(n_94), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_95), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_96), .B(n_283), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_97), .A2(n_130), .B1(n_131), .B2(n_134), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_97), .Y(n_134) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_98), .B(n_201), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_100), .B(n_309), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_101), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_102), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_103), .B(n_170), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_117), .B(n_911), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_106), .Y(n_915) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g122 ( .A(n_108), .B(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_109), .B(n_116), .Y(n_895) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_896), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B(n_883), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx5_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g894 ( .A(n_124), .Y(n_894) );
BUFx3_ASAP7_75t_L g910 ( .A(n_125), .Y(n_910) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_126), .B(n_888), .Y(n_887) );
CKINVDCx11_ASAP7_75t_R g899 ( .A(n_126), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B1(n_135), .B2(n_136), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_537), .Y(n_136) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_138), .Y(n_538) );
CKINVDCx10_ASAP7_75t_R g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g535 ( .A(n_142), .Y(n_535) );
NOR2x1_ASAP7_75t_L g142 ( .A(n_143), .B(n_461), .Y(n_142) );
NAND4xp25_ASAP7_75t_L g143 ( .A(n_144), .B(n_369), .C(n_410), .D(n_443), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_344), .Y(n_144) );
OAI222xp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_249), .B1(n_312), .B2(n_327), .C1(n_332), .C2(n_339), .Y(n_145) );
NOR2xp67_ASAP7_75t_SL g146 ( .A(n_147), .B(n_227), .Y(n_146) );
AND2x2_ASAP7_75t_L g444 ( .A(n_147), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_185), .Y(n_147) );
AND2x2_ASAP7_75t_L g378 ( .A(n_148), .B(n_230), .Y(n_378) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_148), .Y(n_395) );
INVx1_ASAP7_75t_L g416 ( .A(n_148), .Y(n_416) );
INVx1_ASAP7_75t_L g465 ( .A(n_148), .Y(n_465) );
AND2x2_ASAP7_75t_L g505 ( .A(n_148), .B(n_436), .Y(n_505) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g247 ( .A(n_149), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g408 ( .A(n_149), .B(n_187), .Y(n_408) );
AND2x2_ASAP7_75t_L g479 ( .A(n_149), .B(n_331), .Y(n_479) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g366 ( .A(n_150), .Y(n_366) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_156), .B(n_181), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_152), .A2(n_178), .B(n_586), .Y(n_589) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g386 ( .A(n_153), .Y(n_386) );
BUFx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_154), .Y(n_191) );
INVxp33_ASAP7_75t_L g588 ( .A(n_154), .Y(n_588) );
INVx1_ASAP7_75t_L g292 ( .A(n_155), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_168), .B(n_178), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_162), .B(n_165), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g283 ( .A(n_160), .Y(n_283) );
INVx1_ASAP7_75t_L g298 ( .A(n_160), .Y(n_298) );
INVx2_ASAP7_75t_L g307 ( .A(n_160), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_160), .B(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g164 ( .A(n_161), .Y(n_164) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
INVx1_ASAP7_75t_L g235 ( .A(n_164), .Y(n_235) );
INVx2_ASAP7_75t_L g277 ( .A(n_164), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_165), .A2(n_234), .B(n_236), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_165), .A2(n_262), .B(n_265), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_165), .A2(n_305), .B(n_308), .Y(n_304) );
AO21x1_ASAP7_75t_L g578 ( .A1(n_165), .A2(n_579), .B(n_580), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_165), .A2(n_612), .B(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_165), .A2(n_623), .B(n_625), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_165), .A2(n_632), .B(n_633), .Y(n_631) );
BUFx10_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g286 ( .A(n_167), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_176), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
INVx2_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
INVx2_ASAP7_75t_L g281 ( .A(n_171), .Y(n_281) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
INVx3_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
INVx2_ASAP7_75t_L g555 ( .A(n_175), .Y(n_555) );
INVx2_ASAP7_75t_L g584 ( .A(n_175), .Y(n_584) );
INVx2_ASAP7_75t_L g614 ( .A(n_175), .Y(n_614) );
AO21x1_ASAP7_75t_L g581 ( .A1(n_176), .A2(n_582), .B(n_583), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_176), .A2(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g195 ( .A(n_177), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_177), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
AOI211x1_ASAP7_75t_L g607 ( .A1(n_177), .A2(n_606), .B(n_608), .C(n_611), .Y(n_607) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_178), .A2(n_193), .B(n_202), .Y(n_192) );
INVx1_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_178), .A2(n_593), .B(n_596), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_178), .A2(n_605), .B(n_606), .Y(n_604) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_178), .A2(n_619), .B(n_622), .Y(n_618) );
BUFx6f_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
INVx2_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
INVx1_ASAP7_75t_L g288 ( .A(n_179), .Y(n_288) );
INVx1_ASAP7_75t_L g552 ( .A(n_179), .Y(n_552) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_183), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g377 ( .A(n_185), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g396 ( .A(n_185), .B(n_365), .Y(n_396) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g469 ( .A(n_186), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_211), .Y(n_186) );
INVx2_ASAP7_75t_L g248 ( .A(n_187), .Y(n_248) );
AND2x4_ASAP7_75t_SL g343 ( .A(n_187), .B(n_246), .Y(n_343) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_187), .Y(n_354) );
INVx1_ASAP7_75t_L g368 ( .A(n_187), .Y(n_368) );
INVxp67_ASAP7_75t_L g437 ( .A(n_187), .Y(n_437) );
INVx1_ASAP7_75t_L g454 ( .A(n_187), .Y(n_454) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_192), .B(n_210), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVxp33_ASAP7_75t_L g224 ( .A(n_191), .Y(n_224) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_191), .Y(n_254) );
INVx1_ASAP7_75t_L g323 ( .A(n_191), .Y(n_323) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_191), .Y(n_605) );
NOR2xp67_ASAP7_75t_SL g661 ( .A(n_191), .B(n_288), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_198), .Y(n_193) );
INVx1_ASAP7_75t_L g567 ( .A(n_195), .Y(n_567) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
AOI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B(n_207), .Y(n_202) );
INVx1_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_207), .A2(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g260 ( .A(n_208), .Y(n_260) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx3_ASAP7_75t_L g216 ( .A(n_209), .Y(n_216) );
INVx2_ASAP7_75t_L g246 ( .A(n_211), .Y(n_246) );
INVx1_ASAP7_75t_L g331 ( .A(n_211), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_211), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g423 ( .A(n_211), .B(n_330), .Y(n_423) );
OR2x2_ASAP7_75t_L g458 ( .A(n_211), .B(n_230), .Y(n_458) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_217), .B(n_223), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g222 ( .A(n_216), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_216), .B(n_389), .C(n_551), .Y(n_556) );
O2A1O1Ixp5_ASAP7_75t_L g634 ( .A1(n_216), .A2(n_297), .B(n_635), .C(n_636), .Y(n_634) );
NOR2xp67_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AOI21xp33_ASAP7_75t_L g223 ( .A1(n_218), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_222), .A2(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g315 ( .A(n_226), .B(n_316), .C(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_247), .Y(n_228) );
AND2x2_ASAP7_75t_L g405 ( .A(n_229), .B(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g426 ( .A(n_229), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_229), .B(n_416), .Y(n_507) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_246), .Y(n_229) );
INVx3_ASAP7_75t_L g330 ( .A(n_230), .Y(n_330) );
INVx1_ASAP7_75t_L g341 ( .A(n_230), .Y(n_341) );
AND2x2_ASAP7_75t_L g436 ( .A(n_230), .B(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_230), .Y(n_442) );
INVx1_ASAP7_75t_L g503 ( .A(n_230), .Y(n_503) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_240), .B(n_244), .Y(n_232) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g564 ( .A(n_238), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_238), .B(n_575), .Y(n_574) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g264 ( .A(n_239), .Y(n_264) );
BUFx2_ASAP7_75t_L g394 ( .A(n_246), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_247), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g488 ( .A(n_247), .Y(n_488) );
AND2x2_ASAP7_75t_L g533 ( .A(n_247), .B(n_503), .Y(n_533) );
AND2x2_ASAP7_75t_L g476 ( .A(n_248), .B(n_366), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_250), .B(n_269), .Y(n_249) );
INVx2_ASAP7_75t_L g347 ( .A(n_250), .Y(n_347) );
AND2x2_ASAP7_75t_L g409 ( .A(n_250), .B(n_357), .Y(n_409) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g392 ( .A(n_251), .B(n_338), .Y(n_392) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g398 ( .A(n_252), .B(n_314), .Y(n_398) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_255), .B(n_268), .Y(n_252) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_253), .A2(n_295), .B(n_311), .Y(n_294) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_253), .A2(n_295), .B(n_311), .Y(n_336) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_253), .A2(n_255), .B(n_268), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_253), .A2(n_618), .B(n_626), .Y(n_617) );
OAI21x1_ASAP7_75t_L g629 ( .A1(n_253), .A2(n_630), .B(n_637), .Y(n_629) );
OAI21x1_ASAP7_75t_L g653 ( .A1(n_253), .A2(n_618), .B(n_626), .Y(n_653) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_261), .B(n_266), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g553 ( .A(n_260), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_263), .A2(n_609), .B(n_610), .Y(n_608) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_264), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g573 ( .A(n_264), .Y(n_573) );
INVx2_ASAP7_75t_L g624 ( .A(n_264), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_266), .A2(n_631), .B(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g310 ( .A(n_267), .Y(n_310) );
AND2x2_ASAP7_75t_L g455 ( .A(n_269), .B(n_398), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_269), .B(n_347), .Y(n_466) );
AND2x2_ASAP7_75t_L g471 ( .A(n_269), .B(n_365), .Y(n_471) );
AND2x2_ASAP7_75t_L g485 ( .A(n_269), .B(n_392), .Y(n_485) );
AND2x2_ASAP7_75t_L g515 ( .A(n_269), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_293), .Y(n_269) );
INVx1_ASAP7_75t_L g499 ( .A(n_270), .Y(n_499) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g326 ( .A(n_271), .Y(n_326) );
INVx2_ASAP7_75t_L g349 ( .A(n_271), .Y(n_349) );
AND2x2_ASAP7_75t_L g357 ( .A(n_271), .B(n_294), .Y(n_357) );
AND2x2_ASAP7_75t_L g497 ( .A(n_271), .B(n_335), .Y(n_497) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_273), .B(n_385), .C(n_387), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_280), .C(n_287), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_278), .C(n_279), .Y(n_274) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_279), .A2(n_594), .B(n_595), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_279), .A2(n_667), .B(n_668), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_283), .B2(n_284), .C(n_285), .Y(n_280) );
INVx2_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_286), .A2(n_297), .B1(n_299), .B2(n_303), .Y(n_296) );
INVx2_ASAP7_75t_SL g302 ( .A(n_286), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g389 ( .A(n_289), .Y(n_389) );
AOI21x1_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_289) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_290), .A2(n_291), .B(n_292), .Y(n_320) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g348 ( .A(n_294), .B(n_349), .Y(n_348) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_304), .B(n_310), .Y(n_295) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_310), .B(n_320), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_324), .Y(n_312) );
AND2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_334), .Y(n_350) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g338 ( .A(n_314), .Y(n_338) );
AND2x2_ASAP7_75t_L g359 ( .A(n_314), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g473 ( .A(n_314), .Y(n_473) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_320), .B(n_321), .Y(n_314) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_315), .B(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_320), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g570 ( .A(n_320), .Y(n_570) );
NOR2xp33_ASAP7_75t_R g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_325), .Y(n_412) );
AND2x2_ASAP7_75t_L g486 ( .A(n_325), .B(n_359), .Y(n_486) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_326), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g351 ( .A(n_328), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
AND2x2_ASAP7_75t_L g358 ( .A(n_333), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g391 ( .A(n_334), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g494 ( .A(n_334), .Y(n_494) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
AND2x4_ASAP7_75t_L g516 ( .A(n_338), .B(n_432), .Y(n_516) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g445 ( .A(n_340), .Y(n_445) );
AOI32xp33_ASAP7_75t_L g470 ( .A1(n_340), .A2(n_471), .A3(n_472), .B1(n_474), .B2(n_475), .Y(n_470) );
AND2x4_ASAP7_75t_L g512 ( .A(n_340), .B(n_469), .Y(n_512) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g453 ( .A(n_341), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g419 ( .A(n_342), .Y(n_419) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g372 ( .A(n_343), .B(n_365), .Y(n_372) );
AND2x2_ASAP7_75t_L g403 ( .A(n_343), .B(n_364), .Y(n_403) );
AND2x2_ASAP7_75t_L g441 ( .A(n_343), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_355), .Y(n_344) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_350), .B(n_351), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g356 ( .A(n_347), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g528 ( .A(n_347), .B(n_460), .Y(n_528) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_398), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_348), .A2(n_378), .B1(n_405), .B2(n_409), .Y(n_404) );
AND2x2_ASAP7_75t_L g474 ( .A(n_348), .B(n_359), .Y(n_474) );
AND2x2_ASAP7_75t_L g482 ( .A(n_348), .B(n_392), .Y(n_482) );
AND2x4_ASAP7_75t_SL g534 ( .A(n_348), .B(n_516), .Y(n_534) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g422 ( .A(n_354), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_362), .Y(n_355) );
AND2x2_ASAP7_75t_L g428 ( .A(n_357), .B(n_398), .Y(n_428) );
INVx1_ASAP7_75t_L g446 ( .A(n_357), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_359), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g432 ( .A(n_360), .Y(n_432) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g530 ( .A(n_365), .B(n_423), .Y(n_530) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g464 ( .A(n_367), .B(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_399), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B1(n_376), .B2(n_379), .C(n_390), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g397 ( .A(n_374), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
OR2x2_ASAP7_75t_L g460 ( .A(n_375), .B(n_384), .Y(n_460) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g447 ( .A(n_381), .Y(n_447) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g439 ( .A(n_382), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g433 ( .A(n_384), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g440 ( .A(n_384), .Y(n_440) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_386), .A2(n_592), .B(n_599), .Y(n_591) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_389), .B(n_551), .C(n_553), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_396), .B2(n_397), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_391), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
AND2x2_ASAP7_75t_L g475 ( .A(n_394), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g451 ( .A(n_395), .Y(n_451) );
AND2x2_ASAP7_75t_L g498 ( .A(n_398), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_398), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g525 ( .A(n_398), .B(n_497), .Y(n_525) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_402), .B(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_403), .B(n_445), .Y(n_492) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g502 ( .A(n_408), .B(n_503), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_424), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .C(n_420), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g456 ( .A(n_415), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B1(n_429), .B2(n_435), .C(n_438), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_430), .B(n_468), .Y(n_467) );
NOR2x1p5_ASAP7_75t_SL g430 ( .A(n_431), .B(n_433), .Y(n_430) );
AND2x2_ASAP7_75t_L g496 ( .A(n_431), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_431), .B(n_471), .Y(n_510) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_439), .A2(n_518), .B(n_521), .Y(n_517) );
AOI322xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .A3(n_447), .B1(n_448), .B2(n_455), .C1(n_456), .C2(n_459), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g480 ( .A(n_452), .Y(n_480) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g484 ( .A(n_458), .Y(n_484) );
INVx1_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
INVx2_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_458), .B(n_476), .Y(n_527) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_460), .B(n_507), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_490), .C(n_508), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .Y(n_462) );
OAI211xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B(n_467), .C(n_470), .Y(n_463) );
INVx2_ASAP7_75t_L g532 ( .A(n_464), .Y(n_532) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI221x1_ASAP7_75t_L g495 ( .A1(n_475), .A2(n_496), .B1(n_498), .B2(n_500), .C(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g521 ( .A(n_476), .B(n_522), .Y(n_521) );
OAI21xp33_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_481), .B(n_483), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_486), .B(n_494), .Y(n_493) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B(n_495), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI21xp33_ASAP7_75t_SL g509 ( .A1(n_493), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g520 ( .A(n_499), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_502), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR3xp33_ASAP7_75t_SL g508 ( .A(n_509), .B(n_513), .C(n_523), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_528), .B2(n_529), .C(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
XNOR2xp5_ASAP7_75t_L g902 ( .A(n_535), .B(n_903), .Y(n_902) );
XOR2xp5_ASAP7_75t_L g905 ( .A(n_535), .B(n_903), .Y(n_905) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_787), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_696), .C(n_760), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_600), .B1(n_638), .B2(n_649), .C(n_654), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_558), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g708 ( .A(n_545), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g723 ( .A(n_545), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g796 ( .A(n_545), .B(n_576), .Y(n_796) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g646 ( .A(n_546), .Y(n_646) );
INVx1_ASAP7_75t_L g675 ( .A(n_546), .Y(n_675) );
AND2x2_ASAP7_75t_L g694 ( .A(n_546), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g721 ( .A(n_546), .B(n_711), .Y(n_721) );
INVxp67_ASAP7_75t_L g736 ( .A(n_546), .Y(n_736) );
AND2x2_ASAP7_75t_L g759 ( .A(n_546), .B(n_591), .Y(n_759) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_546), .Y(n_786) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B1(n_556), .B2(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_558), .A2(n_765), .B(n_769), .Y(n_764) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_576), .Y(n_558) );
AND2x2_ASAP7_75t_L g866 ( .A(n_559), .B(n_759), .Y(n_866) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g642 ( .A(n_561), .Y(n_642) );
INVx1_ASAP7_75t_L g677 ( .A(n_561), .Y(n_677) );
AND2x2_ASAP7_75t_L g705 ( .A(n_561), .B(n_645), .Y(n_705) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_561), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_562), .B(n_571), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_562), .B(n_571), .Y(n_695) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .B(n_569), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_567), .A2(n_597), .B(n_598), .Y(n_596) );
OR2x2_ASAP7_75t_L g571 ( .A(n_568), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g693 ( .A(n_576), .B(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g882 ( .A(n_576), .Y(n_882) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_590), .Y(n_576) );
INVx2_ASAP7_75t_L g645 ( .A(n_577), .Y(n_645) );
AND2x2_ASAP7_75t_L g676 ( .A(n_577), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g687 ( .A(n_577), .Y(n_687) );
OR2x2_ASAP7_75t_L g725 ( .A(n_577), .B(n_695), .Y(n_725) );
AND2x2_ASAP7_75t_L g737 ( .A(n_577), .B(n_695), .Y(n_737) );
AND2x2_ASAP7_75t_L g807 ( .A(n_577), .B(n_591), .Y(n_807) );
AO31x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .A3(n_585), .B(n_589), .Y(n_577) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
INVx1_ASAP7_75t_L g711 ( .A(n_591), .Y(n_711) );
AND2x2_ASAP7_75t_L g733 ( .A(n_591), .B(n_646), .Y(n_733) );
AND2x2_ASAP7_75t_L g816 ( .A(n_591), .B(n_710), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_615), .Y(n_600) );
AND2x2_ASAP7_75t_L g739 ( .A(n_601), .B(n_730), .Y(n_739) );
OR2x2_ASAP7_75t_L g755 ( .A(n_601), .B(n_690), .Y(n_755) );
INVx2_ASAP7_75t_L g767 ( .A(n_601), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_601), .B(n_703), .Y(n_770) );
AND2x2_ASAP7_75t_L g867 ( .A(n_601), .B(n_782), .Y(n_867) );
BUFx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g650 ( .A(n_602), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g777 ( .A(n_602), .B(n_682), .Y(n_777) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g670 ( .A(n_603), .B(n_617), .Y(n_670) );
INVx2_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
BUFx2_ASAP7_75t_L g728 ( .A(n_603), .Y(n_728) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_603), .Y(n_745) );
INVx1_ASAP7_75t_L g752 ( .A(n_603), .Y(n_752) );
AND2x2_ASAP7_75t_L g811 ( .A(n_603), .B(n_754), .Y(n_811) );
INVx1_ASAP7_75t_L g872 ( .A(n_603), .Y(n_872) );
OR2x6_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_627), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_616), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g681 ( .A(n_617), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g837 ( .A(n_627), .Y(n_837) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g754 ( .A(n_628), .Y(n_754) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g680 ( .A(n_629), .Y(n_680) );
INVx1_ASAP7_75t_L g717 ( .A(n_629), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_638), .A2(n_761), .B(n_764), .C(n_771), .Y(n_760) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_642), .Y(n_684) );
AND2x2_ASAP7_75t_L g803 ( .A(n_642), .B(n_733), .Y(n_803) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
AND2x2_ASAP7_75t_L g713 ( .A(n_644), .B(n_709), .Y(n_713) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g774 ( .A(n_645), .Y(n_774) );
INVx2_ASAP7_75t_L g747 ( .A(n_647), .Y(n_747) );
BUFx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_648), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_648), .Y(n_849) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g703 ( .A(n_651), .B(n_680), .Y(n_703) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g716 ( .A(n_652), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g730 ( .A(n_652), .B(n_659), .Y(n_730) );
AND2x2_ASAP7_75t_L g853 ( .A(n_652), .B(n_680), .Y(n_853) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g691 ( .A(n_653), .B(n_659), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_671), .B1(n_678), .B2(n_683), .C(n_688), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_655), .A2(n_783), .B1(n_846), .B2(n_851), .C1(n_854), .C2(n_855), .Y(n_845) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_670), .Y(n_656) );
INVx4_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_658), .B(n_746), .Y(n_763) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g682 ( .A(n_659), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_659), .B(n_680), .Y(n_690) );
AND2x4_ASAP7_75t_L g751 ( .A(n_659), .B(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_665), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_661), .A2(n_666), .B(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g706 ( .A(n_670), .Y(n_706) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_676), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_673), .B(n_859), .C(n_862), .Y(n_858) );
OR2x2_ASAP7_75t_L g874 ( .A(n_673), .B(n_862), .Y(n_874) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_674), .A2(n_744), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g808 ( .A(n_675), .B(n_695), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_676), .B(n_759), .Y(n_779) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
OR2x2_ASAP7_75t_L g822 ( .A(n_679), .B(n_691), .Y(n_822) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g800 ( .A(n_681), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_681), .B(n_727), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_681), .B(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_681), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_681), .B(n_837), .Y(n_865) );
AND2x4_ASAP7_75t_SL g700 ( .A(n_682), .B(n_701), .Y(n_700) );
NOR2x1p5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
BUFx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g758 ( .A(n_687), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_687), .B(n_849), .Y(n_848) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx4_ASAP7_75t_L g782 ( .A(n_691), .Y(n_782) );
NOR2x1_ASAP7_75t_L g879 ( .A(n_691), .B(n_871), .Y(n_879) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g814 ( .A(n_694), .B(n_807), .Y(n_814) );
INVx2_ASAP7_75t_L g710 ( .A(n_695), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_740), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_718), .C(n_731), .Y(n_697) );
OAI322xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .A3(n_704), .B1(n_706), .B2(n_707), .C1(n_712), .C2(n_714), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g838 ( .A(n_700), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_702), .A2(n_813), .B1(n_815), .B2(n_817), .Y(n_812) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_703), .B(n_751), .Y(n_856) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_SL g720 ( .A(n_705), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g801 ( .A(n_705), .B(n_759), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_705), .B(n_736), .Y(n_877) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g833 ( .A(n_708), .B(n_774), .Y(n_833) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI322xp5_ASAP7_75t_L g771 ( .A1(n_714), .A2(n_751), .A3(n_772), .B1(n_775), .B2(n_778), .C1(n_780), .C2(n_783), .Y(n_771) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp33_ASAP7_75t_L g776 ( .A(n_715), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g768 ( .A(n_716), .Y(n_768) );
OR2x2_ASAP7_75t_L g791 ( .A(n_716), .B(n_777), .Y(n_791) );
BUFx2_ASAP7_75t_L g746 ( .A(n_717), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B(n_726), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_719), .A2(n_749), .B1(n_755), .B2(n_756), .Y(n_748) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g841 ( .A(n_721), .Y(n_841) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g744 ( .A(n_725), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g784 ( .A(n_725), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g824 ( .A(n_725), .B(n_825), .Y(n_824) );
OR2x2_ASAP7_75t_L g840 ( .A(n_725), .B(n_841), .Y(n_840) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_728), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g799 ( .A(n_728), .Y(n_799) );
OR2x2_ASAP7_75t_L g817 ( .A(n_729), .B(n_753), .Y(n_817) );
OR2x2_ASAP7_75t_L g843 ( .A(n_729), .B(n_837), .Y(n_843) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B(n_738), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_733), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g862 ( .A(n_737), .Y(n_862) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_747), .B(n_748), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_746), .Y(n_742) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_751), .B(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_752), .Y(n_828) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g871 ( .A(n_754), .B(n_872), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_756), .B(n_840), .Y(n_839) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g794 ( .A(n_758), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_759), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g825 ( .A(n_759), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_761), .B(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g844 ( .A(n_767), .Y(n_844) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_767), .B(n_782), .C(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVxp67_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g881 ( .A(n_785), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR3xp33_ASAP7_75t_SL g787 ( .A(n_788), .B(n_829), .C(n_857), .Y(n_787) );
NAND3xp33_ASAP7_75t_SL g788 ( .A(n_789), .B(n_802), .C(n_818), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_792), .B1(n_797), .B2(n_801), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_795), .Y(n_792) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_796), .A2(n_864), .B1(n_866), .B2(n_867), .Y(n_863) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OR2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_804), .B1(n_806), .B2(n_809), .C(n_812), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g820 ( .A(n_806), .Y(n_820) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx2_ASAP7_75t_L g850 ( .A(n_808), .Y(n_850) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVxp33_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g878 ( .A(n_817), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_821), .B1(n_823), .B2(n_826), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI211xp5_ASAP7_75t_SL g829 ( .A1(n_830), .A2(n_832), .B(n_834), .C(n_845), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_833), .A2(n_835), .B1(n_839), .B2(n_842), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g861 ( .A(n_837), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_843), .B(n_844), .Y(n_842) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
INVxp67_ASAP7_75t_SL g854 ( .A(n_848), .Y(n_854) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVxp67_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_858), .B(n_863), .C(n_868), .D(n_875), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_873), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
BUFx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
BUFx3_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_889), .B(n_910), .Y(n_909) );
NOR2x1_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AND2x4_ASAP7_75t_L g898 ( .A(n_892), .B(n_899), .Y(n_898) );
INVx2_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
NOR2x1p5_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
OAI21x1_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_900), .B(n_909), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g908 ( .A(n_901), .Y(n_908) );
NOR2xp33_ASAP7_75t_R g911 ( .A(n_912), .B(n_913), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_914), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_915), .Y(n_914) );
endmodule