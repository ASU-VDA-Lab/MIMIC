module fake_netlist_5_2092_n_1710 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1710);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1710;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_76),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_64),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_81),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_127),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_35),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_83),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_43),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_97),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_71),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_34),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_24),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_4),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_73),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_31),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_67),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_114),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_22),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_22),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_82),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_38),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_20),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_161),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_142),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_78),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_140),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_79),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_88),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_16),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_139),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_92),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_80),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_24),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_102),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_32),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_126),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_119),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_56),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_31),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_135),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_62),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_144),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_84),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_8),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_105),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_49),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_0),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_63),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_104),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_48),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_150),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_39),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_163),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_116),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_13),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_47),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_28),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_85),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_66),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_33),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_19),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_40),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_123),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_20),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_143),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_23),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_30),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_29),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_52),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_162),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_61),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_93),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_125),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_52),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_17),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_56),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_106),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_34),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_44),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_122),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_164),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_155),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_30),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_86),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_50),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_49),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_74),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_44),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_130),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_151),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_89),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_146),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_43),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_45),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_111),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_41),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_19),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_37),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_69),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_153),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_55),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_54),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_60),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_179),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_202),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_180),
.B(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_196),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_181),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_203),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_204),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_207),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_211),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_1),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_183),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_225),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_216),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_218),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_323),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_213),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_219),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_2),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_220),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_231),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_196),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_323),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_251),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_251),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_221),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_222),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_179),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_226),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_228),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_237),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_229),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_230),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_251),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_331),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_251),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_251),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_258),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_286),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_258),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_233),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_3),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_6),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_242),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_R g381 ( 
.A(n_243),
.B(n_98),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_258),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_244),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_247),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_250),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_200),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_168),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_168),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_253),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_269),
.B(n_6),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_258),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_260),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_267),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_270),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_272),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_174),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_291),
.B(n_8),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_258),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_290),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_297),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_297),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_297),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_299),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_297),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_297),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_254),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_274),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_291),
.B(n_9),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_205),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_169),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_274),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_254),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_R g415 ( 
.A(n_410),
.B(n_169),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_283),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_170),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_333),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_336),
.Y(n_430)
);

CKINVDCx8_ASAP7_75t_R g431 ( 
.A(n_375),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_340),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_359),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_341),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_359),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_342),
.B(n_317),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_343),
.B(n_317),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_347),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_369),
.B(n_167),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_348),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_350),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_358),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_353),
.B(n_210),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_339),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_334),
.B(n_186),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_355),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_361),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_399),
.B(n_193),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_362),
.B(n_174),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_398),
.A2(n_201),
.B(n_198),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_364),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_365),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_367),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_413),
.B(n_283),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_375),
.B(n_329),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_405),
.B(n_170),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_368),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_405),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_383),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_385),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_386),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_428),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_444),
.B(n_354),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_465),
.B(n_413),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_414),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_418),
.B1(n_419),
.B2(n_466),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_206),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_468),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_179),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_452),
.B(n_394),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_446),
.A2(n_419),
.B1(n_466),
.B2(n_417),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_438),
.A2(n_335),
.B1(n_354),
.B2(n_398),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_439),
.B(n_395),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_451),
.B(n_396),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_337),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_455),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_446),
.B(n_352),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_420),
.B(n_446),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_424),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_461),
.Y(n_521)
);

BUFx4f_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_461),
.B(n_412),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_424),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_461),
.B(n_215),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_377),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_461),
.B(n_352),
.Y(n_530)
);

AND3x2_ASAP7_75t_L g531 ( 
.A(n_474),
.B(n_391),
.C(n_256),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_473),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_421),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_380),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_473),
.B(n_388),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_476),
.B(n_241),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_474),
.B(n_409),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_427),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_476),
.B(n_252),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_466),
.B(n_389),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_429),
.B(n_311),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_415),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_432),
.B(n_390),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_434),
.B(n_409),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_425),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_453),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_441),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_456),
.A2(n_344),
.B1(n_378),
.B2(n_379),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_421),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_393),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_429),
.B(n_227),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_423),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_485),
.B(n_397),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_436),
.B(n_234),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_456),
.A2(n_344),
.B1(n_378),
.B2(n_379),
.Y(n_558)
);

INVx4_ASAP7_75t_SL g559 ( 
.A(n_456),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_436),
.B(n_236),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_437),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_485),
.B(n_246),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_437),
.B(n_442),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_486),
.B(n_487),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_448),
.B(n_279),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_457),
.B(n_188),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_440),
.Y(n_573)
);

OR2x2_ASAP7_75t_SL g574 ( 
.A(n_440),
.B(n_199),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_458),
.B(n_400),
.Y(n_575)
);

INVx4_ASAP7_75t_SL g576 ( 
.A(n_456),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_455),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_469),
.B(n_281),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_449),
.B(n_287),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_423),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_470),
.A2(n_235),
.B1(n_209),
.B2(n_223),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_463),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_472),
.B(n_404),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_477),
.A2(n_345),
.B1(n_370),
.B2(n_366),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_486),
.B(n_289),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_431),
.B(n_346),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_459),
.B(n_296),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_479),
.A2(n_356),
.B1(n_195),
.B2(n_192),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_482),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_463),
.B(n_314),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_316),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_423),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_440),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_471),
.B(n_327),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_423),
.Y(n_599)
);

BUFx8_ASAP7_75t_SL g600 ( 
.A(n_484),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_431),
.Y(n_601)
);

BUFx4f_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_440),
.B(n_248),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_384),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_423),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_481),
.B(n_328),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_433),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_456),
.A2(n_298),
.B1(n_214),
.B2(n_224),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_450),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_480),
.B(n_179),
.Y(n_612)
);

OAI21xp33_ASAP7_75t_SL g613 ( 
.A1(n_443),
.A2(n_310),
.B(n_285),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_450),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_450),
.B(n_384),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_443),
.B(n_334),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_450),
.B(n_171),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_450),
.B(n_171),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_450),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_443),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_454),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_454),
.B(n_334),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_454),
.B(n_172),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_460),
.B(n_172),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_483),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_460),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_460),
.B(n_239),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_467),
.A2(n_313),
.B1(n_276),
.B2(n_264),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_467),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_480),
.B(n_179),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_478),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_518),
.B(n_480),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_512),
.B(n_173),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_494),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_511),
.B(n_478),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_529),
.A2(n_190),
.B1(n_184),
.B2(n_176),
.Y(n_639)
);

AND2x6_ASAP7_75t_SL g640 ( 
.A(n_536),
.B(n_278),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_544),
.B(n_173),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_506),
.B(n_483),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_497),
.B(n_303),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_626),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_510),
.A2(n_190),
.B1(n_184),
.B2(n_176),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_626),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_537),
.B(n_178),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_544),
.B(n_175),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_514),
.B(n_175),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_509),
.B(n_179),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_631),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_600),
.B(n_208),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_538),
.B(n_483),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_510),
.A2(n_191),
.B1(n_195),
.B2(n_192),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_541),
.B(n_182),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_499),
.B(n_182),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_542),
.A2(n_300),
.B1(n_217),
.B2(n_282),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_498),
.B(n_185),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_615),
.B(n_189),
.Y(n_659)
);

OR2x2_ASAP7_75t_SL g660 ( 
.A(n_548),
.B(n_532),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_488),
.B(n_189),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_522),
.B(n_179),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_600),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_631),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_500),
.B(n_179),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_489),
.B(n_491),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_492),
.B(n_191),
.Y(n_667)
);

AOI221xp5_ASAP7_75t_L g668 ( 
.A1(n_490),
.A2(n_582),
.B1(n_539),
.B2(n_510),
.C(n_315),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_522),
.B(n_249),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_537),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_249),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_566),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_495),
.B(n_259),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_521),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_604),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_259),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_539),
.B(n_306),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_546),
.B(n_549),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_566),
.B(n_306),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_522),
.A2(n_312),
.B1(n_268),
.B2(n_257),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_521),
.B(n_602),
.Y(n_681)
);

AND2x6_ASAP7_75t_SL g682 ( 
.A(n_545),
.B(n_232),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_556),
.B(n_325),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_293),
.C(n_240),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_632),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_490),
.A2(n_546),
.B1(n_500),
.B2(n_516),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_566),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_552),
.A2(n_363),
.B(n_307),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_602),
.B(n_307),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_602),
.B(n_309),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_520),
.B(n_526),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_516),
.B(n_318),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_556),
.B(n_318),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_527),
.B(n_319),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_540),
.B(n_381),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_523),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_562),
.B(n_363),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_523),
.B(n_528),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_363),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_632),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_500),
.A2(n_530),
.B1(n_633),
.B2(n_612),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_523),
.B(n_255),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_568),
.B(n_245),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_569),
.B(n_261),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_612),
.A2(n_320),
.B1(n_326),
.B2(n_187),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_570),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_569),
.B(n_262),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_578),
.B(n_263),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_528),
.A2(n_288),
.B(n_265),
.C(n_266),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_528),
.B(n_551),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_496),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_571),
.B(n_593),
.Y(n_712)
);

AND2x4_ASAP7_75t_SL g713 ( 
.A(n_620),
.B(n_255),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_596),
.B(n_271),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_273),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_558),
.B(n_255),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_603),
.B(n_275),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_628),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_633),
.B(n_277),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_616),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_599),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_531),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_617),
.B(n_301),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_616),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_587),
.A2(n_604),
.B1(n_573),
.B2(n_595),
.Y(n_726)
);

INVx8_ASAP7_75t_L g727 ( 
.A(n_604),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_500),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_500),
.B(n_302),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_502),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_501),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_500),
.A2(n_178),
.B1(n_187),
.B2(n_324),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_620),
.Y(n_733)
);

INVx6_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_618),
.B(n_304),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_607),
.B(n_305),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_599),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_554),
.A2(n_197),
.B1(n_308),
.B2(n_324),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_605),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_590),
.B(n_329),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_577),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_578),
.B(n_295),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_563),
.A2(n_294),
.B(n_280),
.C(n_284),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_564),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_583),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_624),
.B(n_292),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_623),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_563),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_625),
.B(n_197),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_543),
.B(n_308),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_563),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_504),
.B(n_321),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_592),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_553),
.B(n_329),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_530),
.A2(n_589),
.B1(n_586),
.B2(n_610),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_592),
.B(n_321),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_515),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_572),
.Y(n_758)
);

INVxp67_ASAP7_75t_SL g759 ( 
.A(n_599),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_581),
.B(n_315),
.Y(n_760)
);

AND2x6_ASAP7_75t_L g761 ( 
.A(n_623),
.B(n_325),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_557),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_504),
.B(n_157),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_502),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_586),
.B(n_10),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_517),
.B(n_154),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_554),
.A2(n_152),
.B1(n_148),
.B2(n_147),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_611),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_561),
.B(n_11),
.Y(n_769)
);

AND2x6_ASAP7_75t_SL g770 ( 
.A(n_575),
.B(n_13),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_614),
.A2(n_121),
.B(n_117),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_517),
.B(n_108),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_554),
.A2(n_101),
.B1(n_96),
.B2(n_95),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_580),
.B(n_14),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_505),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_SL g776 ( 
.A(n_504),
.B(n_14),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_504),
.B(n_94),
.Y(n_777)
);

O2A1O1Ixp5_ASAP7_75t_L g778 ( 
.A1(n_588),
.A2(n_91),
.B(n_90),
.C(n_77),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_507),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_517),
.B(n_75),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_601),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_519),
.B(n_68),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_519),
.B(n_65),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_584),
.B(n_15),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_591),
.B(n_15),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_601),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_519),
.B(n_58),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_507),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_508),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_554),
.A2(n_503),
.B1(n_634),
.B2(n_560),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_611),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_585),
.B(n_17),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_18),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_534),
.B(n_21),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_608),
.A2(n_26),
.B(n_27),
.C(n_29),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_629),
.B(n_32),
.C(n_33),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_534),
.B(n_37),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_534),
.B(n_57),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_508),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_721),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_L g801 ( 
.A1(n_704),
.A2(n_595),
.B(n_573),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_710),
.A2(n_513),
.B(n_535),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_649),
.A2(n_613),
.B(n_503),
.C(n_550),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_594),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_663),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_710),
.A2(n_513),
.B(n_535),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_650),
.A2(n_622),
.B(n_630),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_744),
.B(n_634),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_698),
.A2(n_579),
.B(n_555),
.Y(n_809)
);

BUFx12f_ASAP7_75t_L g810 ( 
.A(n_757),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_680),
.A2(n_574),
.B1(n_550),
.B2(n_604),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_739),
.B(n_577),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_745),
.B(n_594),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_642),
.B(n_594),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_698),
.A2(n_579),
.B(n_513),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_674),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_731),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_681),
.A2(n_535),
.B(n_579),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_650),
.A2(n_627),
.B(n_533),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_681),
.A2(n_555),
.B(n_504),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_704),
.A2(n_708),
.B(n_707),
.Y(n_821)
);

OA22x2_ASAP7_75t_L g822 ( 
.A1(n_645),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_725),
.Y(n_823)
);

OR2x2_ASAP7_75t_SL g824 ( 
.A(n_792),
.B(n_42),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_686),
.B(n_619),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_674),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_674),
.Y(n_827)
);

BUFx12f_ASAP7_75t_L g828 ( 
.A(n_660),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_747),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_676),
.A2(n_621),
.B(n_609),
.C(n_565),
.Y(n_830)
);

OAI22x1_ASAP7_75t_L g831 ( 
.A1(n_654),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_638),
.A2(n_555),
.B(n_619),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_636),
.B(n_554),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_683),
.B(n_621),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_768),
.A2(n_619),
.B(n_599),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_636),
.A2(n_554),
.B1(n_606),
.B2(n_547),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_674),
.B(n_606),
.Y(n_837)
);

AO21x1_ASAP7_75t_L g838 ( 
.A1(n_662),
.A2(n_525),
.B(n_565),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_747),
.B(n_524),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_791),
.A2(n_524),
.B(n_560),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_672),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_680),
.A2(n_547),
.B1(n_525),
.B2(n_53),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_722),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_677),
.A2(n_559),
.B(n_576),
.C(n_53),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_740),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_L g846 ( 
.A1(n_707),
.A2(n_46),
.B(n_50),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_653),
.A2(n_559),
.B(n_576),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_701),
.A2(n_54),
.B1(n_57),
.B2(n_559),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_790),
.A2(n_759),
.B(n_662),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_790),
.A2(n_559),
.B(n_576),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_666),
.A2(n_576),
.B(n_691),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_687),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_755),
.A2(n_678),
.B1(n_708),
.B2(n_742),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_670),
.B(n_647),
.Y(n_854)
);

AOI21x1_ASAP7_75t_L g855 ( 
.A1(n_697),
.A2(n_699),
.B(n_669),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_696),
.B(n_753),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_669),
.A2(n_799),
.B(n_775),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_786),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_656),
.A2(n_778),
.B(n_668),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_655),
.B(n_677),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_705),
.A2(n_732),
.B1(n_738),
.B2(n_742),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_706),
.B(n_712),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_711),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_644),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_722),
.A2(n_737),
.B(n_665),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_646),
.Y(n_866)
);

INVx11_ASAP7_75t_L g867 ( 
.A(n_761),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_722),
.A2(n_737),
.B(n_651),
.Y(n_868)
);

O2A1O1Ixp5_ASAP7_75t_L g869 ( 
.A1(n_720),
.A2(n_735),
.B(n_724),
.C(n_690),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_722),
.A2(n_737),
.B(n_664),
.Y(n_870)
);

AOI21x1_ASAP7_75t_L g871 ( 
.A1(n_764),
.A2(n_689),
.B(n_690),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_748),
.B(n_751),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_659),
.B(n_746),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_719),
.B(n_769),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_760),
.A2(n_714),
.B(n_685),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_724),
.A2(n_735),
.B(n_772),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_700),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_705),
.B(n_648),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_723),
.A2(n_758),
.B1(n_720),
.B2(n_692),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_692),
.A2(n_635),
.B1(n_702),
.B2(n_761),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_695),
.A2(n_729),
.B(n_679),
.Y(n_881)
);

O2A1O1Ixp5_ASAP7_75t_L g882 ( 
.A1(n_702),
.A2(n_798),
.B(n_797),
.C(n_794),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_781),
.B(n_754),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_766),
.A2(n_783),
.B(n_782),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_750),
.B(n_749),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_762),
.A2(n_795),
.B(n_769),
.C(n_793),
.Y(n_886)
);

OAI321xp33_ASAP7_75t_L g887 ( 
.A1(n_732),
.A2(n_738),
.A3(n_657),
.B1(n_784),
.B2(n_765),
.C(n_796),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_780),
.A2(n_671),
.B(n_667),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_643),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_774),
.A2(n_785),
.B(n_793),
.C(n_756),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_657),
.A2(n_717),
.B1(n_639),
.B2(n_765),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_661),
.A2(n_673),
.B(n_789),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_728),
.B(n_767),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_774),
.A2(n_785),
.B(n_756),
.C(n_717),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_730),
.A2(n_788),
.B(n_779),
.Y(n_895)
);

INVx11_ASAP7_75t_L g896 ( 
.A(n_761),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_743),
.A2(n_709),
.B(n_688),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_658),
.A2(n_777),
.B(n_763),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_763),
.A2(n_777),
.B(n_728),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_703),
.A2(n_718),
.B(n_736),
.Y(n_901)
);

CKINVDCx10_ASAP7_75t_R g902 ( 
.A(n_733),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_643),
.A2(n_716),
.B(n_715),
.C(n_693),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_761),
.A2(n_684),
.B1(n_752),
.B2(n_787),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_641),
.B(n_786),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_694),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_726),
.B(n_675),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_734),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_635),
.B(n_726),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_752),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_771),
.A2(n_773),
.B(n_675),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_761),
.A2(n_776),
.B(n_741),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_652),
.A2(n_640),
.B(n_682),
.C(n_675),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_713),
.B(n_727),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_727),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_733),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_SL g917 ( 
.A(n_734),
.B(n_727),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_713),
.B(n_680),
.C(n_649),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_770),
.A2(n_522),
.B(n_650),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_649),
.B(n_744),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_686),
.A2(n_636),
.B1(n_745),
.B2(n_744),
.Y(n_922)
);

CKINVDCx8_ASAP7_75t_R g923 ( 
.A(n_682),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_704),
.A2(n_708),
.B(n_707),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_757),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_650),
.A2(n_522),
.B(n_662),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_733),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_757),
.B(n_465),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_676),
.A2(n_542),
.B(n_656),
.C(n_678),
.Y(n_930)
);

OAI321xp33_ASAP7_75t_L g931 ( 
.A1(n_705),
.A2(n_680),
.A3(n_668),
.B1(n_649),
.B2(n_645),
.C(n_654),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_680),
.B(n_649),
.C(n_704),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_676),
.A2(n_542),
.B(n_656),
.C(n_678),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_757),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_739),
.B(n_544),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_649),
.B(n_744),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_649),
.B(n_744),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_662),
.A2(n_650),
.B(n_518),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_637),
.B(n_444),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_649),
.B(n_744),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_649),
.A2(n_677),
.B(n_707),
.C(n_704),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_672),
.B(n_687),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_739),
.B(n_544),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_670),
.B(n_465),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_637),
.B(n_444),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_739),
.B(n_544),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_674),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_674),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_649),
.B(n_744),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_649),
.B(n_744),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_649),
.B(n_744),
.Y(n_956)
);

BUFx4f_ASAP7_75t_L g957 ( 
.A(n_734),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_757),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_649),
.B(n_744),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_757),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_649),
.B(n_744),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_662),
.A2(n_650),
.B(n_518),
.Y(n_963)
);

BUFx12f_ASAP7_75t_L g964 ( 
.A(n_757),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_680),
.A2(n_509),
.B1(n_499),
.B2(n_686),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_649),
.B(n_744),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_649),
.B(n_744),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_649),
.B(n_744),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_705),
.B(n_544),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_662),
.A2(n_650),
.B(n_518),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_674),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_649),
.A2(n_677),
.B(n_707),
.C(n_704),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_744),
.B(n_745),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_710),
.A2(n_698),
.B(n_509),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_674),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_821),
.A2(n_924),
.B1(n_932),
.B2(n_942),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_958),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_972),
.A2(n_929),
.B(n_920),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_SL g980 ( 
.A1(n_890),
.A2(n_894),
.B(n_861),
.C(n_803),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_938),
.A2(n_947),
.B(n_945),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_805),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_940),
.B(n_948),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_965),
.A2(n_861),
.B1(n_853),
.B2(n_974),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_872),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_SL g986 ( 
.A1(n_974),
.A2(n_922),
.B(n_965),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_950),
.A2(n_959),
.B(n_954),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_973),
.A2(n_975),
.B(n_849),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_856),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_L g991 ( 
.A1(n_891),
.A2(n_931),
.B(n_887),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_908),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_859),
.A2(n_926),
.B(n_930),
.Y(n_993)
);

AO21x2_ASAP7_75t_L g994 ( 
.A1(n_859),
.A2(n_825),
.B(n_880),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_819),
.A2(n_875),
.B(n_865),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_935),
.B(n_944),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_900),
.A2(n_850),
.B(n_898),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_921),
.A2(n_962),
.B1(n_956),
.B2(n_960),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_SL g999 ( 
.A1(n_926),
.A2(n_833),
.B(n_933),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_816),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_881),
.A2(n_884),
.B(n_888),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_856),
.B(n_915),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_936),
.B(n_937),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_908),
.Y(n_1004)
);

O2A1O1Ixp5_ASAP7_75t_L g1005 ( 
.A1(n_882),
.A2(n_860),
.B(n_953),
.C(n_967),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_941),
.B(n_955),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_819),
.A2(n_807),
.B(n_855),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_939),
.A2(n_963),
.B(n_970),
.Y(n_1008)
);

OA21x2_ASAP7_75t_L g1009 ( 
.A1(n_869),
.A2(n_807),
.B(n_804),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_908),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_886),
.A2(n_848),
.B(n_842),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_927),
.Y(n_1012)
);

INVxp33_ASAP7_75t_SL g1013 ( 
.A(n_812),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_857),
.A2(n_871),
.B(n_876),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_832),
.A2(n_901),
.B(n_814),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_966),
.B(n_968),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_830),
.A2(n_840),
.B(n_815),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_949),
.B(n_885),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_892),
.A2(n_809),
.B(n_873),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_931),
.A2(n_887),
.B(n_897),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_851),
.A2(n_838),
.B(n_870),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_862),
.A2(n_808),
.B(n_911),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_835),
.A2(n_868),
.B(n_820),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_848),
.A2(n_842),
.A3(n_844),
.B(n_903),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_946),
.B(n_845),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_879),
.A2(n_878),
.B(n_909),
.C(n_906),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_895),
.A2(n_839),
.B(n_837),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_808),
.B(n_834),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_813),
.A2(n_847),
.B(n_877),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_897),
.A2(n_919),
.B(n_910),
.Y(n_1030)
);

AO21x1_ASAP7_75t_L g1031 ( 
.A1(n_969),
.A2(n_874),
.B(n_907),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_836),
.A2(n_904),
.B(n_826),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_810),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_961),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_SL g1035 ( 
.A1(n_951),
.A2(n_827),
.B(n_816),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_845),
.B(n_854),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_952),
.A2(n_976),
.B(n_971),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_943),
.B(n_858),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_907),
.A2(n_883),
.B1(n_905),
.B2(n_811),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_843),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_919),
.A2(n_846),
.B(n_801),
.C(n_852),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_843),
.A2(n_829),
.B(n_823),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_961),
.Y(n_1043)
);

OAI22x1_ASAP7_75t_L g1044 ( 
.A1(n_914),
.A2(n_925),
.B1(n_824),
.B2(n_863),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_841),
.B(n_943),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_831),
.A2(n_811),
.A3(n_866),
.B(n_864),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_951),
.A2(n_827),
.B(n_957),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_917),
.B(n_899),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_912),
.A2(n_822),
.B(n_893),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_817),
.B(n_934),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_928),
.B(n_964),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_912),
.A2(n_822),
.B(n_867),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_893),
.B(n_899),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_913),
.A2(n_957),
.B(n_916),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_L g1055 ( 
.A(n_893),
.B(n_896),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_893),
.A2(n_828),
.B(n_927),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_923),
.B(n_902),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_940),
.B(n_465),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_821),
.A2(n_924),
.B(n_972),
.C(n_942),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_SL g1062 ( 
.A1(n_919),
.A2(n_938),
.B(n_920),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_974),
.B(n_921),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_965),
.A2(n_942),
.B1(n_972),
.B2(n_932),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1066)
);

AOI211x1_ASAP7_75t_L g1067 ( 
.A1(n_861),
.A2(n_924),
.B(n_821),
.C(n_932),
.Y(n_1067)
);

XOR2xp5_ASAP7_75t_L g1068 ( 
.A(n_805),
.B(n_453),
.Y(n_1068)
);

AOI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_932),
.A2(n_861),
.B(n_821),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_974),
.B(n_921),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_SL g1072 ( 
.A1(n_965),
.A2(n_972),
.B(n_942),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_974),
.B(n_921),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_908),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_821),
.A2(n_924),
.B(n_972),
.C(n_942),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_821),
.A2(n_924),
.B1(n_932),
.B2(n_942),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_942),
.A2(n_972),
.A3(n_838),
.B(n_890),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_965),
.A2(n_942),
.B1(n_972),
.B2(n_932),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_974),
.B(n_921),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_805),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_919),
.A2(n_938),
.B(n_920),
.Y(n_1082)
);

AO21x2_ASAP7_75t_L g1083 ( 
.A1(n_859),
.A2(n_972),
.B(n_942),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_810),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_942),
.A2(n_972),
.A3(n_838),
.B(n_890),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_889),
.B(n_856),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_816),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_800),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_974),
.B(n_921),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_974),
.B(n_921),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_974),
.B(n_921),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_872),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_940),
.B(n_465),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_974),
.B(n_921),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_942),
.A2(n_972),
.B(n_890),
.C(n_894),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_932),
.A2(n_861),
.B(n_821),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_872),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_940),
.B(n_465),
.Y(n_1103)
);

AOI221x1_ASAP7_75t_L g1104 ( 
.A1(n_942),
.A2(n_972),
.B1(n_924),
.B2(n_821),
.C(n_932),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_821),
.A2(n_924),
.B(n_972),
.C(n_942),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_872),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_800),
.Y(n_1107)
);

AOI21xp33_ASAP7_75t_L g1108 ( 
.A1(n_932),
.A2(n_861),
.B(n_821),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_974),
.B(n_921),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_917),
.B(n_951),
.Y(n_1111)
);

OAI22x1_ASAP7_75t_L g1112 ( 
.A1(n_932),
.A2(n_853),
.B1(n_918),
.B2(n_879),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_816),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_920),
.A2(n_938),
.B(n_929),
.Y(n_1114)
);

AOI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_932),
.A2(n_861),
.B(n_821),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_802),
.A2(n_806),
.B(n_818),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_942),
.A2(n_972),
.B(n_932),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1038),
.B(n_1002),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1060),
.B(n_1097),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_991),
.A2(n_1061),
.B(n_1076),
.C(n_1105),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1043),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1001),
.A2(n_1019),
.B(n_1072),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_982),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1034),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_L g1128 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_978),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1103),
.B(n_983),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1015),
.A2(n_1022),
.B(n_999),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1073),
.B(n_1080),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1073),
.B(n_1080),
.Y(n_1133)
);

CKINVDCx11_ASAP7_75t_R g1134 ( 
.A(n_1012),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_1040),
.B(n_992),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1090),
.B(n_1093),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1090),
.A2(n_1095),
.B1(n_1109),
.B2(n_1093),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1095),
.B(n_1099),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1089),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1020),
.A2(n_1100),
.B(n_1064),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_SL g1141 ( 
.A(n_1053),
.B(n_985),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1107),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1081),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1069),
.A2(n_1115),
.B(n_1108),
.C(n_1101),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1038),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1018),
.B(n_996),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_987),
.A2(n_1058),
.B(n_1091),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_998),
.A2(n_1115),
.B(n_1108),
.C(n_1101),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_1039),
.B(n_1055),
.Y(n_1149)
);

BUFx8_ASAP7_75t_SL g1150 ( 
.A(n_1033),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1003),
.B(n_1006),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1064),
.A2(n_1079),
.B1(n_984),
.B2(n_1013),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1004),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1099),
.B(n_1109),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_1025),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1003),
.B(n_1006),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1036),
.B(n_1016),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1119),
.A2(n_986),
.B(n_984),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1096),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1059),
.A2(n_1075),
.B(n_1065),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_1004),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1002),
.B(n_990),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_990),
.B(n_1087),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1016),
.B(n_998),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1011),
.A2(n_1112),
.B1(n_1031),
.B2(n_1083),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1102),
.B(n_1106),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1070),
.A2(n_1110),
.B(n_1114),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_1010),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1035),
.B(n_1053),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_989),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1028),
.B(n_1026),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_1010),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_977),
.A2(n_1077),
.B1(n_1067),
.B2(n_1028),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1087),
.B(n_1050),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1049),
.A2(n_1041),
.B1(n_993),
.B2(n_979),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1068),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1051),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1088),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1104),
.A2(n_997),
.A3(n_1032),
.B(n_1029),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1046),
.B(n_1083),
.Y(n_1181)
);

CKINVDCx11_ASAP7_75t_R g1182 ( 
.A(n_1084),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_1046),
.B(n_1044),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1010),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1074),
.B(n_1056),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1074),
.B(n_1113),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1030),
.B(n_1054),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_979),
.A2(n_994),
.B1(n_1030),
.B2(n_1082),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1088),
.B(n_1113),
.Y(n_1189)
);

BUFx4_ASAP7_75t_SL g1190 ( 
.A(n_1054),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_981),
.A2(n_980),
.B(n_994),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1047),
.B(n_1052),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1000),
.B(n_1085),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1048),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_981),
.B(n_1085),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_SL g1196 ( 
.A(n_1057),
.B(n_1042),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1007),
.A2(n_995),
.B(n_1005),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1062),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1021),
.A2(n_1014),
.B(n_1008),
.C(n_1037),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1057),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_988),
.A2(n_1118),
.B(n_1117),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1009),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1024),
.B(n_1078),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1024),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1027),
.B(n_1017),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1066),
.A2(n_1086),
.B(n_1092),
.C(n_1094),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1116),
.A2(n_1098),
.B(n_1023),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1018),
.B(n_821),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1001),
.A2(n_1019),
.B(n_1072),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1001),
.A2(n_1019),
.B(n_1072),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1034),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1018),
.B(n_996),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_982),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1043),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1060),
.B(n_1097),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_991),
.A2(n_932),
.B1(n_924),
.B2(n_821),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1111),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1060),
.B(n_1097),
.Y(n_1219)
);

OAI221xp5_ASAP7_75t_L g1220 ( 
.A1(n_991),
.A2(n_924),
.B1(n_821),
.B2(n_932),
.C(n_861),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1001),
.A2(n_1019),
.B(n_1072),
.Y(n_1221)
);

BUFx4_ASAP7_75t_SL g1222 ( 
.A(n_1084),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_993),
.A2(n_1007),
.B(n_979),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1034),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1063),
.A2(n_965),
.B1(n_1073),
.B2(n_1071),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1001),
.A2(n_1019),
.B(n_1072),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1018),
.B(n_972),
.C(n_942),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_SL g1228 ( 
.A1(n_996),
.A2(n_824),
.B1(n_861),
.B2(n_680),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1060),
.B(n_1097),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_982),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1039),
.A2(n_969),
.B1(n_932),
.B2(n_474),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1018),
.B(n_996),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1111),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1038),
.B(n_1002),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_982),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1038),
.B(n_1002),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1018),
.B(n_972),
.C(n_942),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1063),
.A2(n_965),
.B1(n_1073),
.B2(n_1071),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1242)
);

BUFx8_ASAP7_75t_L g1243 ( 
.A(n_1033),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1045),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1034),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1043),
.Y(n_1246)
);

AO21x1_ASAP7_75t_L g1247 ( 
.A1(n_991),
.A2(n_1079),
.B(n_1064),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1204),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1193),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1143),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1154),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1228),
.A2(n_1213),
.B1(n_1146),
.B2(n_1235),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1246),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_1126),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1160),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1123),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1234),
.A2(n_1153),
.B1(n_1240),
.B2(n_1227),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1162),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1144),
.A2(n_1148),
.B(n_1220),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_1134),
.Y(n_1260)
);

AO21x1_ASAP7_75t_L g1261 ( 
.A1(n_1176),
.A2(n_1122),
.B(n_1140),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1215),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1157),
.B(n_1187),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1152),
.B(n_1167),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1141),
.A2(n_1172),
.B(n_1247),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1220),
.A2(n_1149),
.B1(n_1208),
.B2(n_1159),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1169),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1159),
.A2(n_1217),
.B1(n_1140),
.B2(n_1128),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1124),
.B(n_1132),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1151),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_R g1271 ( 
.A(n_1214),
.B(n_1238),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1127),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1174),
.A2(n_1194),
.B1(n_1183),
.B2(n_1203),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1230),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1216),
.B(n_1219),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1130),
.B(n_1124),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1174),
.A2(n_1203),
.B1(n_1165),
.B2(n_1137),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1137),
.A2(n_1225),
.B1(n_1241),
.B2(n_1242),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1132),
.A2(n_1155),
.B1(n_1231),
.B2(n_1232),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1176),
.A2(n_1190),
.B1(n_1232),
.B2(n_1231),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1156),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1192),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1181),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1201),
.A2(n_1207),
.B(n_1131),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1133),
.B(n_1136),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1171),
.A2(n_1168),
.B(n_1147),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1201),
.A2(n_1207),
.B(n_1131),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1192),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1225),
.A2(n_1241),
.B1(n_1198),
.B2(n_1175),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1172),
.A2(n_1196),
.B1(n_1166),
.B2(n_1164),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1192),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1195),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1173),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1170),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1121),
.A2(n_1229),
.B1(n_1136),
.B2(n_1138),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1170),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1182),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1170),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1195),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1129),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1211),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1133),
.A2(n_1212),
.B1(n_1155),
.B2(n_1242),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1224),
.Y(n_1303)
);

INVx4_ASAP7_75t_SL g1304 ( 
.A(n_1185),
.Y(n_1304)
);

OR2x6_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_1209),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1120),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_L g1307 ( 
.A(n_1163),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1245),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1138),
.A2(n_1233),
.B1(n_1212),
.B2(n_1158),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1180),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1233),
.A2(n_1125),
.B(n_1226),
.Y(n_1311)
);

AOI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1205),
.A2(n_1209),
.B(n_1210),
.Y(n_1312)
);

BUFx8_ASAP7_75t_L g1313 ( 
.A(n_1145),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1180),
.Y(n_1314)
);

CKINVDCx16_ASAP7_75t_R g1315 ( 
.A(n_1120),
.Y(n_1315)
);

BUFx2_ASAP7_75t_SL g1316 ( 
.A(n_1185),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1200),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1244),
.B(n_1223),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1150),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1191),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1191),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1178),
.B(n_1164),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1188),
.B(n_1142),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1199),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1177),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1210),
.A2(n_1221),
.B(n_1226),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1237),
.B(n_1239),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1202),
.B(n_1236),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1237),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1221),
.A2(n_1147),
.B(n_1161),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1139),
.B(n_1218),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1197),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1197),
.B(n_1161),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1222),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1243),
.A2(n_1186),
.B1(n_1189),
.B2(n_1179),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1206),
.B(n_1135),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1189),
.Y(n_1337)
);

AO21x1_ASAP7_75t_L g1338 ( 
.A1(n_1184),
.A2(n_991),
.B(n_1064),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1243),
.Y(n_1339)
);

AOI222xp33_ASAP7_75t_L g1340 ( 
.A1(n_1228),
.A2(n_861),
.B1(n_1146),
.B2(n_1235),
.C1(n_1213),
.C2(n_932),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1228),
.A2(n_932),
.B1(n_924),
.B2(n_821),
.Y(n_1341)
);

NAND2x1_ASAP7_75t_L g1342 ( 
.A(n_1192),
.B(n_1170),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1192),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1134),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1228),
.A2(n_932),
.B1(n_924),
.B2(n_821),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1201),
.A2(n_997),
.B(n_1207),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1248),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1269),
.B(n_1285),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1318),
.B(n_1292),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1262),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1330),
.A2(n_1311),
.B(n_1259),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1318),
.B(n_1292),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1312),
.A2(n_1326),
.B(n_1347),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1282),
.B(n_1288),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1299),
.B(n_1283),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1332),
.Y(n_1357)
);

BUFx2_ASAP7_75t_SL g1358 ( 
.A(n_1258),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1299),
.B(n_1249),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1269),
.B(n_1285),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1321),
.A2(n_1287),
.B(n_1284),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1296),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1309),
.B(n_1279),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1333),
.A2(n_1342),
.B(n_1324),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1310),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1284),
.A2(n_1287),
.B(n_1324),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1314),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1282),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1288),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1288),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1257),
.A2(n_1340),
.B(n_1341),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1302),
.B(n_1343),
.Y(n_1372)
);

BUFx12f_ASAP7_75t_L g1373 ( 
.A(n_1260),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1291),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1291),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1344),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1263),
.B(n_1278),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1286),
.B(n_1278),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1344),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_1338),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1343),
.B(n_1264),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1250),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1274),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1261),
.B(n_1323),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1305),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1262),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1281),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1265),
.A2(n_1257),
.B(n_1323),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1294),
.B(n_1298),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1305),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1265),
.A2(n_1294),
.B(n_1298),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1305),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1298),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1355),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1355),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1371),
.B(n_1295),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1364),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1350),
.B(n_1277),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1350),
.B(n_1336),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1371),
.A2(n_1252),
.B1(n_1346),
.B2(n_1266),
.Y(n_1401)
);

OAI222xp33_ASAP7_75t_L g1402 ( 
.A1(n_1363),
.A2(n_1280),
.B1(n_1268),
.B2(n_1273),
.C1(n_1290),
.C2(n_1276),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1363),
.B(n_1270),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1372),
.B(n_1381),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1378),
.B(n_1352),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1356),
.B(n_1270),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1256),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1353),
.B(n_1384),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1384),
.B(n_1328),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1385),
.B(n_1304),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1348),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1380),
.A2(n_1335),
.B1(n_1275),
.B2(n_1315),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1352),
.B(n_1255),
.Y(n_1413)
);

INVx2_ASAP7_75t_R g1414 ( 
.A(n_1365),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1356),
.B(n_1377),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1380),
.A2(n_1271),
.B(n_1258),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1381),
.A2(n_1322),
.B1(n_1253),
.B2(n_1272),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1378),
.B(n_1316),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1357),
.B(n_1367),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1372),
.A2(n_1317),
.B1(n_1329),
.B2(n_1335),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1357),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1357),
.B(n_1331),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1377),
.B(n_1304),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1366),
.B(n_1361),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1397),
.B(n_1375),
.C(n_1369),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1397),
.A2(n_1387),
.B(n_1392),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1403),
.B(n_1360),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1401),
.B(n_1369),
.C(n_1368),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1360),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1412),
.B(n_1390),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_SL g1433 ( 
.A(n_1412),
.B(n_1382),
.C(n_1250),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1401),
.A2(n_1387),
.B(n_1392),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1411),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1420),
.B(n_1390),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1407),
.B(n_1389),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1420),
.B(n_1417),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1417),
.B(n_1390),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1402),
.A2(n_1388),
.B(n_1339),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1408),
.B(n_1359),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1416),
.A2(n_1388),
.B1(n_1315),
.B2(n_1307),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1405),
.B(n_1370),
.C(n_1368),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1405),
.B(n_1376),
.C(n_1370),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1410),
.A2(n_1383),
.B1(n_1319),
.B2(n_1339),
.Y(n_1445)
);

OAI221xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1405),
.A2(n_1388),
.B1(n_1300),
.B2(n_1362),
.C(n_1393),
.Y(n_1446)
);

OAI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1407),
.A2(n_1394),
.B(n_1386),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1415),
.B(n_1389),
.Y(n_1448)
);

NAND3xp33_ASAP7_75t_SL g1449 ( 
.A(n_1407),
.B(n_1301),
.C(n_1303),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1413),
.B(n_1379),
.C(n_1376),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1406),
.B(n_1389),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1406),
.B(n_1389),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1399),
.A2(n_1373),
.B1(n_1385),
.B2(n_1391),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1418),
.A2(n_1393),
.B1(n_1391),
.B2(n_1374),
.C(n_1301),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1421),
.A2(n_1354),
.B(n_1364),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1402),
.B(n_1374),
.Y(n_1456)
);

OA211x2_ASAP7_75t_L g1457 ( 
.A1(n_1424),
.A2(n_1358),
.B(n_1373),
.C(n_1327),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1399),
.A2(n_1334),
.B(n_1393),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1421),
.A2(n_1354),
.B(n_1364),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1424),
.A2(n_1307),
.B1(n_1306),
.B2(n_1308),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1413),
.B(n_1351),
.C(n_1386),
.D(n_1251),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1413),
.B(n_1390),
.Y(n_1462)
);

OAI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1418),
.A2(n_1391),
.B1(n_1306),
.B2(n_1307),
.C(n_1337),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1411),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1399),
.A2(n_1390),
.B(n_1373),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1435),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1464),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1441),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1448),
.B(n_1425),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1450),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1451),
.B(n_1425),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1443),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1445),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1432),
.B(n_1398),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1462),
.B(n_1414),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1455),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1444),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1462),
.B(n_1414),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1455),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1455),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1459),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1437),
.B(n_1419),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1427),
.B(n_1422),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1428),
.B(n_1410),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1429),
.B(n_1423),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1431),
.B(n_1423),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1426),
.B(n_1422),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1432),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1434),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1439),
.B(n_1419),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1400),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1436),
.B(n_1398),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1447),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1491),
.B(n_1395),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1467),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1493),
.B(n_1396),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1488),
.B(n_1423),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1488),
.B(n_1469),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1494),
.B(n_1456),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1476),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1466),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1491),
.B(n_1395),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1476),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1491),
.B(n_1395),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1466),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1469),
.B(n_1454),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1481),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1474),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1494),
.B(n_1456),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1297),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1495),
.B(n_1409),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1471),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1473),
.A2(n_1440),
.B1(n_1438),
.B2(n_1433),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1486),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1468),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1468),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1472),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1481),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1486),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1486),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1487),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1471),
.B(n_1418),
.Y(n_1530)
);

NAND2x1_ASAP7_75t_L g1531 ( 
.A(n_1493),
.B(n_1398),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1487),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1497),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1524),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1497),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1524),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1489),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

NOR2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1345),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1519),
.B(n_1477),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_1489),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1518),
.A2(n_1490),
.B1(n_1485),
.B2(n_1438),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1498),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1515),
.A2(n_1490),
.B1(n_1474),
.B2(n_1477),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1520),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1470),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1520),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1521),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1492),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1500),
.B(n_1471),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1526),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1527),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1527),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1502),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1528),
.B(n_1483),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1528),
.B(n_1483),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_1492),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1478),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1532),
.A2(n_1485),
.B1(n_1446),
.B2(n_1442),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1496),
.B(n_1493),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1496),
.B(n_1493),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1499),
.B(n_1492),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1505),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1502),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1505),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1543),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1517),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1563),
.Y(n_1578)
);

AO21x2_ASAP7_75t_L g1579 ( 
.A1(n_1554),
.A2(n_1504),
.B(n_1502),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1580)
);

OAI21xp33_ASAP7_75t_L g1581 ( 
.A1(n_1546),
.A2(n_1430),
.B(n_1436),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1536),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1569),
.A2(n_1457),
.B1(n_1460),
.B2(n_1458),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1563),
.Y(n_1586)
);

NAND2x1_ASAP7_75t_L g1587 ( 
.A(n_1547),
.B(n_1475),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1574),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1542),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1548),
.A2(n_1453),
.B1(n_1461),
.B2(n_1463),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1574),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1533),
.B(n_1499),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.B(n_1531),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1535),
.B(n_1507),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1537),
.B(n_1541),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1538),
.B(n_1465),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1551),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1535),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1535),
.B(n_1507),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1545),
.B(n_1531),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1534),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1534),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1560),
.B(n_1509),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1555),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1506),
.Y(n_1611)
);

XNOR2x1_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1589),
.Y(n_1612)
);

O2A1O1Ixp5_ASAP7_75t_L g1613 ( 
.A1(n_1587),
.A2(n_1539),
.B(n_1561),
.C(n_1550),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1582),
.B(n_1558),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1581),
.B(n_1557),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1581),
.A2(n_1562),
.B(n_1271),
.Y(n_1616)
);

CKINVDCx16_ASAP7_75t_R g1617 ( 
.A(n_1589),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1609),
.A2(n_1566),
.B(n_1557),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1584),
.A2(n_1609),
.B1(n_1598),
.B2(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1590),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1598),
.A2(n_1572),
.B1(n_1530),
.B2(n_1517),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1585),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1567),
.Y(n_1624)
);

OAI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1595),
.A2(n_1567),
.B(n_1545),
.C(n_1559),
.Y(n_1625)
);

OAI322xp33_ASAP7_75t_L g1626 ( 
.A1(n_1576),
.A2(n_1575),
.A3(n_1573),
.B1(n_1530),
.B2(n_1478),
.C1(n_1565),
.C2(n_1564),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1585),
.Y(n_1627)
);

OAI32xp33_ASAP7_75t_L g1628 ( 
.A1(n_1600),
.A2(n_1559),
.A3(n_1480),
.B1(n_1482),
.B2(n_1478),
.Y(n_1628)
);

INVxp67_ASAP7_75t_SL g1629 ( 
.A(n_1595),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1592),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1592),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1610),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1598),
.A2(n_1565),
.B1(n_1564),
.B2(n_1479),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1591),
.A2(n_1571),
.B1(n_1570),
.B2(n_1484),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1603),
.B(n_1506),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1617),
.B(n_1580),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1631),
.B(n_1580),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1629),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1612),
.B(n_1345),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1618),
.B(n_1583),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1621),
.B(n_1583),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1635),
.B(n_1598),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1614),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1614),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1620),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1594),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1615),
.A2(n_1616),
.B1(n_1636),
.B2(n_1625),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1619),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1613),
.B(n_1598),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1637),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1623),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1594),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1630),
.B(n_1577),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1637),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1632),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1650),
.A2(n_1622),
.B(n_1600),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1648),
.A2(n_1650),
.B1(n_1641),
.B2(n_1651),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1648),
.B(n_1633),
.C(n_1634),
.Y(n_1661)
);

AOI222xp33_ASAP7_75t_L g1662 ( 
.A1(n_1652),
.A2(n_1603),
.B1(n_1604),
.B2(n_1628),
.C1(n_1597),
.C2(n_1599),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_R g1663 ( 
.A(n_1652),
.B(n_1297),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1649),
.A2(n_1626),
.B(n_1604),
.C(n_1597),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1640),
.A2(n_1606),
.B1(n_1605),
.B2(n_1599),
.C(n_1587),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1638),
.A2(n_1577),
.B1(n_1606),
.B2(n_1605),
.C(n_1596),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1645),
.A2(n_1601),
.B1(n_1596),
.B2(n_1579),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1586),
.C(n_1578),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1644),
.A2(n_1579),
.B(n_1607),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1645),
.A2(n_1601),
.B1(n_1579),
.B2(n_1602),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1659),
.B(n_1647),
.C(n_1655),
.Y(n_1671)
);

NAND4xp75_ASAP7_75t_L g1672 ( 
.A(n_1660),
.B(n_1647),
.C(n_1643),
.D(n_1642),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1661),
.B(n_1656),
.Y(n_1673)
);

NOR4xp75_ASAP7_75t_L g1674 ( 
.A(n_1666),
.B(n_1639),
.C(n_1643),
.D(n_1642),
.Y(n_1674)
);

NAND5xp2_ASAP7_75t_L g1675 ( 
.A(n_1662),
.B(n_1639),
.C(n_1657),
.D(n_1658),
.E(n_1654),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1668),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1664),
.A2(n_1653),
.B(n_1658),
.C(n_1654),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1669),
.B(n_1653),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1665),
.Y(n_1679)
);

AOI322xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1667),
.A3(n_1670),
.B1(n_1663),
.B2(n_1602),
.C1(n_1607),
.C2(n_1608),
.Y(n_1680)
);

OR3x1_ASAP7_75t_L g1681 ( 
.A(n_1675),
.B(n_1579),
.C(n_1510),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1677),
.B(n_1586),
.C(n_1578),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1678),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1673),
.B(n_1607),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1681),
.A2(n_1672),
.B1(n_1676),
.B2(n_1671),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1683),
.A2(n_1682),
.B1(n_1684),
.B2(n_1674),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1680),
.A2(n_1602),
.B1(n_1586),
.B2(n_1588),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_L g1688 ( 
.A(n_1683),
.B(n_1325),
.C(n_1267),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1682),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1681),
.A2(n_1588),
.B1(n_1593),
.B2(n_1578),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1688),
.B(n_1608),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1267),
.C(n_1251),
.Y(n_1692)
);

XNOR2x1_ASAP7_75t_L g1693 ( 
.A(n_1686),
.B(n_1293),
.Y(n_1693)
);

NAND5xp2_ASAP7_75t_L g1694 ( 
.A(n_1689),
.B(n_1254),
.C(n_1293),
.D(n_1570),
.E(n_1571),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1687),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_L g1696 ( 
.A(n_1693),
.B(n_1588),
.Y(n_1696)
);

XOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1254),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1691),
.Y(n_1698)
);

XOR2xp5_ASAP7_75t_L g1699 ( 
.A(n_1697),
.B(n_1690),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1692),
.B1(n_1698),
.B2(n_1694),
.C(n_1696),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1593),
.B1(n_1694),
.B2(n_1611),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1700),
.A2(n_1593),
.B(n_1611),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1701),
.A2(n_1611),
.B1(n_1254),
.B2(n_1512),
.Y(n_1703)
);

AO21x2_ASAP7_75t_L g1704 ( 
.A1(n_1702),
.A2(n_1611),
.B(n_1508),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1704),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1703),
.A2(n_1508),
.B(n_1504),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1705),
.B(n_1313),
.C(n_1504),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1706),
.B1(n_1508),
.B2(n_1525),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1525),
.B1(n_1523),
.B2(n_1512),
.C(n_1510),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1525),
.B(n_1523),
.C(n_1512),
.Y(n_1710)
);


endmodule