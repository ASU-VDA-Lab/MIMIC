module fake_jpeg_10928_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx8_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_53),
.Y(n_107)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_81),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_23),
.Y(n_71)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_75),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_87),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_27),
.B(n_5),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_84),
.Y(n_138)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_27),
.A2(n_35),
.B(n_33),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_36),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_29),
.B(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_92),
.Y(n_137)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_36),
.B1(n_42),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_122),
.B1(n_133),
.B2(n_135),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_111),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_30),
.Y(n_111)
);

BUFx2_ASAP7_75t_R g113 ( 
.A(n_49),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_51),
.B(n_38),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_142),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_50),
.A2(n_42),
.B1(n_32),
.B2(n_46),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_35),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_38),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_20),
.B1(n_32),
.B2(n_46),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_20),
.B1(n_45),
.B2(n_18),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_84),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_69),
.B1(n_60),
.B2(n_80),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_167),
.B1(n_173),
.B2(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_146),
.B(n_149),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_104),
.C(n_110),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.B(n_171),
.CI(n_112),
.CON(n_195),
.SN(n_195)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_150),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_19),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_45),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_155),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_37),
.B(n_19),
.Y(n_153)
);

NOR2x1_ASAP7_75t_R g186 ( 
.A(n_153),
.B(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_37),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_73),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_73),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_166),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_91),
.B1(n_85),
.B2(n_66),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_178),
.B1(n_135),
.B2(n_122),
.Y(n_183)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_77),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_65),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_106),
.A2(n_65),
.B1(n_63),
.B2(n_105),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_52),
.C(n_78),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_97),
.A2(n_63),
.B1(n_78),
.B2(n_72),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_89),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_130),
.B(n_112),
.Y(n_188)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_156),
.B1(n_112),
.B2(n_103),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_102),
.B(n_6),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_114),
.B1(n_117),
.B2(n_98),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_96),
.B1(n_176),
.B2(n_145),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_200),
.B1(n_165),
.B2(n_138),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_159),
.B1(n_139),
.B2(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_163),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_139),
.A3(n_128),
.B1(n_138),
.B2(n_130),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_114),
.B1(n_117),
.B2(n_98),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

CKINVDCx11_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_163),
.B(n_166),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_222),
.B(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_219),
.B1(n_159),
.B2(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_218),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_184),
.B1(n_175),
.B2(n_145),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_221),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_147),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_165),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_195),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_233),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_212),
.B(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_182),
.B1(n_195),
.B2(n_145),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_175),
.B1(n_201),
.B2(n_193),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_155),
.C(n_171),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_207),
.C(n_204),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_186),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_238),
.B1(n_213),
.B2(n_181),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_202),
.B1(n_213),
.B2(n_199),
.Y(n_245)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_186),
.A3(n_184),
.B1(n_187),
.B2(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_211),
.B1(n_222),
.B2(n_215),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_244),
.C(n_232),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_243),
.B(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_249),
.B1(n_230),
.B2(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_198),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_263),
.B1(n_264),
.B2(n_248),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_226),
.C(n_228),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_223),
.C(n_224),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_267),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_234),
.B1(n_223),
.B2(n_233),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_234),
.B1(n_239),
.B2(n_238),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_262),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_251),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_257),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_278),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_245),
.B1(n_242),
.B2(n_235),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_241),
.B1(n_252),
.B2(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_282),
.Y(n_294)
);

BUFx12f_ASAP7_75t_SL g280 ( 
.A(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_281),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_259),
.C(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_201),
.C(n_198),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_287),
.B1(n_268),
.B2(n_202),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_199),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_277),
.CI(n_8),
.CON(n_289),
.SN(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_164),
.B1(n_162),
.B2(n_172),
.Y(n_290)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_119),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_286),
.C(n_287),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_284),
.C(n_127),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_300),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_158),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_289),
.B(n_99),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_304),
.B(n_299),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_99),
.B(n_128),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_308),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_11),
.C(n_12),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_11),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_13),
.Y(n_314)
);


endmodule