module real_jpeg_13291_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_5),
.A2(n_18),
.B(n_19),
.C(n_25),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_5),
.B(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_32),
.C(n_54),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_69),
.B(n_71),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_65)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_73),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_62),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_62),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_39),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_27),
.Y(n_16)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_18),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_18),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_21),
.B(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_21),
.B(n_28),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_22),
.A2(n_23),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_23),
.B(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B(n_35),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_28),
.A2(n_35),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_29),
.B(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_29),
.A2(n_36),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_32),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_31),
.B(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_46),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2x1_ASAP7_75t_R g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_57),
.B2(n_59),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_56),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_65),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.C(n_68),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_86),
.B(n_104),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_83),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_94),
.B(n_103),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_92),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_98),
.B(n_102),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);


endmodule