module fake_jpeg_7390_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_18),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_59),
.C(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_55),
.B1(n_17),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_22),
.B1(n_18),
.B2(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_60),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_22),
.B1(n_24),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_64),
.B1(n_33),
.B2(n_20),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_33),
.B1(n_28),
.B2(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_84),
.B1(n_88),
.B2(n_30),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_86),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_28),
.B1(n_20),
.B2(n_21),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_34),
.B1(n_65),
.B2(n_31),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_90),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_21),
.B1(n_30),
.B2(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_13),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_23),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_34),
.B1(n_29),
.B2(n_26),
.Y(n_146)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_97),
.B(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_104),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_45),
.B(n_59),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_110),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_114),
.B1(n_71),
.B2(n_79),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_65),
.B1(n_47),
.B2(n_51),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_119),
.B1(n_74),
.B2(n_68),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_51),
.B(n_67),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_56),
.B(n_27),
.C(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_117),
.B1(n_94),
.B2(n_101),
.Y(n_147)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_10),
.Y(n_149)
);

OAI22x1_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_23),
.B1(n_31),
.B2(n_46),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_60),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_129),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_134),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_132),
.B1(n_147),
.B2(n_94),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_0),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_136),
.B(n_110),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_78),
.B1(n_70),
.B2(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_130),
.B1(n_137),
.B2(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_68),
.B1(n_86),
.B2(n_90),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_0),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_29),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_113),
.B1(n_111),
.B2(n_118),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_70),
.B1(n_34),
.B2(n_29),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_95),
.B1(n_98),
.B2(n_109),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_26),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_149),
.C(n_96),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_126),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_116),
.C(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_157),
.C(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_163),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_99),
.C(n_100),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_118),
.A3(n_110),
.B1(n_95),
.B2(n_109),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_167),
.B(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_169),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_119),
.C(n_110),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_143),
.B(n_139),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_109),
.B1(n_29),
.B2(n_26),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_178),
.B1(n_129),
.B2(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_26),
.B1(n_29),
.B2(n_1),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_131),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_181),
.B(n_198),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_186),
.B(n_189),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_183),
.A2(n_197),
.B1(n_204),
.B2(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_194),
.B1(n_172),
.B2(n_180),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_137),
.B(n_121),
.Y(n_186)
);

XOR2x1_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_207),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_126),
.B1(n_139),
.B2(n_144),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_151),
.B(n_149),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_135),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_2),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_159),
.C(n_160),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_212),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_153),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_221),
.C(n_224),
.Y(n_252)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_222),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_217),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_172),
.B1(n_152),
.B2(n_168),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_174),
.C(n_179),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_170),
.B(n_150),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_197),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_186),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_159),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_199),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_176),
.B1(n_173),
.B2(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_247),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_198),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_209),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_197),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_214),
.B1(n_226),
.B2(n_221),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_216),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g254 ( 
.A(n_252),
.B(n_216),
.C(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_236),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_224),
.C(n_208),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_238),
.Y(n_269)
);

NOR4xp25_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_203),
.C(n_208),
.D(n_231),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_4),
.C(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_4),
.C(n_6),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_6),
.C(n_7),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_6),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_276),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_255),
.B1(n_233),
.B2(n_259),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_253),
.A2(n_249),
.B(n_240),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_241),
.B(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_236),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_267),
.Y(n_284)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_283),
.B(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_286),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_287),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_250),
.B1(n_244),
.B2(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_266),
.C(n_237),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_260),
.B1(n_8),
.B2(n_9),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_7),
.Y(n_296)
);

OAI21x1_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_298),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_290),
.Y(n_300)
);

NOR2x1_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_273),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_8),
.B(n_10),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_283),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.C(n_296),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_288),
.C(n_13),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_307),
.A2(n_302),
.B(n_295),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_306),
.B(n_308),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_12),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_12),
.Y(n_313)
);


endmodule