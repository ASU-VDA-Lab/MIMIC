module fake_jpeg_31798_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_58),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_61),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_25),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_25),
.B(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_66),
.B(n_70),
.Y(n_158)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_15),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_74),
.B(n_77),
.Y(n_160)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_89),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_42),
.Y(n_138)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_101),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_39),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_108),
.B(n_138),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_48),
.B1(n_39),
.B2(n_43),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_128),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_42),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_119),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_24),
.B1(n_49),
.B2(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_116),
.A2(n_146),
.B1(n_122),
.B2(n_164),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_60),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_24),
.B1(n_49),
.B2(n_22),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_120),
.A2(n_24),
.B1(n_49),
.B2(n_62),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_46),
.B1(n_49),
.B2(n_24),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_71),
.B(n_67),
.Y(n_171)
);

AND2x4_ASAP7_75t_SL g128 ( 
.A(n_66),
.B(n_46),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_43),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_46),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_53),
.A2(n_49),
.B1(n_24),
.B2(n_19),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_151),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_68),
.A2(n_48),
.B(n_19),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_174),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_171),
.A2(n_116),
.B(n_120),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_34),
.B1(n_19),
.B2(n_28),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_173),
.B(n_178),
.Y(n_242)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_180),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_185),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_131),
.B(n_34),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_34),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_188),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_189),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_47),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_203),
.Y(n_243)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx5_ASAP7_75t_SL g268 ( 
.A(n_193),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_123),
.A2(n_124),
.B1(n_75),
.B2(n_127),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_195),
.B1(n_225),
.B2(n_226),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_89),
.B1(n_24),
.B2(n_49),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_196),
.A2(n_210),
.B1(n_216),
.B2(n_224),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_128),
.B(n_83),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_202),
.Y(n_253)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_91),
.B1(n_92),
.B2(n_85),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_212),
.Y(n_259)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_28),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_211),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_133),
.A2(n_59),
.B1(n_56),
.B2(n_80),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_141),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_214),
.Y(n_252)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_51),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_219),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_150),
.A2(n_69),
.B1(n_102),
.B2(n_104),
.Y(n_216)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_145),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_110),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

CKINVDCx12_ASAP7_75t_R g256 ( 
.A(n_221),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_137),
.B(n_51),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_30),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_150),
.A2(n_26),
.B1(n_47),
.B2(n_38),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_118),
.B1(n_166),
.B2(n_159),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_227),
.A2(n_225),
.B1(n_191),
.B2(n_189),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_125),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_172),
.B(n_38),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_217),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_164),
.B1(n_118),
.B2(n_122),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_198),
.B(n_9),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_202),
.B(n_9),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_155),
.B1(n_89),
.B2(n_146),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_249),
.A2(n_261),
.B1(n_269),
.B2(n_211),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_0),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_173),
.B(n_13),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_258),
.B(n_11),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_179),
.A2(n_144),
.B1(n_134),
.B2(n_26),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_177),
.B(n_199),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_199),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_177),
.A2(n_135),
.B1(n_126),
.B2(n_36),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_192),
.B1(n_175),
.B2(n_193),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_187),
.A2(n_135),
.B1(n_36),
.B2(n_32),
.Y(n_269)
);

CKINVDCx12_ASAP7_75t_R g270 ( 
.A(n_183),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_270),
.Y(n_295)
);

AO22x2_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_259),
.B1(n_253),
.B2(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_279),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_168),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_280),
.B(n_256),
.Y(n_353)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_171),
.B(n_218),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_282),
.A2(n_264),
.B(n_252),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_283),
.A2(n_315),
.B(n_264),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g284 ( 
.A1(n_231),
.A2(n_204),
.B(n_195),
.C(n_214),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_284),
.A2(n_277),
.B(n_282),
.Y(n_344)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_296),
.B1(n_307),
.B2(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_169),
.B1(n_207),
.B2(n_200),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_291),
.B1(n_310),
.B2(n_266),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_205),
.B1(n_184),
.B2(n_182),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_230),
.B(n_36),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_292),
.B(n_312),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_245),
.A2(n_201),
.B1(n_220),
.B2(n_32),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_293),
.A2(n_300),
.B1(n_303),
.B2(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_298),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_253),
.A2(n_263),
.B1(n_235),
.B2(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_32),
.B1(n_21),
.B2(n_11),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_228),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_259),
.A2(n_242),
.B1(n_235),
.B2(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_271),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_242),
.A2(n_21),
.B1(n_10),
.B2(n_46),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_243),
.A2(n_21),
.B1(n_46),
.B2(n_51),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_10),
.B1(n_46),
.B2(n_2),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_308),
.A2(n_268),
.B1(n_251),
.B2(n_232),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_229),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_311),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_268),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_51),
.Y(n_312)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_258),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_232),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_243),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_257),
.B1(n_273),
.B2(n_251),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_341),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_318),
.B(n_340),
.Y(n_377)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_247),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_328),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_296),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_272),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_335),
.Y(n_374)
);

OAI22x1_ASAP7_75t_SL g334 ( 
.A1(n_278),
.A2(n_239),
.B1(n_256),
.B2(n_272),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_347),
.B1(n_288),
.B2(n_306),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_230),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_275),
.B(n_228),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_299),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_350),
.B1(n_287),
.B2(n_314),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_346),
.A2(n_349),
.B(n_352),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_277),
.A2(n_264),
.B1(n_252),
.B2(n_257),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_348),
.A2(n_300),
.B1(n_295),
.B2(n_311),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_246),
.B(n_233),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_303),
.A2(n_274),
.B1(n_246),
.B2(n_260),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_316),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_278),
.A2(n_285),
.B(n_281),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_334),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_280),
.B(n_278),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_354),
.A2(n_382),
.B(n_320),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_358),
.A2(n_371),
.B1(n_387),
.B2(n_347),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_278),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_378),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_348),
.Y(n_392)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_376),
.B1(n_343),
.B2(n_329),
.Y(n_404)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_380),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_308),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_385),
.C(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_284),
.B1(n_275),
.B2(n_313),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_373),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_307),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_379),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_338),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_346),
.A2(n_302),
.B(n_295),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_381),
.A2(n_339),
.B(n_351),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_297),
.B(n_289),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_386),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_350),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_274),
.B1(n_255),
.B2(n_260),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_389),
.A2(n_364),
.B(n_375),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_376),
.B1(n_369),
.B2(n_378),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_327),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_392),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_333),
.Y(n_393)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_361),
.Y(n_396)
);

INVx13_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_319),
.Y(n_397)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_377),
.B(n_340),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_402),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_415),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_372),
.Y(n_402)
);

OA21x2_ASAP7_75t_L g403 ( 
.A1(n_355),
.A2(n_319),
.B(n_321),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_358),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_407),
.B1(n_409),
.B2(n_371),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_321),
.Y(n_405)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_365),
.A2(n_351),
.B(n_349),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_418),
.B(n_357),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_372),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_357),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_359),
.B(n_320),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_412),
.A2(n_354),
.B(n_382),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_335),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_365),
.A2(n_329),
.B(n_331),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_439),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_420),
.A2(n_441),
.B1(n_414),
.B2(n_400),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_423),
.B(n_436),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_434),
.Y(n_459)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_412),
.A2(n_364),
.B(n_375),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_433),
.B(n_437),
.Y(n_446)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_362),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_438),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_SL g439 ( 
.A(n_393),
.B(n_325),
.C(n_384),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_389),
.A2(n_387),
.B(n_373),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_403),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_390),
.A2(n_325),
.B1(n_341),
.B2(n_317),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_443),
.A2(n_417),
.B1(n_416),
.B2(n_400),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_392),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_449),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_399),
.C(n_410),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_452),
.C(n_460),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_428),
.A2(n_404),
.B1(n_414),
.B2(n_388),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_401),
.C(n_415),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_432),
.B1(n_424),
.B2(n_430),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_454),
.A2(n_463),
.B1(n_465),
.B2(n_440),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_466),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_401),
.C(n_421),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_426),
.A2(n_400),
.B1(n_418),
.B2(n_391),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_441),
.A2(n_417),
.B1(n_411),
.B2(n_318),
.Y(n_464)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_464),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_403),
.B1(n_406),
.B2(n_337),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_465),
.B(n_463),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_455),
.B(n_454),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_337),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_451),
.A2(n_420),
.B1(n_436),
.B2(n_422),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_466),
.B1(n_446),
.B2(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

OAI21xp33_ASAP7_75t_SL g475 ( 
.A1(n_450),
.A2(n_421),
.B(n_438),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_475),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_342),
.Y(n_476)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_433),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_479),
.C(n_255),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_443),
.C(n_437),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_480),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_429),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_481),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_453),
.A2(n_439),
.B1(n_381),
.B2(n_423),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_482),
.A2(n_483),
.B1(n_233),
.B2(n_304),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_449),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_490),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_487),
.Y(n_500)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_452),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_479),
.A2(n_445),
.B(n_429),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_495),
.B(n_496),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_494),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_301),
.C(n_274),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_273),
.C(n_266),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_484),
.A2(n_473),
.B1(n_468),
.B2(n_467),
.Y(n_502)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_477),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_494),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_472),
.B(n_470),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_506),
.Y(n_516)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_491),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_471),
.B1(n_470),
.B2(n_273),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_507),
.A2(n_489),
.B1(n_493),
.B2(n_266),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_486),
.A2(n_266),
.B(n_240),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_238),
.Y(n_518)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_497),
.C(n_498),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_496),
.C(n_487),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_512),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_513),
.A2(n_518),
.B(n_509),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_515),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_505),
.A2(n_238),
.B1(n_240),
.B2(n_5),
.Y(n_515)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_519),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_499),
.B(n_508),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_523),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_516),
.B(n_501),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_SL g524 ( 
.A1(n_521),
.A2(n_517),
.B(n_518),
.C(n_501),
.Y(n_524)
);

OAI221xp5_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_526),
.B1(n_507),
.B2(n_240),
.C(n_238),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_522),
.Y(n_527)
);

OAI311xp33_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.A3(n_1),
.B1(n_4),
.C1(n_5),
.Y(n_529)
);

OA21x2_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_7),
.B(n_8),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_7),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_7),
.B(n_8),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_8),
.C(n_402),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_533),
.Y(n_534)
);


endmodule