module fake_jpeg_11497_n_144 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx9p33_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_32),
.B(n_35),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_6),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_38),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_4),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_40),
.B(n_46),
.Y(n_86)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_5),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_12),
.B(n_5),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_58),
.Y(n_83)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_12),
.A2(n_5),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_21),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_16),
.B1(n_11),
.B2(n_30),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_70),
.B(n_79),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_16),
.B1(n_11),
.B2(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_59),
.B1(n_33),
.B2(n_55),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_31),
.B1(n_34),
.B2(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_78),
.B1(n_75),
.B2(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_47),
.B1(n_37),
.B2(n_44),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_56),
.B(n_57),
.C(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_96),
.Y(n_115)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_79),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_85),
.B1(n_74),
.B2(n_80),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_103),
.B(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_102),
.B(n_105),
.Y(n_110)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_83),
.B(n_60),
.C(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_117),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_104),
.B1(n_99),
.B2(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_69),
.C(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_74),
.B1(n_85),
.B2(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_121),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_106),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_124),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_93),
.B(n_100),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_93),
.C(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_106),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_129),
.B1(n_117),
.B2(n_116),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_112),
.B1(n_115),
.B2(n_113),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_125),
.B1(n_121),
.B2(n_109),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_125),
.B1(n_114),
.B2(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_134),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_129),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_108),
.A3(n_116),
.B1(n_80),
.B2(n_67),
.C(n_101),
.Y(n_134)
);

OAI31xp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_127),
.A3(n_67),
.B(n_105),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_131),
.A3(n_127),
.B1(n_133),
.B2(n_89),
.C1(n_67),
.C2(n_108),
.Y(n_138)
);

OAI31xp33_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_139),
.A3(n_135),
.B(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_140),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);


endmodule