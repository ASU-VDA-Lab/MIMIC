module real_aes_1359_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
HB1xp67_ASAP7_75t_L g6 ( .A(n_0), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g9 ( .A(n_3), .B(n_7), .Y(n_9) );
AOI32xp33_ASAP7_75t_L g4 ( .A1(n_5), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .Y(n_4) );
CKINVDCx20_ASAP7_75t_R g5 ( .A(n_6), .Y(n_5) );
endmodule