module fake_jpeg_2896_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_13),
.C(n_28),
.Y(n_43)
);

NAND2x1_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_47),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_56),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_38),
.B1(n_34),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_42),
.B1(n_45),
.B2(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_34),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_31),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_70),
.B(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_45),
.B1(n_32),
.B2(n_39),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_57),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_31),
.B1(n_30),
.B2(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_6),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_48),
.B(n_16),
.C(n_17),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_58),
.B1(n_57),
.B2(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_81),
.B1(n_63),
.B2(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_6),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_10),
.B(n_11),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_15),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_79),
.B1(n_81),
.B2(n_71),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_20),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_12),
.B1(n_25),
.B2(n_27),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_97),
.B(n_101),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_86),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_96),
.Y(n_109)
);

AOI321xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_106),
.A3(n_99),
.B1(n_91),
.B2(n_95),
.C(n_104),
.Y(n_110)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_98),
.A3(n_90),
.B1(n_102),
.B2(n_88),
.C(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_83),
.Y(n_112)
);


endmodule