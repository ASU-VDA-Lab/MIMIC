module real_jpeg_23373_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_SL g85 ( 
.A(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_6),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_8),
.B(n_39),
.C(n_65),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_8),
.B(n_55),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_8),
.A2(n_36),
.B1(n_136),
.B2(n_139),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_57),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_104),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_103),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_71),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_18),
.B(n_71),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_51),
.C(n_58),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_19),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_34),
.B2(n_35),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B(n_27),
.C(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_22),
.A2(n_23),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.CON(n_28),
.SN(n_28)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_29),
.A2(n_33),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_31),
.B(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_31),
.B(n_41),
.Y(n_141)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_42),
.B(n_44),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_36),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_36),
.A2(n_48),
.B1(n_129),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_37),
.B(n_45),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_37),
.A2(n_118),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_38),
.B(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_40),
.Y(n_139)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_42),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_50),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_51),
.B(n_58),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_60),
.A2(n_63),
.B1(n_67),
.B2(n_113),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_68),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_94),
.B2(n_95),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_87),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_93),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_145),
.B(n_149),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_125),
.B(n_144),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_110),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_121),
.C(n_124),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_132),
.B(n_143),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_131),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_137),
.B(n_142),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_148),
.Y(n_149)
);


endmodule