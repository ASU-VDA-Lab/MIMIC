module fake_jpeg_1569_n_578 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_578);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g177 ( 
.A(n_59),
.Y(n_177)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_61),
.Y(n_185)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_65),
.B(n_107),
.Y(n_158)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_20),
.A2(n_18),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_70),
.B(n_9),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_78),
.Y(n_138)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_77),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_80),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_81),
.Y(n_167)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_93),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_96),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_97),
.B(n_103),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_43),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_38),
.Y(n_104)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_31),
.B(n_18),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_43),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_113),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_45),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_49),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_121),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_51),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_33),
.Y(n_172)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_32),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_14),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_59),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_128),
.A2(n_137),
.B1(n_147),
.B2(n_154),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_62),
.B(n_19),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_130),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_56),
.B1(n_22),
.B2(n_32),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_22),
.B1(n_46),
.B2(n_21),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_66),
.A2(n_50),
.B1(n_46),
.B2(n_21),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_151),
.A2(n_164),
.B1(n_181),
.B2(n_199),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_22),
.B1(n_29),
.B2(n_40),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_91),
.A2(n_50),
.B1(n_40),
.B2(n_35),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_165),
.B(n_192),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_97),
.B(n_35),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_198),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_203),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_74),
.A2(n_26),
.B1(n_19),
.B2(n_45),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_176),
.A2(n_196),
.B1(n_214),
.B2(n_128),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_58),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_124),
.A2(n_23),
.B1(n_26),
.B2(n_19),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_64),
.A2(n_26),
.B1(n_2),
.B2(n_4),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_71),
.A2(n_26),
.B1(n_4),
.B2(n_5),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_72),
.A2(n_26),
.B1(n_17),
.B2(n_16),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_79),
.B(n_17),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_75),
.A2(n_1),
.B1(n_6),
.B2(n_8),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_83),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_103),
.B(n_14),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_80),
.A2(n_1),
.B1(n_6),
.B2(n_8),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_86),
.A2(n_106),
.B1(n_123),
.B2(n_120),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_200),
.A2(n_184),
.B1(n_183),
.B2(n_84),
.Y(n_294)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_101),
.Y(n_206)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_113),
.B(n_110),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_207),
.B(n_210),
.Y(n_268)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_116),
.B(n_6),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_122),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_87),
.B(n_9),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_217),
.B(n_202),
.Y(n_241)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_105),
.C(n_127),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_221),
.B(n_254),
.C(n_291),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_222),
.B(n_232),
.Y(n_315)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_223),
.Y(n_296)
);

NAND2x1_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_110),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_224),
.B(n_241),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_90),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_226),
.B(n_235),
.Y(n_311)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_227),
.Y(n_298)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_228),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_180),
.B1(n_152),
.B2(n_146),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_229),
.A2(n_276),
.B1(n_275),
.B2(n_219),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_93),
.A3(n_95),
.B1(n_108),
.B2(n_10),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_263),
.B(n_282),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_160),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_234),
.A2(n_240),
.B(n_275),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_11),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_167),
.A2(n_11),
.B1(n_174),
.B2(n_175),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_138),
.B(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_242),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_129),
.A2(n_187),
.B1(n_148),
.B2(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_155),
.B(n_143),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_243),
.B(n_278),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_244),
.B(n_246),
.Y(n_319)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_157),
.Y(n_245)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_204),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_159),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_248),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_159),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_130),
.B(n_134),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_256),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_149),
.Y(n_257)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_139),
.Y(n_258)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_135),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

O2A1O1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_183),
.A2(n_184),
.B(n_176),
.C(n_147),
.Y(n_263)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_264),
.Y(n_349)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_137),
.A2(n_193),
.B1(n_189),
.B2(n_179),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_279),
.B1(n_289),
.B2(n_294),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_142),
.Y(n_271)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_163),
.Y(n_272)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_176),
.A2(n_162),
.B1(n_168),
.B2(n_190),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_274),
.A2(n_280),
.B1(n_283),
.B2(n_266),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_195),
.A2(n_201),
.B1(n_132),
.B2(n_150),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_131),
.Y(n_277)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_140),
.A2(n_196),
.B1(n_154),
.B2(n_135),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_178),
.B(n_186),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_161),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_281),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_188),
.A2(n_214),
.B(n_131),
.C(n_203),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_149),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_131),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_284),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_161),
.A2(n_166),
.B1(n_169),
.B2(n_173),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_285),
.A2(n_292),
.B1(n_289),
.B2(n_286),
.Y(n_346)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_290),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g289 ( 
.A1(n_212),
.A2(n_99),
.B1(n_112),
.B2(n_98),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_158),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_146),
.B(n_152),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_183),
.A2(n_184),
.B1(n_210),
.B2(n_180),
.Y(n_292)
);

NOR2x1_ASAP7_75t_R g293 ( 
.A(n_217),
.B(n_202),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_224),
.C(n_269),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_323),
.B1(n_342),
.B2(n_346),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_225),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_302),
.B(n_306),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_291),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_332),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_221),
.B(n_278),
.C(n_293),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_308),
.B(n_326),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_230),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_329),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_263),
.A2(n_278),
.B(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_317),
.A2(n_252),
.B(n_272),
.Y(n_357)
);

OAI22x1_ASAP7_75t_SL g323 ( 
.A1(n_276),
.A2(n_236),
.B1(n_243),
.B2(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_267),
.C(n_273),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_251),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_243),
.B(n_267),
.C(n_262),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_331),
.C(n_341),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_262),
.B(n_236),
.C(n_220),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_236),
.B(n_270),
.C(n_255),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_231),
.A2(n_236),
.B1(n_234),
.B2(n_240),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_312),
.A2(n_223),
.B1(n_245),
.B2(n_285),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_350),
.A2(n_370),
.B1(n_378),
.B2(n_381),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_265),
.B(n_249),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_351),
.A2(n_367),
.B(n_391),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_302),
.B(n_253),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_360),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_315),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_358),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_253),
.B1(n_255),
.B2(n_257),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_356),
.B1(n_363),
.B2(n_368),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_237),
.B1(n_256),
.B2(n_250),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_357),
.A2(n_367),
.B(n_391),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_329),
.B(n_288),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_261),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_374),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_300),
.B(n_328),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_362),
.B(n_382),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_277),
.B1(n_264),
.B2(n_284),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_366),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_347),
.A2(n_228),
.B(n_284),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_228),
.B1(n_305),
.B2(n_297),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_318),
.B1(n_313),
.B2(n_331),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_369),
.A2(n_377),
.B1(n_303),
.B2(n_324),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_305),
.A2(n_347),
.B1(n_346),
.B2(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_347),
.A2(n_295),
.B1(n_306),
.B2(n_312),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g422 ( 
.A1(n_372),
.A2(n_390),
.B(n_351),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_325),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_349),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_380),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_301),
.B1(n_295),
.B2(n_308),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_316),
.A2(n_301),
.B1(n_327),
.B2(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_379),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_298),
.B(n_336),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_309),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_385),
.A2(n_375),
.B1(n_381),
.B2(n_371),
.Y(n_419)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_386),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_340),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_304),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_309),
.B(n_338),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_389),
.Y(n_418)
);

AO22x1_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_304),
.B1(n_296),
.B2(n_345),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_316),
.A2(n_307),
.B(n_299),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_392),
.B(n_414),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_386),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_396),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_386),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_299),
.C(n_314),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_398),
.B(n_424),
.C(n_383),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_364),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_412),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_354),
.A2(n_320),
.B1(n_333),
.B2(n_296),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_405),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_314),
.B(n_337),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_404),
.A2(n_410),
.B(n_417),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_354),
.A2(n_320),
.B1(n_333),
.B2(n_303),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_357),
.A2(n_337),
.B(n_338),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_364),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_358),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_365),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_373),
.A2(n_324),
.B(n_322),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_373),
.B(n_360),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_368),
.A2(n_384),
.B1(n_377),
.B2(n_372),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_390),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_370),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_378),
.Y(n_424)
);

AO21x1_ASAP7_75t_L g469 ( 
.A1(n_426),
.A2(n_429),
.B(n_440),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_402),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_428),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_397),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_422),
.A2(n_373),
.B(n_384),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_393),
.B(n_352),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_442),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_393),
.B(n_376),
.Y(n_433)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_416),
.B(n_376),
.Y(n_436)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_399),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_439),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_369),
.B1(n_355),
.B2(n_356),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_441),
.A2(n_448),
.B1(n_455),
.B2(n_400),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_415),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_423),
.C(n_415),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_399),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_446),
.A2(n_454),
.B1(n_456),
.B2(n_409),
.Y(n_480)
);

AO22x1_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_390),
.B1(n_363),
.B2(n_383),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_447),
.A2(n_426),
.B(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_404),
.B(n_374),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_450),
.B(n_451),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_418),
.B(n_359),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_418),
.B(n_366),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_414),
.B1(n_400),
.B2(n_403),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_466),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_424),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_464),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_398),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_408),
.B1(n_422),
.B2(n_420),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_476),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_470),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_392),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_475),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_423),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_447),
.A2(n_405),
.B1(n_410),
.B2(n_417),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_447),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_478),
.C(n_481),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_447),
.A2(n_407),
.B1(n_394),
.B2(n_396),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_SL g490 ( 
.A(n_479),
.B(n_446),
.C(n_438),
.Y(n_490)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_480),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_409),
.C(n_413),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_432),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_436),
.B(n_413),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_450),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_485),
.B(n_442),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_489),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_490),
.A2(n_502),
.B(n_469),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_460),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_493),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_481),
.B(n_451),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_495),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_444),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_504),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_458),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_498),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_438),
.C(n_426),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_508),
.C(n_475),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_484),
.B(n_462),
.Y(n_501)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_501),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_443),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_433),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_472),
.B(n_443),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_496),
.Y(n_510)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_507),
.A2(n_467),
.B1(n_428),
.B2(n_431),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_SL g508 ( 
.A(n_468),
.B(n_425),
.C(n_454),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_512),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_477),
.Y(n_512)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_513),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_515),
.Y(n_536)
);

MAJx2_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_469),
.C(n_482),
.Y(n_515)
);

BUFx12_ASAP7_75t_L g516 ( 
.A(n_490),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_516),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_517),
.A2(n_486),
.B1(n_499),
.B2(n_483),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_487),
.B(n_479),
.C(n_476),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_525),
.C(n_508),
.Y(n_528)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_522),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_492),
.B(n_458),
.C(n_459),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_504),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_526),
.B(n_528),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_511),
.B(n_474),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_529),
.B(n_531),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_520),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_500),
.C(n_494),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_505),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_538),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_521),
.A2(n_497),
.B1(n_457),
.B2(n_483),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_537),
.A2(n_419),
.B1(n_467),
.B2(n_453),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_517),
.A2(n_497),
.B1(n_480),
.B2(n_425),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_518),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_411),
.Y(n_552)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_465),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_541),
.B(n_551),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_537),
.A2(n_497),
.B1(n_524),
.B2(n_519),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_544),
.B(n_545),
.Y(n_555)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_527),
.B(n_515),
.CI(n_516),
.CON(n_545),
.SN(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_523),
.C(n_514),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_531),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_530),
.A2(n_532),
.B(n_516),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_SL g554 ( 
.A(n_548),
.B(n_543),
.C(n_545),
.Y(n_554)
);

AOI21xp33_ASAP7_75t_L g549 ( 
.A1(n_536),
.A2(n_453),
.B(n_470),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_549),
.A2(n_536),
.B(n_489),
.Y(n_558)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_379),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_547),
.C(n_542),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_554),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_540),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_556),
.A2(n_558),
.B(n_548),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_557),
.B(n_560),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_562),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_543),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_559),
.B(n_541),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_561),
.B(n_535),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_535),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_568),
.A2(n_456),
.B(n_430),
.Y(n_571)
);

AOI321xp33_ASAP7_75t_SL g569 ( 
.A1(n_565),
.A2(n_545),
.A3(n_555),
.B1(n_538),
.B2(n_510),
.C(n_533),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_569),
.B(n_571),
.C(n_572),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_568),
.A2(n_550),
.B(n_533),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_567),
.C(n_523),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_512),
.B1(n_427),
.B2(n_494),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_575),
.A2(n_573),
.B(n_473),
.Y(n_576)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_452),
.B(n_449),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_455),
.Y(n_578)
);


endmodule