module fake_jpeg_20411_n_261 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_20),
.B(n_28),
.Y(n_38)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_35),
.B1(n_30),
.B2(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_16),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_47),
.B(n_60),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_58),
.C(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_57),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_37),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_35),
.B1(n_27),
.B2(n_23),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_19),
.B1(n_34),
.B2(n_20),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_31),
.B1(n_34),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_40),
.B1(n_42),
.B2(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_86),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_61),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_77),
.B1(n_105),
.B2(n_61),
.Y(n_115)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_40),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_37),
.C(n_41),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_102),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_98),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_33),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_37),
.A3(n_21),
.B1(n_32),
.B2(n_24),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_68),
.B(n_67),
.C(n_50),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_33),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_7),
.B(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_51),
.B(n_48),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_113),
.B(n_81),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_117),
.B1(n_124),
.B2(n_79),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_61),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_119),
.B1(n_120),
.B2(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_41),
.B1(n_36),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_26),
.B1(n_36),
.B2(n_32),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_41),
.B1(n_36),
.B2(n_26),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_75),
.A2(n_33),
.B1(n_21),
.B2(n_24),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_17),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_17),
.B1(n_32),
.B2(n_24),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_83),
.B1(n_91),
.B2(n_86),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_33),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_17),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_93),
.B1(n_88),
.B2(n_3),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_156),
.B(n_108),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_76),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_148),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_102),
.C(n_89),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_113),
.C(n_110),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_112),
.B1(n_117),
.B2(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_111),
.B(n_12),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_159),
.C(n_161),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_96),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_125),
.B1(n_123),
.B2(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_79),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_71),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_114),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_158),
.B1(n_139),
.B2(n_144),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_130),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_172),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_132),
.C(n_108),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_156),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_113),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_113),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_174),
.B(n_137),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_106),
.C(n_120),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_125),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_182),
.B1(n_153),
.B2(n_157),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_190),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_191),
.A2(n_197),
.B1(n_199),
.B2(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

AO21x2_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_141),
.B(n_146),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_171),
.B1(n_155),
.B2(n_72),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_173),
.B(n_184),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_198),
.B(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_149),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_147),
.B1(n_139),
.B2(n_143),
.C(n_152),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_203),
.B1(n_159),
.B2(n_165),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_136),
.C(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_177),
.C(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_175),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_208),
.B1(n_191),
.B2(n_190),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_193),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_181),
.B1(n_178),
.B2(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_211),
.C(n_202),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_171),
.C(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_196),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_72),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_155),
.C(n_4),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_201),
.C(n_4),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_187),
.B(n_198),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_231),
.B(n_212),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_228),
.C(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_195),
.C(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_215),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_234),
.B(n_241),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_212),
.B1(n_213),
.B2(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_193),
.B1(n_186),
.B2(n_222),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_9),
.B(n_5),
.Y(n_247)
);

OAI221xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_205),
.B1(n_207),
.B2(n_230),
.C(n_221),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_243),
.B(n_247),
.Y(n_250)
);

OAI221xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_204),
.B1(n_222),
.B2(n_227),
.C(n_193),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_237),
.B1(n_238),
.B2(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_9),
.C(n_5),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_239),
.C(n_6),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_6),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_15),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_246),
.C(n_8),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_250),
.C(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

OAI211xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_15),
.B(n_13),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_256),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_258),
.B(n_0),
.Y(n_261)
);


endmodule