module fake_aes_7953_n_748 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_748);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_748;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_37), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_11), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_15), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_10), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_10), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_17), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_44), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_58), .Y(n_92) );
BUFx3_ASAP7_75t_L g93 ( .A(n_3), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_24), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_77), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_31), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_72), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_69), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_79), .Y(n_100) );
BUFx2_ASAP7_75t_L g101 ( .A(n_78), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_61), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_11), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_80), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_52), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_13), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_32), .Y(n_112) );
INVxp33_ASAP7_75t_L g113 ( .A(n_47), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_50), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_9), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_35), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_45), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_9), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_41), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_34), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_6), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_65), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_7), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
INVxp33_ASAP7_75t_SL g128 ( .A(n_13), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_5), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_73), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_21), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_40), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_101), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
XNOR2x2_ASAP7_75t_L g137 ( .A(n_88), .B(n_1), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_93), .B(n_1), .Y(n_142) );
BUFx8_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_113), .B(n_2), .Y(n_144) );
BUFx12f_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_93), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_109), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_148) );
INVx5_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_109), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
BUFx8_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_89), .B(n_8), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_123), .B(n_8), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_121), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_95), .B(n_53), .Y(n_159) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_96), .A2(n_54), .B(n_81), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_123), .B(n_12), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_128), .A2(n_14), .B1(n_19), .B2(n_20), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_97), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_102), .A2(n_55), .B(n_23), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_104), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_105), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_103), .B(n_14), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g171 ( .A1(n_128), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_112), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_114), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_110), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_116), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_120), .B(n_28), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_127), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_177), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g187 ( .A(n_154), .B(n_117), .C(n_131), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_161), .B(n_134), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_142), .B(n_134), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_161), .B(n_84), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_161), .B(n_132), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_144), .B(n_132), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_169), .B(n_92), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_177), .B(n_92), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
AND3x1_ASAP7_75t_L g200 ( .A(n_163), .B(n_130), .C(n_121), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_162), .B(n_126), .C(n_108), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
INVx5_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_144), .B(n_179), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_175), .B(n_126), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_142), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_169), .B(n_107), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_142), .B(n_130), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_173), .B(n_122), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_115), .B1(n_111), .B2(n_100), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_153), .B(n_99), .C(n_98), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_179), .B(n_94), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_142), .B(n_30), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_173), .B(n_36), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_149), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_177), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_177), .Y(n_228) );
AND2x4_ASAP7_75t_SL g229 ( .A(n_170), .B(n_38), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_143), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_175), .B(n_39), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_176), .B(n_42), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_176), .B(n_46), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_145), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_136), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_147), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_139), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_177), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_174), .B(n_48), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_174), .B(n_49), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_180), .B(n_56), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_140), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_159), .A2(n_57), .B1(n_59), .B2(n_60), .Y(n_246) );
INVx4_ASAP7_75t_L g247 ( .A(n_159), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_140), .Y(n_248) );
AND2x6_ASAP7_75t_SL g249 ( .A(n_211), .B(n_137), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
NAND2x1_ASAP7_75t_L g251 ( .A(n_217), .B(n_159), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_206), .B(n_155), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_206), .B(n_180), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_216), .B(n_177), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_182), .B(n_178), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_216), .B(n_172), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_195), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_135), .B1(n_163), .B2(n_171), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_230), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_211), .A2(n_150), .B1(n_148), .B2(n_155), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_L g261 ( .A1(n_182), .A2(n_146), .B(n_167), .C(n_158), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_233), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_237), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_195), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_208), .B(n_146), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_235), .B(n_172), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_209), .A2(n_167), .B1(n_151), .B2(n_158), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_192), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_235), .B(n_151), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_192), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_240), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_196), .B(n_143), .Y(n_274) );
BUFx6f_ASAP7_75t_SL g275 ( .A(n_192), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_188), .B(n_240), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_187), .A2(n_150), .B1(n_141), .B2(n_165), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_229), .B(n_157), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_182), .B(n_143), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_191), .B(n_143), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_229), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
NAND2x1_ASAP7_75t_L g284 ( .A(n_217), .B(n_141), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_194), .B(n_152), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_230), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_224), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_186), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_210), .B(n_152), .Y(n_289) );
NOR3xp33_ASAP7_75t_L g290 ( .A(n_203), .B(n_157), .C(n_168), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_209), .A2(n_137), .B1(n_168), .B2(n_165), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_186), .B(n_152), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_183), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_190), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_209), .A2(n_156), .B1(n_157), .B2(n_160), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_215), .B(n_156), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_212), .B(n_152), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_217), .B(n_62), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_193), .B(n_166), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_199), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_214), .B(n_166), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_225), .A2(n_160), .B1(n_166), .B2(n_66), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_225), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_197), .B(n_166), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_236), .A2(n_160), .B1(n_64), .B2(n_67), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_244), .B(n_63), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_244), .B(n_68), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_236), .B(n_70), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_238), .B(n_82), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_239), .A2(n_75), .B1(n_76), .B2(n_248), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_245), .B(n_248), .Y(n_315) );
AO22x1_ASAP7_75t_L g316 ( .A1(n_200), .A2(n_247), .B1(n_199), .B2(n_205), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_199), .B(n_247), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_205), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_245), .B(n_239), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_245), .B(n_205), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_247), .B(n_205), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_242), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_275), .Y(n_323) );
INVx11_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_270), .A2(n_219), .B(n_234), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_257), .A2(n_227), .B1(n_232), .B2(n_205), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_288), .B(n_231), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_300), .A2(n_200), .B1(n_246), .B2(n_227), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_251), .A2(n_227), .B(n_241), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_265), .B(n_226), .Y(n_331) );
O2A1O1Ixp5_ASAP7_75t_L g332 ( .A1(n_303), .A2(n_243), .B(n_218), .C(n_222), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_288), .B(n_241), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_282), .B(n_228), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_312), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_301), .A2(n_227), .B(n_228), .Y(n_338) );
AO22x1_ASAP7_75t_L g339 ( .A1(n_300), .A2(n_227), .B1(n_226), .B2(n_185), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_277), .B(n_185), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_250), .Y(n_341) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_279), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_222), .B(n_218), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_252), .B(n_204), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_255), .A2(n_204), .B(n_223), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_258), .A2(n_202), .B1(n_213), .B2(n_207), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_255), .A2(n_223), .B(n_202), .Y(n_347) );
BUFx4f_ASAP7_75t_L g348 ( .A(n_279), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_253), .B(n_213), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_279), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_300), .A2(n_207), .B1(n_221), .B2(n_220), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_268), .B(n_220), .Y(n_352) );
INVx4_ASAP7_75t_L g353 ( .A(n_288), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_284), .A2(n_181), .B(n_184), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_256), .B(n_220), .Y(n_355) );
INVx6_ASAP7_75t_L g356 ( .A(n_249), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_322), .A2(n_181), .B(n_184), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_271), .B(n_220), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_309), .A2(n_220), .B1(n_221), .B2(n_201), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_189), .B(n_198), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_260), .B(n_221), .Y(n_362) );
O2A1O1Ixp5_ASAP7_75t_L g363 ( .A1(n_303), .A2(n_189), .B(n_198), .C(n_201), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_278), .B(n_221), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_295), .A2(n_221), .B(n_307), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_269), .B(n_266), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_269), .B(n_290), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_261), .A2(n_310), .B(n_267), .C(n_273), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_296), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_291), .A2(n_315), .B(n_319), .C(n_254), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_291), .B(n_316), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_285), .A2(n_274), .B(n_292), .C(n_280), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_283), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_259), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_297), .A2(n_286), .B1(n_305), .B2(n_287), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_317), .B(n_296), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_317), .A2(n_299), .B1(n_289), .B2(n_302), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_321), .A2(n_292), .B(n_280), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_321), .A2(n_317), .B(n_281), .Y(n_379) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_262), .B(n_263), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_262), .B(n_263), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_365), .A2(n_304), .B(n_308), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_372), .A2(n_320), .B(n_302), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_338), .A2(n_304), .B(n_313), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g386 ( .A1(n_365), .A2(n_308), .B(n_264), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_363), .A2(n_311), .B(n_264), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_314), .B(n_293), .C(n_294), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_379), .A2(n_318), .B(n_293), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
AO31x2_ASAP7_75t_L g393 ( .A1(n_368), .A2(n_276), .A3(n_294), .B(n_298), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_362), .B(n_314), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_341), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_361), .B(n_318), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_328), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_329), .A2(n_276), .B1(n_298), .B2(n_318), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_330), .A2(n_378), .B(n_360), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_366), .B(n_364), .C(n_358), .Y(n_402) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_323), .B(n_350), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_377), .A2(n_357), .B(n_351), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_349), .A2(n_352), .B(n_340), .C(n_374), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_332), .A2(n_371), .B(n_346), .C(n_325), .Y(n_406) );
NOR2xp67_ASAP7_75t_SL g407 ( .A(n_336), .B(n_369), .Y(n_407) );
AO21x1_ASAP7_75t_L g408 ( .A1(n_359), .A2(n_327), .B(n_343), .Y(n_408) );
NAND3x1_ASAP7_75t_L g409 ( .A(n_356), .B(n_324), .C(n_375), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_355), .B(n_331), .Y(n_410) );
BUFx2_ASAP7_75t_R g411 ( .A(n_373), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_348), .B(n_353), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_348), .B(n_336), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_345), .A2(n_347), .B(n_339), .Y(n_414) );
AO31x2_ASAP7_75t_L g415 ( .A1(n_354), .A2(n_334), .A3(n_343), .B(n_380), .Y(n_415) );
AOI21x1_ASAP7_75t_SL g416 ( .A1(n_326), .A2(n_333), .B(n_381), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
BUFx12f_ASAP7_75t_L g419 ( .A(n_391), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_389), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_401), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_383), .A2(n_336), .B(n_369), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_385), .A2(n_399), .B(n_383), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_400), .B(n_369), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_414), .A2(n_387), .B(n_416), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_406), .A2(n_394), .B(n_388), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_382), .B(n_392), .Y(n_429) );
OAI21x1_ASAP7_75t_L g430 ( .A1(n_386), .A2(n_404), .B(n_408), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_393), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_410), .B(n_396), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_386), .A2(n_398), .B(n_384), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_415), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_398), .A2(n_402), .B(n_390), .Y(n_438) );
AOI21xp33_ASAP7_75t_SL g439 ( .A1(n_412), .A2(n_403), .B(n_413), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_415), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_405), .A2(n_418), .B(n_397), .Y(n_441) );
OAI21x1_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_415), .B(n_407), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_411), .A2(n_383), .B(n_406), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_417), .A2(n_385), .B(n_399), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_400), .A2(n_260), .B1(n_356), .B2(n_329), .Y(n_445) );
AO31x2_ASAP7_75t_L g446 ( .A1(n_406), .A2(n_408), .A3(n_394), .B(n_404), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_300), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_400), .B(n_206), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_400), .B(n_211), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_440), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_440), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_431), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_433), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_419), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_436), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_431), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_432), .B(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_436), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_442), .B(n_433), .Y(n_460) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_444), .B(n_427), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_421), .Y(n_462) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_424), .A2(n_430), .B(n_427), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_432), .B(n_428), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_447), .B(n_441), .Y(n_466) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_444), .A2(n_430), .B(n_426), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_428), .B(n_447), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_447), .B(n_425), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_425), .B(n_441), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_437), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_434), .Y(n_473) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_430), .A2(n_426), .B(n_435), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_445), .B(n_443), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_442), .B(n_437), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_421), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_443), .B(n_429), .Y(n_481) );
OR2x6_ASAP7_75t_L g482 ( .A(n_442), .B(n_443), .Y(n_482) );
AOI21x1_ASAP7_75t_L g483 ( .A1(n_426), .A2(n_443), .B(n_423), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_419), .B(n_429), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_443), .B(n_429), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_458), .B(n_446), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_455), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_458), .B(n_448), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_476), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_454), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_450), .B(n_446), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_460), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_465), .B(n_446), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_469), .B(n_446), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_469), .B(n_446), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_454), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_450), .B(n_446), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_460), .B(n_419), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_452), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_451), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_451), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_454), .B(n_448), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_456), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_468), .B(n_429), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_456), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_468), .B(n_446), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_475), .B(n_422), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_456), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_466), .B(n_422), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_481), .B(n_422), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_457), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_475), .B(n_438), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_485), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_462), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_464), .B(n_449), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_470), .B(n_439), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_473), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_460), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_471), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_462), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_470), .B(n_439), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_473), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_501), .B(n_466), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_488), .B(n_472), .Y(n_538) );
NAND2x1_ASAP7_75t_L g539 ( .A(n_507), .B(n_460), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_495), .Y(n_540) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_492), .B(n_478), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_487), .B(n_486), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_490), .B(n_479), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_487), .B(n_486), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_511), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_500), .B(n_472), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_493), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_500), .B(n_479), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_481), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_515), .B(n_471), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_502), .B(n_478), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_532), .B(n_482), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_489), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_507), .B(n_478), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_494), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_503), .B(n_480), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_494), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_503), .B(n_461), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_515), .B(n_480), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_532), .B(n_482), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_528), .B(n_461), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_518), .B(n_480), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_509), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_505), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_518), .B(n_473), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_524), .B(n_463), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_520), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_524), .B(n_463), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_522), .B(n_463), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_522), .B(n_463), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_522), .B(n_474), .Y(n_583) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_507), .B(n_482), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_497), .B(n_461), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_522), .B(n_474), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_532), .B(n_491), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_520), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_497), .B(n_474), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_508), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_506), .B(n_474), .Y(n_592) );
NOR2x1p5_ASAP7_75t_L g593 ( .A(n_492), .B(n_483), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_525), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_506), .B(n_484), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_529), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_550), .B(n_533), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_553), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_590), .B(n_533), .Y(n_600) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_593), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_555), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
NOR2x1_ASAP7_75t_L g604 ( .A(n_594), .B(n_507), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_549), .B(n_534), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_545), .B(n_535), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_549), .B(n_534), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_550), .B(n_529), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_590), .B(n_521), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_546), .B(n_517), .Y(n_610) );
NAND2xp67_ASAP7_75t_L g611 ( .A(n_584), .B(n_530), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_538), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_546), .B(n_527), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_560), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_542), .B(n_534), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_551), .B(n_521), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_559), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_548), .B(n_513), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_565), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_571), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_547), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_542), .B(n_504), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_544), .B(n_504), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_584), .B(n_516), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_558), .B(n_499), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_559), .B(n_499), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_592), .B(n_508), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_585), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_539), .B(n_508), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_576), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_570), .A2(n_482), .B1(n_491), .B2(n_526), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_577), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_592), .B(n_536), .Y(n_637) );
AND2x2_ASAP7_75t_SL g638 ( .A(n_570), .B(n_491), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
BUFx12f_ASAP7_75t_L g640 ( .A(n_541), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_538), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_558), .B(n_491), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_564), .B(n_536), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_564), .B(n_536), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_569), .B(n_482), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_563), .B(n_531), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_552), .B(n_531), .Y(n_648) );
OR2x2_ASAP7_75t_SL g649 ( .A(n_585), .B(n_531), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_569), .B(n_512), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_598), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_599), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_641), .B(n_580), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_602), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_603), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_606), .A2(n_567), .B1(n_552), .B2(n_586), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_606), .B(n_543), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_641), .B(n_575), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_614), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_628), .A2(n_541), .B1(n_556), .B2(n_537), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_632), .B(n_575), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_625), .B(n_583), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_600), .B(n_580), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_618), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_617), .Y(n_665) );
AND2x4_ASAP7_75t_SL g666 ( .A(n_626), .B(n_567), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_620), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_621), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_640), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_622), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_632), .B(n_568), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_624), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_612), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_634), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_605), .B(n_583), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_636), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_639), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_597), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_607), .B(n_586), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_608), .Y(n_680) );
OR2x6_ASAP7_75t_L g681 ( .A(n_604), .B(n_567), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_610), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_609), .B(n_616), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_615), .B(n_582), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_613), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_644), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_647), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_633), .A2(n_556), .B(n_588), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_681), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_664), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_660), .A2(n_628), .B1(n_638), .B2(n_601), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_687), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_660), .B(n_601), .C(n_630), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_661), .B(n_631), .Y(n_694) );
NOR4xp25_ASAP7_75t_SL g695 ( .A(n_688), .B(n_630), .C(n_611), .D(n_649), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_669), .B(n_619), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_688), .A2(n_633), .B1(n_648), .B2(n_635), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_671), .B(n_650), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_671), .B(n_631), .Y(n_699) );
AOI211xp5_ASAP7_75t_L g700 ( .A1(n_657), .A2(n_635), .B(n_588), .C(n_582), .Y(n_700) );
AOI32xp33_ASAP7_75t_L g701 ( .A1(n_666), .A2(n_629), .A3(n_646), .B1(n_642), .B2(n_581), .Y(n_701) );
OAI21x1_ASAP7_75t_SL g702 ( .A1(n_656), .A2(n_638), .B(n_637), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_652), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_681), .B(n_581), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_654), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_661), .B(n_637), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_655), .Y(n_707) );
OA21x2_ASAP7_75t_L g708 ( .A1(n_653), .A2(n_643), .B(n_627), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_681), .A2(n_648), .B(n_595), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_659), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_694), .B(n_663), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_692), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_703), .Y(n_713) );
OAI32xp33_ASAP7_75t_L g714 ( .A1(n_693), .A2(n_683), .A3(n_658), .B1(n_682), .B2(n_685), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_697), .A2(n_651), .B1(n_665), .B2(n_672), .C1(n_677), .C2(n_676), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_708), .Y(n_716) );
OAI22x1_ASAP7_75t_L g717 ( .A1(n_691), .A2(n_673), .B1(n_680), .B2(n_678), .Y(n_717) );
OAI322xp33_ASAP7_75t_L g718 ( .A1(n_691), .A2(n_667), .A3(n_668), .B1(n_670), .B2(n_674), .C1(n_686), .C2(n_645), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g719 ( .A1(n_700), .A2(n_589), .B(n_579), .C(n_596), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_708), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_699), .B(n_662), .Y(n_721) );
AOI322xp5_ASAP7_75t_L g722 ( .A1(n_696), .A2(n_679), .A3(n_675), .B1(n_684), .B2(n_574), .C1(n_627), .C2(n_623), .Y(n_722) );
OAI21xp33_ASAP7_75t_SL g723 ( .A1(n_701), .A2(n_476), .B(n_587), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_698), .B(n_591), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g725 ( .A1(n_702), .A2(n_467), .B(n_484), .Y(n_725) );
OAI21x1_ASAP7_75t_SL g726 ( .A1(n_709), .A2(n_573), .B(n_566), .Y(n_726) );
XNOR2x1_ASAP7_75t_L g727 ( .A(n_690), .B(n_573), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_695), .A2(n_566), .B(n_554), .Y(n_728) );
OAI221xp5_ASAP7_75t_SL g729 ( .A1(n_689), .A2(n_476), .B1(n_526), .B2(n_523), .C(n_514), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_704), .A2(n_523), .B(n_519), .Y(n_730) );
XOR2x1_ASAP7_75t_L g731 ( .A(n_727), .B(n_716), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_720), .Y(n_732) );
NAND4xp25_ASAP7_75t_SL g733 ( .A(n_715), .B(n_723), .C(n_722), .D(n_728), .Y(n_733) );
NOR2xp67_ASAP7_75t_L g734 ( .A(n_717), .B(n_712), .Y(n_734) );
AOI221x1_ASAP7_75t_L g735 ( .A1(n_719), .A2(n_713), .B1(n_725), .B2(n_726), .C(n_707), .Y(n_735) );
NOR2x1_ASAP7_75t_L g736 ( .A(n_733), .B(n_718), .Y(n_736) );
BUFx2_ASAP7_75t_L g737 ( .A(n_732), .Y(n_737) );
NAND4xp25_ASAP7_75t_L g738 ( .A(n_735), .B(n_715), .C(n_714), .D(n_729), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_737), .B(n_736), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_738), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_740), .Y(n_741) );
NAND3x1_ASAP7_75t_L g742 ( .A(n_739), .B(n_731), .C(n_734), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_741), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_743), .A2(n_742), .B(n_721), .Y(n_744) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_744), .B(n_704), .Y(n_745) );
AOI21xp33_ASAP7_75t_SL g746 ( .A1(n_745), .A2(n_711), .B(n_710), .Y(n_746) );
OR2x6_ASAP7_75t_L g747 ( .A(n_746), .B(n_705), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_747), .A2(n_724), .B1(n_706), .B2(n_730), .Y(n_748) );
endmodule