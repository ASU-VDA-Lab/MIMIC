module fake_jpeg_30610_n_456 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_456);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_456;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_49),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_59),
.Y(n_110)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_81),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_73),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_79),
.Y(n_141)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_85),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_90),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_89),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g88 ( 
.A(n_36),
.B(n_0),
.CON(n_88),
.SN(n_88)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_21),
.B(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_15),
.Y(n_136)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_91),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_33),
.B1(n_39),
.B2(n_21),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_106),
.B1(n_120),
.B2(n_121),
.Y(n_155)
);

OR2x2_ASAP7_75t_SL g192 ( 
.A(n_102),
.B(n_23),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_48),
.A2(n_33),
.B1(n_39),
.B2(n_21),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_103),
.A2(n_111),
.B1(n_124),
.B2(n_140),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_62),
.B1(n_58),
.B2(n_46),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_107),
.B(n_114),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_50),
.A2(n_88),
.B1(n_64),
.B2(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_49),
.A2(n_33),
.B1(n_46),
.B2(n_17),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_112),
.A2(n_144),
.B(n_10),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_74),
.B(n_44),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_17),
.B1(n_40),
.B2(n_38),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_40),
.B1(n_38),
.B2(n_28),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_137),
.B1(n_139),
.B2(n_142),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_77),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_87),
.B1(n_96),
.B2(n_45),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_151),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_84),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_86),
.A2(n_19),
.B1(n_18),
.B2(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_59),
.A2(n_19),
.B1(n_18),
.B2(n_45),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_19),
.C(n_45),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_153),
.Y(n_234)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_157),
.Y(n_244)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_160),
.B(n_162),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_45),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

OR2x4_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_90),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_164),
.A2(n_179),
.B(n_143),
.C(n_132),
.Y(n_223)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_169),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_45),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_178),
.Y(n_209)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_198),
.B1(n_100),
.B2(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_0),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_23),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_184),
.Y(n_220)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_186),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_193),
.Y(n_242)
);

BUFx8_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_104),
.B(n_1),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_202),
.C(n_125),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_23),
.Y(n_193)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_201),
.Y(n_232)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_199),
.B(n_150),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_194),
.B1(n_185),
.B2(n_157),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_200),
.Y(n_241)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

OR2x2_ASAP7_75t_SL g202 ( 
.A(n_113),
.B(n_2),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_127),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_206),
.B1(n_213),
.B2(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_161),
.B(n_148),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_175),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_155),
.A2(n_131),
.B1(n_108),
.B2(n_128),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_207),
.A2(n_214),
.B1(n_230),
.B2(n_231),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_105),
.B1(n_151),
.B2(n_147),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_131),
.B1(n_128),
.B2(n_108),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_147),
.B1(n_98),
.B2(n_138),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_147),
.B1(n_98),
.B2(n_138),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_216),
.A2(n_235),
.B1(n_132),
.B2(n_166),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_202),
.B(n_179),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_189),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_157),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_164),
.A2(n_98),
.B1(n_150),
.B2(n_122),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_152),
.B1(n_127),
.B2(n_113),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_156),
.A2(n_133),
.B1(n_125),
.B2(n_130),
.Y(n_235)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_247),
.B(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_168),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_251),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_190),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_253),
.A2(n_6),
.B(n_9),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_239),
.C(n_222),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_186),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_165),
.B1(n_195),
.B2(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_258),
.B(n_261),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_216),
.A2(n_125),
.B1(n_172),
.B2(n_177),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_191),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_229),
.A2(n_183),
.B1(n_181),
.B2(n_154),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_266),
.B1(n_240),
.B2(n_215),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_196),
.B1(n_176),
.B2(n_170),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_208),
.B(n_163),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_269),
.Y(n_295)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_3),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_280),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

BUFx4f_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_3),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_223),
.A2(n_145),
.B(n_132),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_277),
.B(n_231),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_244),
.A2(n_145),
.B(n_188),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_188),
.B(n_5),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_245),
.B(n_226),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_222),
.B(n_4),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_211),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_239),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_280)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_284),
.B(n_311),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_261),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_279),
.C(n_267),
.Y(n_325)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_204),
.B1(n_209),
.B2(n_234),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_308),
.B1(n_248),
.B2(n_271),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_232),
.C(n_241),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_301),
.C(n_309),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_221),
.C(n_234),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_269),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_307),
.B(n_314),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_248),
.A2(n_227),
.B1(n_236),
.B2(n_210),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_306),
.A2(n_266),
.B1(n_265),
.B2(n_250),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_236),
.B(n_221),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_256),
.A2(n_245),
.B1(n_226),
.B2(n_237),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_258),
.B(n_211),
.C(n_237),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_310),
.A2(n_312),
.B(n_307),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_251),
.B(n_238),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_238),
.B(n_218),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_278),
.B(n_274),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_275),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_303),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_291),
.B1(n_297),
.B2(n_306),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_317),
.A2(n_327),
.B1(n_281),
.B2(n_294),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_247),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_331),
.C(n_340),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_255),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_323),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_297),
.B1(n_313),
.B2(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_329),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_328),
.B(n_297),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_252),
.C(n_260),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_252),
.Y(n_332)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_264),
.Y(n_333)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_299),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_337),
.Y(n_368)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_336),
.A2(n_304),
.B(n_314),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_270),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_259),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_338),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_253),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_341),
.A2(n_291),
.B1(n_335),
.B2(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_281),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_342),
.B(n_343),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_289),
.B(n_277),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_338),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_355),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_288),
.C(n_310),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_354),
.C(n_358),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_365),
.B1(n_327),
.B2(n_294),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_356),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_340),
.C(n_339),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_313),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_318),
.B(n_308),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_273),
.C(n_283),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_302),
.C(n_257),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_326),
.C(n_338),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_352),
.B1(n_367),
.B2(n_355),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_321),
.A2(n_316),
.B1(n_343),
.B2(n_317),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_218),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_337),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_326),
.B(n_336),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_388),
.B1(n_359),
.B2(n_347),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_323),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_373),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_379),
.Y(n_393)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_350),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_383),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_320),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_381),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_384),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_357),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_366),
.B(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_316),
.B(n_334),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_389),
.B(n_361),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_292),
.B(n_262),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_390),
.A2(n_351),
.B1(n_358),
.B2(n_356),
.Y(n_398)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_396),
.A2(n_382),
.B1(n_376),
.B2(n_375),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_398),
.A2(n_402),
.B1(n_404),
.B2(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_401),
.B(n_406),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_390),
.A2(n_345),
.B1(n_354),
.B2(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_389),
.A2(n_345),
.B1(n_369),
.B2(n_360),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_349),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_408),
.B(n_412),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_399),
.B(n_374),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_416),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_374),
.C(n_371),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_415),
.C(n_393),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_371),
.C(n_376),
.Y(n_415)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_391),
.B(n_373),
.CI(n_370),
.CON(n_416),
.SN(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_399),
.B(n_384),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_417),
.B(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_268),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_396),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_400),
.A2(n_262),
.B(n_290),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_397),
.B(n_246),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_392),
.B1(n_395),
.B2(n_407),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_422),
.B1(n_410),
.B2(n_404),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_409),
.A2(n_395),
.B1(n_392),
.B2(n_394),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_423),
.B(n_429),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_412),
.B(n_391),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_426),
.C(n_430),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_418),
.C(n_415),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_431),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_405),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_434),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_409),
.B(n_414),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_401),
.B(n_419),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_436),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_426),
.A2(n_408),
.B(n_416),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_437),
.B(n_403),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_424),
.C(n_428),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_439),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_416),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_438),
.A2(n_403),
.B(n_263),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_441),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_445),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_224),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_444),
.A2(n_440),
.B1(n_446),
.B2(n_441),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_447),
.A2(n_448),
.B(n_212),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_433),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_452),
.C(n_450),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g452 ( 
.A(n_449),
.B(n_219),
.C(n_212),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_9),
.B(n_10),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_9),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_455),
.B(n_9),
.Y(n_456)
);


endmodule