module real_aes_7880_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g537 ( .A1(n_0), .A2(n_140), .B(n_538), .C(n_541), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_1), .B(n_482), .Y(n_542) );
INVx1_ASAP7_75t_L g425 ( .A(n_2), .Y(n_425) );
INVx1_ASAP7_75t_L g174 ( .A(n_3), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_4), .B(n_132), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_5), .A2(n_451), .B(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_6), .A2(n_117), .B(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_7), .A2(n_36), .B1(n_126), .B2(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_8), .B(n_117), .Y(n_143) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_10), .A2(n_141), .B(n_441), .C(n_443), .Y(n_440) );
AOI222xp33_ASAP7_75t_L g106 ( .A1(n_11), .A2(n_107), .B1(n_716), .B2(n_717), .C1(n_726), .C2(n_730), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_12), .B(n_37), .Y(n_426) );
INVx1_ASAP7_75t_L g167 ( .A(n_13), .Y(n_167) );
INVx1_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_15), .B(n_130), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_16), .B(n_132), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_17), .B(n_118), .Y(n_179) );
AO32x2_ASAP7_75t_L g201 ( .A1(n_18), .A2(n_117), .A3(n_147), .B1(n_158), .B2(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_19), .B(n_126), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_20), .B(n_118), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_21), .A2(n_56), .B1(n_126), .B2(n_204), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_22), .A2(n_84), .B1(n_126), .B2(n_130), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_23), .B(n_126), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_24), .A2(n_158), .B(n_441), .C(n_502), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_25), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_25), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_26), .A2(n_158), .B(n_441), .C(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_27), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_28), .B(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_29), .A2(n_451), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_30), .B(n_160), .Y(n_198) );
INVx2_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_32), .A2(n_453), .B(n_461), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_33), .B(n_126), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_34), .B(n_160), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_35), .B(n_212), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_38), .B(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_39), .B(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_40), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_41), .A2(n_80), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_41), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_42), .B(n_132), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_43), .B(n_451), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_44), .A2(n_81), .B1(n_420), .B2(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_44), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_45), .A2(n_453), .B(n_455), .C(n_461), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_46), .A2(n_721), .B1(n_724), .B2(n_725), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_46), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_47), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g539 ( .A(n_48), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_49), .A2(n_92), .B1(n_204), .B2(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g456 ( .A(n_50), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_51), .B(n_126), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_52), .B(n_126), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_53), .A2(n_747), .B1(n_748), .B2(n_750), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_53), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_54), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_55), .B(n_138), .Y(n_137) );
AOI22xp33_ASAP7_75t_SL g183 ( .A1(n_57), .A2(n_61), .B1(n_126), .B2(n_130), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_58), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_59), .B(n_126), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_60), .B(n_126), .Y(n_209) );
INVx1_ASAP7_75t_L g142 ( .A(n_62), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_63), .B(n_451), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_64), .B(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_65), .A2(n_138), .B(n_170), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_66), .B(n_126), .Y(n_175) );
INVx1_ASAP7_75t_L g121 ( .A(n_67), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_68), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_69), .B(n_132), .Y(n_492) );
AO32x2_ASAP7_75t_L g222 ( .A1(n_70), .A2(n_117), .A3(n_158), .B1(n_223), .B2(n_227), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_71), .B(n_133), .Y(n_444) );
INVx1_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
INVx1_ASAP7_75t_L g193 ( .A(n_73), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_74), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_75), .B(n_458), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_76), .A2(n_441), .B(n_461), .C(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_77), .B(n_130), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_78), .Y(n_477) );
INVx1_ASAP7_75t_L g738 ( .A(n_79), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_80), .Y(n_722) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_81), .A2(n_109), .B1(n_419), .B2(n_420), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_81), .Y(n_420) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_82), .A2(n_89), .B1(n_520), .B2(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_82), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_83), .B(n_457), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_85), .B(n_204), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_86), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_87), .B(n_130), .Y(n_197) );
INVx2_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_89), .A2(n_105), .B1(n_734), .B2(n_743), .C1(n_761), .C2(n_767), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_89), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_90), .B(n_157), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_91), .B(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g423 ( .A(n_93), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g715 ( .A(n_93), .Y(n_715) );
OR2x2_ASAP7_75t_L g742 ( .A(n_93), .B(n_733), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_94), .A2(n_103), .B1(n_130), .B2(n_131), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_95), .B(n_451), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_96), .Y(n_491) );
INVxp67_ASAP7_75t_L g480 ( .A(n_97), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_98), .B(n_130), .Y(n_151) );
INVx1_ASAP7_75t_L g437 ( .A(n_99), .Y(n_437) );
INVx1_ASAP7_75t_L g515 ( .A(n_100), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_101), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g463 ( .A(n_102), .B(n_160), .Y(n_463) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_421), .B1(n_427), .B2(n_712), .Y(n_107) );
INVx1_ASAP7_75t_L g727 ( .A(n_108), .Y(n_727) );
INVx2_ASAP7_75t_L g419 ( .A(n_109), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_109), .A2(n_419), .B1(n_754), .B2(n_755), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g109 ( .A(n_110), .B(n_343), .Y(n_109) );
AND2x2_ASAP7_75t_SL g110 ( .A(n_111), .B(n_301), .Y(n_110) );
NOR4xp25_ASAP7_75t_L g111 ( .A(n_112), .B(n_241), .C(n_277), .D(n_291), .Y(n_111) );
OAI221xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_185), .B1(n_217), .B2(n_228), .C(n_232), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_113), .B(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_161), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_144), .Y(n_115) );
AND2x2_ASAP7_75t_L g238 ( .A(n_116), .B(n_145), .Y(n_238) );
INVx3_ASAP7_75t_L g246 ( .A(n_116), .Y(n_246) );
AND2x2_ASAP7_75t_L g300 ( .A(n_116), .B(n_164), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_116), .B(n_163), .Y(n_336) );
AND2x2_ASAP7_75t_L g394 ( .A(n_116), .B(n_256), .Y(n_394) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_123), .B(n_143), .Y(n_116) );
INVx4_ASAP7_75t_L g184 ( .A(n_117), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_117), .A2(n_468), .B(n_469), .Y(n_467) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_117), .Y(n_474) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_119), .B(n_120), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_135), .B(n_141), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_132), .Y(n_124) );
INVx3_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_126), .Y(n_517) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g204 ( .A(n_127), .Y(n_204) );
BUFx3_ASAP7_75t_L g225 ( .A(n_127), .Y(n_225) );
AND2x6_ASAP7_75t_L g441 ( .A(n_127), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
INVx1_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
INVx2_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_132), .A2(n_150), .B(n_151), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_SL g191 ( .A1(n_132), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_132), .B(n_480), .Y(n_479) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_133), .A2(n_157), .B1(n_224), .B2(n_226), .Y(n_223) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
AND2x2_ASAP7_75t_L g439 ( .A(n_134), .B(n_139), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_134), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_140), .Y(n_135) );
INVx2_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_140), .A2(n_154), .B(n_174), .C(n_175), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g181 ( .A1(n_140), .A2(n_157), .B1(n_182), .B2(n_183), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_140), .A2(n_157), .B1(n_203), .B2(n_205), .Y(n_202) );
BUFx3_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_141), .A2(n_166), .B(n_173), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_141), .A2(n_191), .B(n_195), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_141), .A2(n_208), .B(n_213), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_141), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g451 ( .A(n_141), .B(n_439), .Y(n_451) );
INVx4_ASAP7_75t_SL g462 ( .A(n_141), .Y(n_462) );
AND2x2_ASAP7_75t_L g229 ( .A(n_144), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g243 ( .A(n_144), .B(n_164), .Y(n_243) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_145), .B(n_164), .Y(n_258) );
AND2x2_ASAP7_75t_L g270 ( .A(n_145), .B(n_246), .Y(n_270) );
OR2x2_ASAP7_75t_L g272 ( .A(n_145), .B(n_230), .Y(n_272) );
AND2x2_ASAP7_75t_L g307 ( .A(n_145), .B(n_230), .Y(n_307) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_145), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_145), .Y(n_360) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_159), .Y(n_145) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_146), .A2(n_165), .B(n_176), .Y(n_164) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_147), .B(n_447), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_158), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_155), .C(n_156), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_154), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_156), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g540 ( .A(n_157), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_158), .B(n_181), .C(n_184), .Y(n_180) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_190), .B(n_198), .Y(n_189) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_160), .A2(n_207), .B(n_216), .Y(n_206) );
INVx2_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_160), .A2(n_450), .B(n_452), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_160), .A2(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g508 ( .A(n_160), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g277 ( .A1(n_161), .A2(n_278), .B1(n_282), .B2(n_286), .C(n_287), .Y(n_277) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g237 ( .A(n_162), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_177), .Y(n_162) );
INVx2_ASAP7_75t_L g236 ( .A(n_163), .Y(n_236) );
AND2x2_ASAP7_75t_L g289 ( .A(n_163), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g308 ( .A(n_163), .B(n_246), .Y(n_308) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g371 ( .A(n_164), .B(n_246), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_169), .C(n_170), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_168), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_168), .A2(n_471), .B(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_170), .A2(n_515), .B(n_516), .C(n_517), .Y(n_514) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_171), .A2(n_196), .B(n_197), .Y(n_195) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g458 ( .A(n_172), .Y(n_458) );
AND2x2_ASAP7_75t_L g293 ( .A(n_177), .B(n_238), .Y(n_293) );
OAI322xp33_ASAP7_75t_L g361 ( .A1(n_177), .A2(n_317), .A3(n_362), .B1(n_364), .B2(n_367), .C1(n_369), .C2(n_373), .Y(n_361) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2x1_ASAP7_75t_L g244 ( .A(n_178), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
AND2x2_ASAP7_75t_L g366 ( .A(n_178), .B(n_246), .Y(n_366) );
AND2x2_ASAP7_75t_L g398 ( .A(n_178), .B(n_270), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_178), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
AO21x1_ASAP7_75t_L g230 ( .A1(n_181), .A2(n_184), .B(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_184), .A2(n_436), .B(n_446), .Y(n_435) );
INVx3_ASAP7_75t_L g482 ( .A(n_184), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_184), .B(n_494), .Y(n_493) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_184), .A2(n_512), .B(n_519), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_184), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_199), .Y(n_186) );
INVx1_ASAP7_75t_L g414 ( .A(n_187), .Y(n_414) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g219 ( .A(n_188), .B(n_206), .Y(n_219) );
INVx2_ASAP7_75t_L g254 ( .A(n_188), .Y(n_254) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_189), .Y(n_284) );
OR2x2_ASAP7_75t_L g408 ( .A(n_189), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g233 ( .A(n_199), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g273 ( .A(n_199), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g325 ( .A(n_199), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_206), .Y(n_199) );
AND2x2_ASAP7_75t_L g220 ( .A(n_200), .B(n_221), .Y(n_220) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_200), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g334 ( .A(n_200), .B(n_222), .Y(n_334) );
OR2x2_ASAP7_75t_L g342 ( .A(n_200), .B(n_276), .Y(n_342) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
AND2x2_ASAP7_75t_L g261 ( .A(n_201), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g285 ( .A(n_201), .B(n_206), .Y(n_285) );
AND2x2_ASAP7_75t_L g349 ( .A(n_201), .B(n_222), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_206), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_206), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g262 ( .A(n_206), .Y(n_262) );
INVx1_ASAP7_75t_L g267 ( .A(n_206), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_206), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_206), .Y(n_357) );
INVx1_ASAP7_75t_L g409 ( .A(n_206), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
AND2x2_ASAP7_75t_L g386 ( .A(n_218), .B(n_295), .Y(n_386) );
INVx2_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g313 ( .A(n_220), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g412 ( .A(n_220), .B(n_347), .Y(n_412) );
INVx1_ASAP7_75t_L g234 ( .A(n_221), .Y(n_234) );
AND2x2_ASAP7_75t_L g260 ( .A(n_221), .B(n_254), .Y(n_260) );
BUFx2_ASAP7_75t_L g319 ( .A(n_221), .Y(n_319) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_222), .Y(n_240) );
INVx1_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_225), .Y(n_460) );
INVx2_ASAP7_75t_L g541 ( .A(n_225), .Y(n_541) );
INVx1_ASAP7_75t_L g505 ( .A(n_227), .Y(n_505) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_228), .B(n_235), .Y(n_388) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI32xp33_ASAP7_75t_L g232 ( .A1(n_229), .A2(n_233), .A3(n_235), .B1(n_237), .B2(n_239), .Y(n_232) );
AND2x2_ASAP7_75t_L g372 ( .A(n_229), .B(n_245), .Y(n_372) );
AND2x2_ASAP7_75t_L g410 ( .A(n_229), .B(n_308), .Y(n_410) );
INVx1_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_234), .B(n_296), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_235), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_235), .B(n_238), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_235), .B(n_307), .Y(n_389) );
OR2x2_ASAP7_75t_L g403 ( .A(n_235), .B(n_272), .Y(n_403) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g330 ( .A(n_236), .B(n_238), .Y(n_330) );
OR2x2_ASAP7_75t_L g339 ( .A(n_236), .B(n_326), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_238), .B(n_289), .Y(n_311) );
INVx2_ASAP7_75t_L g326 ( .A(n_240), .Y(n_326) );
OR2x2_ASAP7_75t_L g341 ( .A(n_240), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g356 ( .A(n_240), .B(n_357), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g413 ( .A1(n_240), .A2(n_333), .B(n_414), .C(n_415), .Y(n_413) );
OAI321xp33_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_247), .A3(n_252), .B1(n_255), .B2(n_259), .C(n_263), .Y(n_241) );
INVx1_ASAP7_75t_L g354 ( .A(n_242), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g365 ( .A(n_243), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g317 ( .A(n_245), .Y(n_317) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_246), .B(n_360), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_247), .A2(n_385), .B1(n_387), .B2(n_389), .C(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND2x2_ASAP7_75t_L g322 ( .A(n_249), .B(n_296), .Y(n_322) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_250), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g295 ( .A(n_251), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_252), .A2(n_293), .B(n_338), .C(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g304 ( .A(n_254), .B(n_261), .Y(n_304) );
BUFx2_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
INVx1_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OR2x2_ASAP7_75t_L g335 ( .A(n_257), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g418 ( .A(n_257), .Y(n_418) );
INVx1_ASAP7_75t_L g411 ( .A(n_258), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_260), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g368 ( .A(n_260), .B(n_285), .Y(n_368) );
INVx1_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_268), .B1(n_271), .B2(n_273), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_265), .B(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_L g333 ( .A(n_266), .B(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_267), .B(n_276), .Y(n_296) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g288 ( .A(n_270), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g298 ( .A(n_272), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_275), .A2(n_393), .B1(n_395), .B2(n_396), .C(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g281 ( .A(n_276), .Y(n_281) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_276), .Y(n_347) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_279), .B(n_398), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_280), .A2(n_285), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_283), .B(n_293), .Y(n_390) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g359 ( .A(n_284), .Y(n_359) );
AND2x2_ASAP7_75t_L g318 ( .A(n_285), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g407 ( .A(n_285), .Y(n_407) );
INVx1_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g378 ( .A(n_289), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B1(n_297), .B2(n_298), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_295), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g363 ( .A(n_296), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_296), .B(n_334), .Y(n_400) );
OR2x2_ASAP7_75t_L g373 ( .A(n_297), .B(n_326), .Y(n_373) );
INVx1_ASAP7_75t_L g312 ( .A(n_298), .Y(n_312) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_300), .B(n_351), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_320), .C(n_331), .Y(n_301) );
OAI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_309), .C(n_315), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_304), .A2(n_375), .B1(n_379), .B2(n_382), .C(n_384), .Y(n_374) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_307), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g370 ( .A(n_307), .B(n_371), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_356), .B(n_358), .C(n_360), .Y(n_355) );
INVx2_ASAP7_75t_L g402 ( .A(n_308), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_312), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g381 ( .A(n_314), .B(n_334), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
OAI21xp5_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_323), .B(n_324), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_327), .B(n_330), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_325), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_330), .B(n_417), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_337), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g358 ( .A(n_334), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND4x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_374), .C(n_391), .D(n_413), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_361), .Y(n_344) );
OAI211xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_350), .B(n_353), .C(n_355), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_349), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_360), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g395 ( .A(n_370), .Y(n_395) );
INVx2_ASAP7_75t_SL g383 ( .A(n_371), .Y(n_383) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g396 ( .A(n_381), .Y(n_396) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_399), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_401), .B1(n_403), .B2(n_404), .C(n_405), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_410), .B1(n_411), .B2(n_412), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g728 ( .A(n_422), .Y(n_728) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g714 ( .A(n_424), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g733 ( .A(n_424), .Y(n_733) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_428), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
OR3x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_610), .C(n_675), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g429 ( .A(n_430), .B(n_551), .C(n_577), .D(n_600), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_483), .B1(n_521), .B2(n_528), .C(n_543), .Y(n_430) );
CKINVDCx14_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_432), .A2(n_544), .B1(n_568), .B2(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_464), .Y(n_432) );
INVx1_ASAP7_75t_SL g604 ( .A(n_433), .Y(n_604) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_448), .Y(n_433) );
OR2x2_ASAP7_75t_L g526 ( .A(n_434), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g546 ( .A(n_434), .B(n_465), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_434), .B(n_473), .Y(n_559) );
AND2x2_ASAP7_75t_L g576 ( .A(n_434), .B(n_448), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_434), .B(n_524), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_434), .B(n_575), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_434), .B(n_464), .Y(n_697) );
AOI211xp5_ASAP7_75t_SL g708 ( .A1(n_434), .A2(n_614), .B(n_709), .C(n_710), .Y(n_708) );
INVx5_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_435), .B(n_465), .Y(n_580) );
AND2x2_ASAP7_75t_L g583 ( .A(n_435), .B(n_466), .Y(n_583) );
OR2x2_ASAP7_75t_L g628 ( .A(n_435), .B(n_465), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_435), .B(n_473), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_440), .Y(n_436) );
INVx5_ASAP7_75t_L g454 ( .A(n_441), .Y(n_454) );
INVx5_ASAP7_75t_SL g527 ( .A(n_448), .Y(n_527) );
AND2x2_ASAP7_75t_L g545 ( .A(n_448), .B(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_448), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g631 ( .A(n_448), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g663 ( .A(n_448), .B(n_473), .Y(n_663) );
OR2x2_ASAP7_75t_L g669 ( .A(n_448), .B(n_559), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_448), .B(n_619), .Y(n_678) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_463), .Y(n_448) );
BUFx2_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_454), .A2(n_462), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_454), .A2(n_462), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_459), .C(n_460), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_457), .A2(n_460), .B(n_491), .C(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
AND2x2_ASAP7_75t_L g560 ( .A(n_465), .B(n_527), .Y(n_560) );
INVx1_ASAP7_75t_SL g573 ( .A(n_465), .Y(n_573) );
OR2x2_ASAP7_75t_L g608 ( .A(n_465), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g614 ( .A(n_465), .B(n_473), .Y(n_614) );
AND2x2_ASAP7_75t_L g672 ( .A(n_465), .B(n_524), .Y(n_672) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_466), .B(n_527), .Y(n_599) );
INVx3_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
OR2x2_ASAP7_75t_L g565 ( .A(n_473), .B(n_527), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_473), .B(n_573), .Y(n_575) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_473), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_473), .B(n_546), .Y(n_632) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_482), .A2(n_534), .B(n_542), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_483), .A2(n_649), .B1(n_651), .B2(n_653), .C(n_656), .Y(n_648) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .Y(n_484) );
AND2x2_ASAP7_75t_L g622 ( .A(n_485), .B(n_603), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_485), .B(n_681), .Y(n_685) );
OR2x2_ASAP7_75t_L g706 ( .A(n_485), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_485), .B(n_711), .Y(n_710) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx5_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
AND2x2_ASAP7_75t_L g630 ( .A(n_486), .B(n_497), .Y(n_630) );
AND2x2_ASAP7_75t_L g691 ( .A(n_486), .B(n_570), .Y(n_691) );
AND2x2_ASAP7_75t_L g704 ( .A(n_486), .B(n_524), .Y(n_704) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_509), .Y(n_495) );
AND2x4_ASAP7_75t_L g531 ( .A(n_496), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g549 ( .A(n_496), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g556 ( .A(n_496), .Y(n_556) );
AND2x2_ASAP7_75t_L g625 ( .A(n_496), .B(n_603), .Y(n_625) );
AND2x2_ASAP7_75t_L g635 ( .A(n_496), .B(n_553), .Y(n_635) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_496), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_496), .B(n_533), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_496), .B(n_587), .Y(n_659) );
AND2x2_ASAP7_75t_L g696 ( .A(n_496), .B(n_691), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_496), .B(n_570), .Y(n_707) );
OR2x2_ASAP7_75t_L g709 ( .A(n_496), .B(n_645), .Y(n_709) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g595 ( .A(n_497), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g605 ( .A(n_497), .B(n_550), .Y(n_605) );
AND2x2_ASAP7_75t_L g617 ( .A(n_497), .B(n_533), .Y(n_617) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_497), .Y(n_647) );
AND2x4_ASAP7_75t_L g681 ( .A(n_497), .B(n_532), .Y(n_681) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_506), .Y(n_497) );
AOI21xp5_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_501), .B(n_505), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
BUFx2_ASAP7_75t_L g530 ( .A(n_509), .Y(n_530) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
AND2x2_ASAP7_75t_L g603 ( .A(n_510), .B(n_533), .Y(n_603) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g550 ( .A(n_511), .B(n_533), .Y(n_550) );
BUFx2_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_523), .B(n_604), .Y(n_683) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_524), .B(n_546), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_524), .B(n_527), .Y(n_585) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_576), .Y(n_640) );
AOI221xp5_ASAP7_75t_SL g577 ( .A1(n_525), .A2(n_578), .B1(n_586), .B2(n_588), .C(n_592), .Y(n_577) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g613 ( .A(n_526), .B(n_614), .Y(n_613) );
OAI321xp33_ASAP7_75t_L g620 ( .A1(n_526), .A2(n_579), .A3(n_621), .B1(n_623), .B2(n_624), .C(n_626), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_527), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_530), .B(n_681), .Y(n_699) );
AND2x2_ASAP7_75t_L g586 ( .A(n_531), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_532), .Y(n_562) );
AND2x2_ASAP7_75t_L g569 ( .A(n_532), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_532), .B(n_644), .Y(n_674) );
INVx1_ASAP7_75t_L g711 ( .A(n_532), .Y(n_711) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B(n_548), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_545), .A2(n_655), .B(n_704), .C(n_705), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_546), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_546), .B(n_584), .Y(n_650) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g593 ( .A(n_550), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_550), .B(n_553), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_550), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_550), .B(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B1(n_566), .B2(n_571), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g567 ( .A(n_553), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_553), .B(n_596), .Y(n_638) );
OR2x2_ASAP7_75t_L g645 ( .A(n_553), .B(n_570), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_553), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g695 ( .A(n_553), .B(n_681), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .B1(n_561), .B2(n_563), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g601 ( .A(n_556), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_559), .A2(n_574), .B1(n_642), .B2(n_646), .Y(n_641) );
INVx1_ASAP7_75t_L g689 ( .A(n_560), .Y(n_689) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_564), .A2(n_601), .B1(n_604), .B2(n_605), .C(n_606), .Y(n_600) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g579 ( .A(n_565), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_569), .B(n_635), .Y(n_667) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_570), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_570), .Y(n_591) );
NAND2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g609 ( .A(n_576), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_576), .B(n_619), .Y(n_618) );
NAND2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g662 ( .A(n_583), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_612), .B1(n_615), .B2(n_618), .C(n_620), .Y(n_611) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_590), .B(n_647), .Y(n_646) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B(n_597), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_597), .Y(n_694) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
OR2x2_ASAP7_75t_L g636 ( .A(n_599), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g657 ( .A(n_602), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_602), .B(n_662), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_605), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_629), .C(n_648), .D(n_661), .Y(n_610) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g619 ( .A(n_614), .Y(n_619) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g652 ( .A(n_623), .B(n_628), .Y(n_652) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_633), .C(n_641), .Y(n_629) );
AOI211xp5_ASAP7_75t_L g700 ( .A1(n_631), .A2(n_673), .B(n_701), .C(n_708), .Y(n_700) );
INVx1_ASAP7_75t_SL g660 ( .A(n_632), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g664 ( .A(n_638), .Y(n_664) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_644), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_644), .B(n_655), .Y(n_688) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g665 ( .A(n_655), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B(n_660), .Y(n_656) );
INVxp33_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .A3(n_665), .B1(n_666), .B2(n_668), .C1(n_670), .C2(n_673), .Y(n_661) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g675 ( .A(n_676), .B(n_693), .C(n_700), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g692 ( .A(n_681), .Y(n_692) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_696), .B2(n_697), .C(n_698), .Y(n_693) );
NAND2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g729 ( .A(n_713), .Y(n_729) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_715), .B(n_733), .Y(n_732) );
CKINVDCx16_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_740), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g736 ( .A(n_737), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_SL g766 ( .A(n_737), .Y(n_766) );
INVx1_ASAP7_75t_L g765 ( .A(n_739), .Y(n_765) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_739), .A2(n_766), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g744 ( .A(n_742), .Y(n_744) );
INVx2_ASAP7_75t_L g760 ( .A(n_742), .Y(n_760) );
BUFx2_ASAP7_75t_L g769 ( .A(n_742), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B(n_757), .Y(n_743) );
XOR2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_751), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
CKINVDCx6p67_ASAP7_75t_R g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
endmodule