module fake_ariane_1554_n_2585 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2585);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2585;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_762;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_59),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_315),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_508),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_127),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_267),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_42),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_167),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_85),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_224),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_195),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_105),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_479),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_244),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_387),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_0),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_349),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_403),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_517),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_295),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_323),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_275),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_382),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_346),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_549),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_446),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_18),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_174),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_129),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_242),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_231),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_270),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_390),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_311),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_520),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_141),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_73),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_410),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_548),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_365),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_426),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_184),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_377),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_254),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_126),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_188),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_454),
.Y(n_606)
);

BUFx2_ASAP7_75t_SL g607 ( 
.A(n_28),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_17),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_498),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_363),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_70),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_285),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_44),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_408),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_237),
.Y(n_615)
);

BUFx8_ASAP7_75t_SL g616 ( 
.A(n_64),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_209),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_170),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_424),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_545),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_450),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_147),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_21),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_546),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_193),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_511),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_31),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_286),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_263),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_481),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_1),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_85),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_521),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_489),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_382),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_529),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_140),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_551),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_206),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_200),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_482),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_426),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_547),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_552),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_190),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_354),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_79),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_543),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g649 ( 
.A(n_480),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_31),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_358),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_205),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_209),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_257),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_392),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_0),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_101),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_540),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_335),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_484),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_194),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_199),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_470),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_465),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_305),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_315),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_516),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_371),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_74),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_9),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_378),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_15),
.Y(n_672)
);

CKINVDCx14_ASAP7_75t_R g673 ( 
.A(n_344),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_329),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_499),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_228),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_42),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_312),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_101),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_200),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_550),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_19),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_34),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_86),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_168),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_412),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_77),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_158),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_278),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_424),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_241),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_338),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_36),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_257),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_453),
.Y(n_697)
);

CKINVDCx16_ASAP7_75t_R g698 ( 
.A(n_110),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_386),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_23),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_176),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_265),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_429),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_374),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_285),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_294),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_555),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_449),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_17),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_297),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_442),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_471),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_468),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_171),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_544),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_162),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_33),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_254),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_201),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_391),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_169),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_466),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_501),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_259),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_252),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_20),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_338),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_48),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_416),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_57),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_414),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_538),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_161),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_477),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_96),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_473),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_542),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_303),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_298),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_513),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_553),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_283),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_415),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_414),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_539),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_367),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_397),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_334),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_62),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_369),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_220),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_231),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_288),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_38),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_485),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_195),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_161),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_541),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_393),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_557),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_160),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_240),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_183),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_206),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_281),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_95),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_413),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_154),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_533),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_383),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_378),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_554),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_556),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_183),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_132),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_323),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_398),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_439),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_300),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_247),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_144),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_333),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_404),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_92),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_63),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_345),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_199),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_534),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_577),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_635),
.Y(n_791)
);

INVxp67_ASAP7_75t_SL g792 ( 
.A(n_635),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_673),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_651),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_651),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_719),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_616),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_645),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_738),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_719),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_756),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_739),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_739),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_561),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_643),
.Y(n_805)
);

INVxp33_ASAP7_75t_SL g806 ( 
.A(n_707),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_563),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_651),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_577),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_760),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_633),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_651),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_677),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_677),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_677),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_677),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_583),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_565),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_564),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_694),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_566),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_607),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_649),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_570),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_571),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_585),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_585),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_573),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_594),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_598),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_602),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_603),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_610),
.Y(n_835)
);

CKINVDCx14_ASAP7_75t_R g836 ( 
.A(n_579),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_611),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_612),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_618),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_619),
.Y(n_840)
);

INVxp33_ASAP7_75t_SL g841 ( 
.A(n_565),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_628),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_664),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_629),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_631),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_637),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_675),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_732),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_640),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_642),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_694),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_694),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_694),
.Y(n_853)
);

INVxp33_ASAP7_75t_L g854 ( 
.A(n_650),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_694),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_576),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_659),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_722),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_610),
.Y(n_859)
);

INVxp33_ASAP7_75t_SL g860 ( 
.A(n_567),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_698),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_732),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_661),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_666),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_668),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_678),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_680),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_699),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_683),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_681),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_686),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_699),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_695),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_700),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_652),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_702),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_705),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_575),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_687),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_718),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_730),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_576),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_733),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_575),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_652),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_716),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_744),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_808),
.Y(n_889)
);

BUFx12f_ASAP7_75t_L g890 ( 
.A(n_797),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_848),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_855),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_805),
.B(n_697),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_805),
.B(n_715),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_848),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_879),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_848),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_879),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_811),
.B(n_717),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_797),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_848),
.Y(n_902)
);

BUFx12f_ASAP7_75t_L g903 ( 
.A(n_793),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_811),
.B(n_717),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_792),
.B(n_745),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_861),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_861),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_806),
.B(n_772),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_794),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_836),
.B(n_755),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_862),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_793),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_875),
.B(n_576),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_806),
.B(n_638),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_862),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_794),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_862),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_862),
.Y(n_918)
);

BUFx8_ASAP7_75t_L g919 ( 
.A(n_810),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_795),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_804),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_795),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_810),
.B(n_708),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_807),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_818),
.B(n_579),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_862),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_817),
.Y(n_927)
);

BUFx8_ASAP7_75t_SL g928 ( 
.A(n_789),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_817),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_885),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_822),
.Y(n_932)
);

BUFx8_ASAP7_75t_SL g933 ( 
.A(n_789),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_852),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_854),
.B(n_653),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_852),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_821),
.Y(n_937)
);

AND2x6_ASAP7_75t_L g938 ( 
.A(n_870),
.B(n_600),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_853),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_791),
.B(n_653),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_885),
.Y(n_941)
);

BUFx8_ASAP7_75t_SL g942 ( 
.A(n_809),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_853),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_790),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_814),
.B(n_601),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_796),
.B(n_653),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_814),
.B(n_767),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_819),
.B(n_737),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_790),
.Y(n_949)
);

NOR2x1_ASAP7_75t_L g950 ( 
.A(n_843),
.B(n_778),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_800),
.B(n_662),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_870),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_812),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_909),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_927),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_909),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_927),
.Y(n_958)
);

BUFx8_ASAP7_75t_L g959 ( 
.A(n_890),
.Y(n_959)
);

INVxp33_ASAP7_75t_SL g960 ( 
.A(n_925),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_916),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_924),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_927),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_889),
.B(n_847),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_916),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_920),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_937),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_892),
.B(n_847),
.Y(n_968)
);

AND2x6_ASAP7_75t_L g969 ( 
.A(n_940),
.B(n_601),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_952),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_952),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_895),
.B(n_818),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_920),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_906),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_927),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_952),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_945),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_922),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_880),
.B(n_813),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_908),
.B(n_825),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_930),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_944),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_900),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_912),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_927),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_893),
.A2(n_841),
.B1(n_860),
.B2(n_819),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_900),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_938),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_896),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_938),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_940),
.B(n_758),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_948),
.B(n_914),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_929),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_946),
.B(n_951),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_900),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_929),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_944),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_904),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_903),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_904),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_904),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_944),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_923),
.B(n_825),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_896),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_947),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_944),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_929),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_947),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_905),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_929),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_944),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_912),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_949),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_946),
.B(n_858),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_896),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_951),
.B(n_823),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_949),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_949),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_949),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_949),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_910),
.B(n_858),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_953),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_953),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_913),
.B(n_824),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_953),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_950),
.B(n_826),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_935),
.B(n_880),
.Y(n_1029)
);

BUFx8_ASAP7_75t_L g1030 ( 
.A(n_890),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_953),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_929),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_935),
.B(n_913),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_928),
.Y(n_1034)
);

XNOR2xp5_ASAP7_75t_L g1035 ( 
.A(n_897),
.B(n_809),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_931),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_953),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_932),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_932),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_903),
.Y(n_1040)
);

OA21x2_ASAP7_75t_L g1041 ( 
.A1(n_938),
.A2(n_813),
.B(n_812),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_932),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_979),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_1033),
.B(n_897),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_956),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1033),
.A2(n_860),
.B1(n_841),
.B2(n_938),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_979),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_995),
.B(n_899),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_995),
.B(n_899),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_979),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_995),
.B(n_993),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_962),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_957),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_957),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_961),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_993),
.B(n_941),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_1029),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_972),
.B(n_856),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1011),
.B(n_569),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_985),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_961),
.Y(n_1061)
);

CKINVDCx6p67_ASAP7_75t_R g1062 ( 
.A(n_1000),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_977),
.B(n_1029),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_965),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_974),
.B(n_799),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_989),
.B(n_569),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_989),
.B(n_991),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_965),
.Y(n_1068)
);

NOR2x1p5_ASAP7_75t_L g1069 ( 
.A(n_1000),
.B(n_901),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_967),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_966),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_1018),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_985),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_966),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_980),
.A2(n_693),
.B1(n_584),
.B2(n_581),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_970),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_971),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_976),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_984),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_969),
.A2(n_938),
.B1(n_801),
.B2(n_798),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_987),
.B(n_1023),
.C(n_1004),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_989),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_988),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_996),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_955),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_991),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_969),
.B(n_883),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_1018),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_969),
.B(n_938),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_991),
.B(n_582),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_973),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_973),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_954),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1026),
.B(n_919),
.C(n_907),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_990),
.Y(n_1095)
);

INVxp67_ASAP7_75t_R g1096 ( 
.A(n_1036),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_954),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_990),
.B(n_582),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_990),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_1040),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_969),
.B(n_919),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_999),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1001),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1005),
.B(n_758),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_969),
.B(n_919),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1005),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1002),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_969),
.A2(n_716),
.B1(n_763),
.B2(n_646),
.Y(n_1108)
);

CKINVDCx6p67_ASAP7_75t_R g1109 ( 
.A(n_1034),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_981),
.Y(n_1111)
);

INVxp33_ASAP7_75t_SL g1112 ( 
.A(n_1035),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_981),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_955),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_982),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1014),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_992),
.B(n_767),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1009),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_992),
.B(n_567),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_992),
.B(n_558),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_1010),
.B(n_901),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_960),
.B(n_907),
.Y(n_1122)
);

NOR2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1016),
.B(n_1018),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_982),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_559),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1005),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_992),
.B(n_562),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1017),
.B(n_732),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_978),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1017),
.B(n_732),
.Y(n_1130)
);

INVx6_ASAP7_75t_L g1131 ( 
.A(n_959),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_964),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_998),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_983),
.A2(n_816),
.B(n_815),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_998),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_1017),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_968),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1014),
.B(n_802),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_SL g1139 ( 
.A(n_992),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1003),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_983),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_974),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1028),
.B(n_803),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_SL g1145 ( 
.A(n_1028),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1003),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_959),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1015),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_959),
.Y(n_1149)
);

INVxp33_ASAP7_75t_L g1150 ( 
.A(n_1035),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1041),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1028),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_955),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1013),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1007),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1007),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_960),
.B(n_593),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1020),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1019),
.B(n_907),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1041),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1020),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1021),
.A2(n_763),
.B1(n_615),
.B2(n_704),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1041),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1025),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1025),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1022),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_955),
.B(n_732),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_958),
.B(n_560),
.Y(n_1169)
);

NOR2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1030),
.B(n_568),
.Y(n_1170)
);

NAND2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1027),
.B(n_568),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1034),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_958),
.B(n_592),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1027),
.B(n_828),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1024),
.B(n_595),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1031),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1037),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1042),
.B(n_599),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1038),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1085),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1079),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1083),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1085),
.Y(n_1184)
);

CKINVDCx16_ASAP7_75t_R g1185 ( 
.A(n_1100),
.Y(n_1185)
);

NOR2xp67_ASAP7_75t_L g1186 ( 
.A(n_1122),
.B(n_827),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1084),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_1073),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1102),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1053),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1143),
.B(n_828),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1081),
.B(n_1039),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1053),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1054),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1116),
.B(n_829),
.Y(n_1195)
);

XNOR2xp5_ASAP7_75t_L g1196 ( 
.A(n_1112),
.B(n_829),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1058),
.B(n_835),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1103),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1051),
.B(n_958),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_1082),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1107),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1110),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_L g1203 ( 
.A(n_1094),
.B(n_830),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1051),
.A2(n_963),
.B(n_958),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1118),
.Y(n_1205)
);

XNOR2xp5_ASAP7_75t_L g1206 ( 
.A(n_1112),
.B(n_835),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_1060),
.B(n_831),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1045),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1044),
.B(n_958),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1052),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1138),
.B(n_859),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1056),
.B(n_859),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1072),
.B(n_994),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1056),
.B(n_868),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1085),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1070),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1093),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1093),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1097),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1097),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1096),
.B(n_1174),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1054),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1147),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1062),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1111),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1065),
.B(n_868),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

INVxp33_ASAP7_75t_L g1228 ( 
.A(n_1150),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1158),
.B(n_872),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1062),
.Y(n_1230)
);

XOR2xp5_ASAP7_75t_L g1231 ( 
.A(n_1150),
.B(n_872),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1055),
.Y(n_1232)
);

CKINVDCx16_ASAP7_75t_R g1233 ( 
.A(n_1147),
.Y(n_1233)
);

INVx4_ASAP7_75t_SL g1234 ( 
.A(n_1139),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1113),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_887),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1098),
.A2(n_1012),
.B(n_1008),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1115),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1115),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1109),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1088),
.B(n_887),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1124),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1088),
.B(n_832),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1124),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1129),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1085),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1109),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1057),
.B(n_833),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1082),
.Y(n_1249)
);

BUFx8_ASAP7_75t_L g1250 ( 
.A(n_1172),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1131),
.B(n_1030),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1057),
.B(n_834),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1129),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1076),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1153),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1055),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1131),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1132),
.B(n_963),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_R g1259 ( 
.A(n_1121),
.B(n_1030),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1048),
.B(n_963),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1077),
.Y(n_1261)
);

XOR2xp5_ASAP7_75t_L g1262 ( 
.A(n_1149),
.B(n_1101),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1078),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1142),
.Y(n_1264)
);

BUFx8_ASAP7_75t_L g1265 ( 
.A(n_1149),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1148),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1152),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1155),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1061),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1167),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1131),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1095),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1176),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1061),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1048),
.B(n_963),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1177),
.Y(n_1276)
);

INVxp67_ASAP7_75t_SL g1277 ( 
.A(n_1082),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1180),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1144),
.B(n_837),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1064),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1049),
.B(n_975),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1064),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1068),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1163),
.B(n_838),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1068),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1069),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1071),
.Y(n_1287)
);

INVxp33_ASAP7_75t_SL g1288 ( 
.A(n_1160),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1063),
.B(n_975),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1071),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1123),
.B(n_839),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1086),
.B(n_975),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1108),
.B(n_840),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1074),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_R g1295 ( 
.A(n_1121),
.B(n_1105),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1121),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1121),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1074),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1091),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1049),
.B(n_842),
.Y(n_1300)
);

XOR2xp5_ASAP7_75t_L g1301 ( 
.A(n_1075),
.B(n_928),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1091),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1178),
.B(n_844),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1092),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1092),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1137),
.B(n_975),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1170),
.B(n_845),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1171),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1099),
.B(n_975),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1086),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1133),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_1059),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1133),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1098),
.A2(n_997),
.B(n_994),
.Y(n_1314)
);

INVxp33_ASAP7_75t_L g1315 ( 
.A(n_1059),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1135),
.Y(n_1316)
);

XOR2x2_ASAP7_75t_L g1317 ( 
.A(n_1080),
.B(n_933),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1135),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1087),
.B(n_942),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1140),
.Y(n_1320)
);

XOR2xp5_ASAP7_75t_L g1321 ( 
.A(n_1046),
.B(n_942),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1140),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1175),
.B(n_846),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1146),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1099),
.B(n_986),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1117),
.B(n_849),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1146),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1156),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1156),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1157),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1114),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1145),
.B(n_725),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1157),
.Y(n_1333)
);

XOR2xp5_ASAP7_75t_L g1334 ( 
.A(n_1120),
.B(n_572),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1159),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1159),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1162),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1171),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1125),
.B(n_850),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1145),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1162),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1166),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1166),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1179),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1127),
.B(n_857),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1179),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1165),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1145),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1165),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1043),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1086),
.B(n_863),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1043),
.B(n_864),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1099),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1047),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1047),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1114),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1050),
.Y(n_1357)
);

AND2x6_ASAP7_75t_L g1358 ( 
.A(n_1139),
.B(n_986),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1106),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1169),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1114),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1106),
.B(n_986),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1050),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1106),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1134),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1104),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1169),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1151),
.A2(n_866),
.B(n_865),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1104),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1151),
.Y(n_1370)
);

XNOR2xp5_ASAP7_75t_L g1371 ( 
.A(n_1173),
.B(n_867),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1151),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1173),
.B(n_869),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1066),
.A2(n_994),
.B(n_986),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1114),
.B(n_986),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1161),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1095),
.B(n_994),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1161),
.Y(n_1378)
);

BUFx5_ASAP7_75t_L g1379 ( 
.A(n_1067),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1161),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1217),
.B(n_1095),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1288),
.B(n_1136),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1186),
.B(n_1188),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1265),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1197),
.B(n_1136),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1212),
.A2(n_1139),
.B1(n_1119),
.B2(n_692),
.Y(n_1386)
);

BUFx4_ASAP7_75t_L g1387 ( 
.A(n_1185),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1279),
.B(n_1126),
.Y(n_1388)
);

BUFx8_ASAP7_75t_L g1389 ( 
.A(n_1195),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1208),
.Y(n_1390)
);

AND2x6_ASAP7_75t_SL g1391 ( 
.A(n_1226),
.B(n_871),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1211),
.B(n_662),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1218),
.B(n_1136),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1210),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1303),
.B(n_1141),
.Y(n_1395)
);

BUFx5_ASAP7_75t_L g1396 ( 
.A(n_1358),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1188),
.B(n_1141),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1248),
.B(n_1141),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1265),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1190),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1252),
.B(n_1141),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1251),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1251),
.B(n_1089),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1229),
.A2(n_1119),
.B1(n_692),
.B2(n_768),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1243),
.B(n_1255),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1191),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1216),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1251),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1182),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1183),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1193),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1293),
.B(n_1154),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1192),
.A2(n_1130),
.B(n_1128),
.C(n_1090),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1321),
.A2(n_774),
.B1(n_766),
.B2(n_574),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1236),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1214),
.B(n_1312),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1300),
.B(n_1066),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1192),
.B(n_1130),
.C(n_1128),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1315),
.B(n_1090),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1187),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1189),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1310),
.A2(n_751),
.B1(n_753),
.B2(n_749),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1198),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1310),
.A2(n_757),
.B1(n_761),
.B2(n_754),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1194),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1284),
.B(n_1164),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1228),
.B(n_1164),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_SL g1429 ( 
.A(n_1257),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1201),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1241),
.B(n_662),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1196),
.B(n_1164),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1291),
.B(n_572),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1224),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_R g1435 ( 
.A(n_1230),
.B(n_574),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1351),
.B(n_578),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1358),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1206),
.B(n_578),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1202),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1332),
.B(n_692),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1250),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1351),
.B(n_580),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1223),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1205),
.B(n_580),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1254),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1326),
.B(n_586),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1339),
.B(n_586),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1345),
.B(n_587),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1219),
.B(n_1067),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1222),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1261),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1207),
.B(n_587),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1308),
.A2(n_1338),
.B1(n_1319),
.B2(n_1360),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1199),
.A2(n_1168),
.B(n_779),
.C(n_783),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1334),
.B(n_588),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1340),
.B(n_1168),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1263),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1307),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1317),
.A2(n_768),
.B1(n_734),
.B2(n_589),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1199),
.A2(n_771),
.B(n_874),
.C(n_873),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1268),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1270),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1371),
.B(n_997),
.Y(n_1463)
);

INVx5_ASAP7_75t_L g1464 ( 
.A(n_1358),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1352),
.B(n_588),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1271),
.Y(n_1466)
);

NOR3xp33_ASAP7_75t_L g1467 ( 
.A(n_1260),
.B(n_780),
.C(n_590),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1260),
.B(n_997),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1264),
.B(n_589),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1232),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1234),
.B(n_886),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1231),
.B(n_590),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1266),
.B(n_1267),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1273),
.B(n_591),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1276),
.B(n_591),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1367),
.A2(n_768),
.B1(n_734),
.B2(n_776),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1256),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1181),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1245),
.A2(n_734),
.B1(n_777),
.B2(n_776),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1204),
.A2(n_877),
.B(n_876),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1278),
.B(n_777),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1259),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1253),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1275),
.A2(n_597),
.B1(n_605),
.B2(n_604),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1233),
.B(n_780),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1368),
.B(n_782),
.C(n_781),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1220),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1340),
.B(n_878),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1250),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1181),
.B(n_997),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1281),
.A2(n_613),
.B1(n_614),
.B2(n_608),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1235),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1238),
.B(n_782),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1269),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1296),
.B(n_784),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1239),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1336),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1242),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1244),
.B(n_784),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1353),
.B(n_785),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1200),
.A2(n_786),
.B1(n_787),
.B2(n_785),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1297),
.B(n_786),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1348),
.B(n_787),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1358),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1281),
.B(n_1008),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1353),
.B(n_1359),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1282),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1283),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1323),
.B(n_881),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1274),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1350),
.B(n_882),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1348),
.B(n_884),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1272),
.B(n_1008),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1290),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1294),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1209),
.B(n_617),
.Y(n_1517)
);

INVx8_ASAP7_75t_L g1518 ( 
.A(n_1240),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1209),
.B(n_1008),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1280),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1301),
.A2(n_623),
.B1(n_625),
.B2(n_622),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1354),
.B(n_1355),
.Y(n_1522)
);

AO22x1_ASAP7_75t_L g1523 ( 
.A1(n_1286),
.A2(n_632),
.B1(n_639),
.B2(n_627),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1285),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1181),
.B(n_1012),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1373),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1287),
.Y(n_1527)
);

BUFx4_ASAP7_75t_L g1528 ( 
.A(n_1247),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1357),
.B(n_888),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_L g1530 ( 
.A(n_1379),
.B(n_1012),
.Y(n_1530)
);

O2A1O1Ixp5_ASAP7_75t_L g1531 ( 
.A1(n_1374),
.A2(n_851),
.B(n_820),
.C(n_886),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1298),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1295),
.A2(n_654),
.B1(n_655),
.B2(n_647),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1184),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1311),
.A2(n_657),
.B1(n_665),
.B2(n_656),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1234),
.B(n_1012),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1299),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1320),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1333),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1364),
.B(n_669),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_L g1541 ( 
.A(n_1379),
.B(n_1012),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1302),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1363),
.B(n_670),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1184),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1184),
.B(n_1032),
.Y(n_1545)
);

NOR3xp33_ASAP7_75t_L g1546 ( 
.A(n_1289),
.B(n_672),
.C(n_671),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_L g1547 ( 
.A(n_1379),
.B(n_1215),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1262),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1304),
.Y(n_1549)
);

INVx8_ASAP7_75t_L g1550 ( 
.A(n_1215),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1341),
.A2(n_676),
.B1(n_679),
.B2(n_674),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_L g1552 ( 
.A(n_1379),
.B(n_1032),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1234),
.B(n_1032),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1368),
.B(n_684),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1258),
.B(n_685),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1305),
.A2(n_689),
.B1(n_690),
.B2(n_688),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1313),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1316),
.A2(n_696),
.B1(n_701),
.B2(n_691),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_SL g1559 ( 
.A(n_1246),
.B(n_703),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1347),
.B(n_706),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1318),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1322),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1324),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1349),
.B(n_709),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1246),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1246),
.Y(n_1566)
);

NOR2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1258),
.B(n_714),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1327),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1306),
.B(n_720),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1328),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1329),
.B(n_1330),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1335),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1200),
.B(n_721),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1337),
.Y(n_1574)
);

BUFx5_ASAP7_75t_L g1575 ( 
.A(n_1370),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1366),
.B(n_724),
.Y(n_1576)
);

AND2x6_ASAP7_75t_SL g1577 ( 
.A(n_1362),
.B(n_820),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1414),
.A2(n_1419),
.B(n_1531),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1458),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1385),
.B(n_1203),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1390),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1530),
.A2(n_1277),
.B(n_1249),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1394),
.Y(n_1583)
);

AO21x1_ASAP7_75t_L g1584 ( 
.A1(n_1517),
.A2(n_1314),
.B(n_1237),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1541),
.A2(n_1552),
.B(n_1377),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1381),
.A2(n_1377),
.B(n_1325),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1438),
.A2(n_1342),
.B1(n_1344),
.B2(n_1343),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1408),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1381),
.A2(n_1325),
.B(n_1309),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1389),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1382),
.B(n_1346),
.Y(n_1591)
);

AO21x1_ASAP7_75t_L g1592 ( 
.A1(n_1519),
.A2(n_1204),
.B(n_1369),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1393),
.A2(n_1309),
.B(n_1362),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1417),
.B(n_1405),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1526),
.B(n_1331),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1466),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1393),
.A2(n_1376),
.B(n_1372),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1547),
.A2(n_1380),
.B(n_1378),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1392),
.B(n_1432),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1464),
.B(n_1437),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1407),
.B(n_1440),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_L g1604 ( 
.A(n_1399),
.B(n_1213),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1410),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1388),
.A2(n_1292),
.B1(n_1361),
.B2(n_1356),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1395),
.B(n_1356),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1455),
.A2(n_727),
.B1(n_728),
.B2(n_726),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1416),
.B(n_729),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1514),
.A2(n_1375),
.B(n_1365),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1570),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1453),
.B(n_1032),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1486),
.A2(n_735),
.B1(n_742),
.B2(n_731),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1411),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1548),
.B(n_1032),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1525),
.A2(n_851),
.B(n_606),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1472),
.A2(n_746),
.B1(n_747),
.B2(n_743),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1498),
.B(n_748),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1420),
.B(n_932),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1545),
.A2(n_609),
.B(n_596),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1502),
.B(n_1447),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1498),
.B(n_750),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1441),
.B(n_932),
.Y(n_1623)
);

NOR2x1_ASAP7_75t_L g1624 ( 
.A(n_1544),
.B(n_934),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1449),
.A2(n_621),
.B(n_620),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1534),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1503),
.A2(n_759),
.B1(n_762),
.B2(n_752),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1459),
.A2(n_765),
.B1(n_770),
.B2(n_764),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1449),
.A2(n_626),
.B(n_624),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1431),
.B(n_775),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1473),
.A2(n_636),
.B(n_630),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1572),
.Y(n_1632)
);

NOR2x2_ASAP7_75t_L g1633 ( 
.A(n_1387),
.B(n_1),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_SL g1634 ( 
.A1(n_1397),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1428),
.B(n_934),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1434),
.B(n_432),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1465),
.B(n_934),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1386),
.B(n_934),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1486),
.A2(n_644),
.B1(n_648),
.B2(n_641),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1468),
.A2(n_660),
.B(n_658),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1480),
.A2(n_911),
.B(n_894),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1464),
.B(n_934),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1506),
.A2(n_667),
.B(n_663),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1398),
.A2(n_711),
.B(n_682),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1421),
.Y(n_1645)
);

BUFx4f_ASAP7_75t_L g1646 ( 
.A(n_1518),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1448),
.B(n_936),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1401),
.A2(n_713),
.B(n_712),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1443),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1404),
.A2(n_736),
.B(n_740),
.C(n_723),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1485),
.B(n_741),
.Y(n_1651)
);

O2A1O1Ixp33_ASAP7_75t_SL g1652 ( 
.A1(n_1573),
.A2(n_1507),
.B(n_1554),
.C(n_1418),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1550),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1427),
.A2(n_773),
.B(n_769),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1422),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1400),
.Y(n_1656)
);

AO21x1_ASAP7_75t_L g1657 ( 
.A1(n_1480),
.A2(n_939),
.B(n_936),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1437),
.Y(n_1658)
);

INVx11_ASAP7_75t_L g1659 ( 
.A(n_1389),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1412),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1489),
.A2(n_788),
.B(n_936),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1391),
.B(n_2),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1489),
.A2(n_1464),
.B(n_1522),
.Y(n_1663)
);

AO21x1_ASAP7_75t_L g1664 ( 
.A1(n_1555),
.A2(n_1569),
.B(n_1413),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1491),
.A2(n_939),
.B(n_936),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1518),
.Y(n_1666)
);

INVx5_ASAP7_75t_L g1667 ( 
.A(n_1505),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1426),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1467),
.B(n_939),
.C(n_898),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1533),
.B(n_939),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1513),
.B(n_1415),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1423),
.B(n_3),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1488),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1550),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1423),
.B(n_4),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1383),
.B(n_5),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1523),
.B(n_5),
.C(n_6),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1425),
.B(n_6),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1415),
.B(n_7),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1435),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_SL g1681 ( 
.A1(n_1501),
.A2(n_1406),
.B(n_1469),
.C(n_1454),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1478),
.B(n_943),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1576),
.A2(n_1510),
.B(n_1425),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1518),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1424),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1550),
.Y(n_1686)
);

XOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1482),
.B(n_433),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1452),
.A2(n_1500),
.B(n_1494),
.C(n_1436),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1504),
.B(n_7),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1460),
.A2(n_943),
.B(n_902),
.C(n_918),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1543),
.A2(n_911),
.B(n_894),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1540),
.A2(n_943),
.B(n_902),
.C(n_918),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1446),
.A2(n_911),
.B(n_894),
.Y(n_1693)
);

INVx11_ASAP7_75t_L g1694 ( 
.A(n_1528),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1430),
.B(n_8),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1439),
.B(n_8),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1396),
.B(n_943),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1445),
.B(n_9),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1451),
.B(n_10),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1433),
.B(n_10),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1457),
.B(n_11),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1450),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1461),
.A2(n_902),
.B(n_891),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1442),
.B(n_11),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1478),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1462),
.A2(n_902),
.B(n_891),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1463),
.B(n_12),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1512),
.B(n_1529),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1470),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1478),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1484),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1711)
);

AND2x2_ASAP7_75t_SL g1712 ( 
.A(n_1490),
.B(n_13),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1560),
.A2(n_911),
.B(n_894),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1566),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1505),
.A2(n_902),
.B(n_891),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1521),
.B(n_14),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_L g1717 ( 
.A(n_1546),
.B(n_1474),
.C(n_1444),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1566),
.Y(n_1718)
);

O2A1O1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1564),
.A2(n_18),
.B(n_15),
.C(n_16),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1566),
.B(n_918),
.Y(n_1720)
);

AND2x6_ASAP7_75t_L g1721 ( 
.A(n_1536),
.B(n_918),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1536),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1471),
.B(n_926),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1544),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1553),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1487),
.A2(n_926),
.B(n_915),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1483),
.B(n_1475),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1481),
.B(n_1493),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1497),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1499),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1567),
.A2(n_926),
.B(n_915),
.C(n_917),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1471),
.B(n_894),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1402),
.B(n_16),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1508),
.A2(n_917),
.B(n_915),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1565),
.A2(n_917),
.B(n_915),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1509),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1409),
.B(n_434),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1384),
.Y(n_1738)
);

NAND2x1p5_ASAP7_75t_L g1739 ( 
.A(n_1553),
.B(n_917),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1515),
.A2(n_19),
.B(n_20),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1477),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1496),
.B(n_21),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1492),
.A2(n_24),
.B(n_25),
.C(n_23),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1479),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1429),
.B(n_22),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1456),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1403),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1495),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1516),
.B(n_26),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1537),
.B(n_26),
.C(n_27),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1476),
.B(n_27),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1511),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1403),
.A2(n_436),
.B(n_435),
.Y(n_1753)
);

AO21x1_ASAP7_75t_L g1754 ( 
.A1(n_1542),
.A2(n_28),
.B(n_29),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1575),
.B(n_29),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1549),
.A2(n_30),
.B(n_32),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1403),
.B(n_437),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1556),
.B(n_30),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1557),
.A2(n_440),
.B(n_438),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1561),
.B(n_32),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1562),
.B(n_33),
.Y(n_1761)
);

O2A1O1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1689),
.A2(n_1558),
.B(n_1551),
.C(n_1535),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1685),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1600),
.B(n_1563),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1651),
.B(n_1429),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1657),
.A2(n_1574),
.B(n_1524),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1580),
.B(n_1575),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_L g1768 ( 
.A(n_1626),
.B(n_1520),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1594),
.B(n_1577),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1602),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1673),
.B(n_1597),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1621),
.A2(n_1456),
.B1(n_1559),
.B2(n_1532),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1680),
.B(n_1596),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1582),
.A2(n_1585),
.B(n_1641),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1641),
.A2(n_1396),
.B(n_1575),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1730),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1727),
.B(n_1527),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1593),
.A2(n_1396),
.B(n_1575),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1581),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1649),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1672),
.A2(n_1396),
.B1(n_1539),
.B2(n_1538),
.Y(n_1782)
);

AO22x1_ASAP7_75t_L g1783 ( 
.A1(n_1662),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1757),
.B(n_35),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1728),
.B(n_37),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1586),
.A2(n_37),
.B(n_38),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1675),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1611),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1589),
.A2(n_39),
.B(n_40),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1757),
.B(n_41),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1579),
.Y(n_1791)
);

OAI21xp33_ASAP7_75t_L g1792 ( 
.A1(n_1700),
.A2(n_43),
.B(n_44),
.Y(n_1792)
);

BUFx8_ASAP7_75t_L g1793 ( 
.A(n_1590),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1708),
.B(n_43),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1671),
.B(n_45),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1603),
.B(n_45),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1598),
.A2(n_46),
.B(n_47),
.Y(n_1797)
);

NAND2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1626),
.B(n_1653),
.Y(n_1798)
);

AOI22x1_ASAP7_75t_L g1799 ( 
.A1(n_1740),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1599),
.A2(n_49),
.B(n_50),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1663),
.A2(n_49),
.B(n_50),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1678),
.A2(n_1742),
.B1(n_1704),
.B2(n_1683),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1722),
.B(n_441),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1583),
.B(n_51),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1684),
.B(n_51),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1588),
.B(n_52),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1713),
.A2(n_52),
.B(n_53),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1743),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1605),
.Y(n_1809)
);

INVx5_ASAP7_75t_L g1810 ( 
.A(n_1721),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1666),
.B(n_1712),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1679),
.B(n_54),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1738),
.B(n_55),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1653),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1614),
.Y(n_1815)
);

NOR3xp33_ASAP7_75t_L g1816 ( 
.A(n_1711),
.B(n_56),
.C(n_57),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1632),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1659),
.B(n_56),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1653),
.B(n_443),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1694),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1646),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1618),
.B(n_58),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1622),
.B(n_60),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1645),
.B(n_61),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1688),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1646),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1676),
.B(n_65),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1674),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1674),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1655),
.B(n_66),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1664),
.B(n_67),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1729),
.B(n_67),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1713),
.A2(n_68),
.B(n_69),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1674),
.Y(n_1834)
);

A2O1A1Ixp33_ASAP7_75t_SL g1835 ( 
.A1(n_1719),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1736),
.B(n_71),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1595),
.B(n_71),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1697),
.A2(n_72),
.B(n_73),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1656),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1660),
.Y(n_1840)
);

O2A1O1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1677),
.A2(n_75),
.B(n_72),
.C(n_74),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_SL g1842 ( 
.A(n_1636),
.B(n_444),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1668),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1697),
.A2(n_1578),
.B(n_1691),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1717),
.B(n_75),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1578),
.A2(n_1691),
.B(n_1652),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1705),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1686),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1734),
.A2(n_76),
.B(n_77),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1734),
.A2(n_1693),
.B(n_1692),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1627),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1702),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1667),
.B(n_78),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1693),
.A2(n_80),
.B(n_81),
.Y(n_1854)
);

OAI21xp33_ASAP7_75t_L g1855 ( 
.A1(n_1740),
.A2(n_80),
.B(n_81),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1587),
.B(n_82),
.Y(n_1856)
);

INVx5_ASAP7_75t_L g1857 ( 
.A(n_1721),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1630),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1667),
.B(n_82),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1758),
.B(n_83),
.Y(n_1860)
);

AO21x1_ASAP7_75t_L g1861 ( 
.A1(n_1756),
.A2(n_83),
.B(n_84),
.Y(n_1861)
);

AOI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1584),
.A2(n_447),
.B(n_445),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1744),
.A2(n_87),
.B(n_84),
.C(n_86),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1686),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1681),
.A2(n_87),
.B(n_88),
.Y(n_1865)
);

NOR3xp33_ASAP7_75t_L g1866 ( 
.A(n_1756),
.B(n_88),
.C(n_89),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1628),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1751),
.B(n_90),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1716),
.B(n_91),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1610),
.A2(n_92),
.B(n_93),
.Y(n_1870)
);

NAND2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1686),
.B(n_448),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1725),
.B(n_1722),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1608),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1709),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1715),
.A2(n_94),
.B(n_96),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1667),
.B(n_97),
.Y(n_1876)
);

O2A1O1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1650),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1741),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1761),
.B(n_98),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_SL g1880 ( 
.A1(n_1750),
.A2(n_102),
.B(n_99),
.C(n_100),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1726),
.A2(n_100),
.B(n_102),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1718),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1745),
.B(n_103),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1695),
.B(n_103),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_SL g1885 ( 
.A(n_1722),
.B(n_451),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1617),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1748),
.Y(n_1887)
);

OR2x6_ASAP7_75t_L g1888 ( 
.A(n_1747),
.B(n_452),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1703),
.A2(n_104),
.B(n_106),
.Y(n_1889)
);

AO21x1_ASAP7_75t_L g1890 ( 
.A1(n_1612),
.A2(n_107),
.B(n_108),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1606),
.B(n_107),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1706),
.A2(n_108),
.B(n_109),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1615),
.B(n_109),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1696),
.B(n_1698),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1699),
.A2(n_1701),
.B1(n_1707),
.B2(n_1749),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1733),
.B(n_110),
.Y(n_1896)
);

AOI22x1_ASAP7_75t_L g1897 ( 
.A1(n_1631),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1760),
.A2(n_1613),
.B1(n_1669),
.B2(n_1755),
.Y(n_1898)
);

AND2x6_ASAP7_75t_L g1899 ( 
.A(n_1747),
.B(n_455),
.Y(n_1899)
);

CKINVDCx11_ASAP7_75t_R g1900 ( 
.A(n_1714),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1661),
.A2(n_111),
.B(n_112),
.Y(n_1901)
);

OAI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1669),
.A2(n_113),
.B(n_114),
.Y(n_1902)
);

BUFx4f_ASAP7_75t_L g1903 ( 
.A(n_1601),
.Y(n_1903)
);

A2O1A1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1625),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1724),
.B(n_115),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1721),
.Y(n_1906)
);

AO32x1_ASAP7_75t_L g1907 ( 
.A1(n_1752),
.A2(n_118),
.A3(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1747),
.B(n_456),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1687),
.B(n_117),
.Y(n_1909)
);

O2A1O1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1634),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_1910)
);

BUFx4_ASAP7_75t_SL g1911 ( 
.A(n_1633),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1710),
.Y(n_1912)
);

NOR2x1p5_ASAP7_75t_SL g1913 ( 
.A(n_1592),
.B(n_457),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1658),
.B(n_120),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1658),
.B(n_121),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1629),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1638),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1746),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1654),
.A2(n_124),
.B(n_125),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1725),
.B(n_125),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1609),
.B(n_126),
.Y(n_1921)
);

AO22x1_ASAP7_75t_L g1922 ( 
.A1(n_1604),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1780),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_SL g1924 ( 
.A(n_1827),
.B(n_1754),
.C(n_1639),
.Y(n_1924)
);

AO31x2_ASAP7_75t_L g1925 ( 
.A1(n_1846),
.A2(n_1731),
.A3(n_1690),
.B(n_1635),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1777),
.B(n_1714),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1802),
.A2(n_1753),
.B(n_1759),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1844),
.A2(n_1619),
.B(n_1720),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1809),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1771),
.B(n_1607),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1815),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1763),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1774),
.A2(n_1670),
.B(n_1682),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1770),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1862),
.A2(n_1665),
.B(n_1624),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1850),
.A2(n_1776),
.B(n_1779),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1810),
.A2(n_1647),
.B(n_1637),
.Y(n_1937)
);

A2O1A1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1762),
.A2(n_1737),
.B(n_1648),
.C(n_1644),
.Y(n_1938)
);

AND3x2_ASAP7_75t_L g1939 ( 
.A(n_1765),
.B(n_1623),
.C(n_1601),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1788),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1791),
.B(n_1723),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1817),
.Y(n_1942)
);

AOI211x1_ASAP7_75t_L g1943 ( 
.A1(n_1783),
.A2(n_1643),
.B(n_1640),
.C(n_1620),
.Y(n_1943)
);

NAND2x1p5_ASAP7_75t_L g1944 ( 
.A(n_1810),
.B(n_1857),
.Y(n_1944)
);

OAI21x1_ASAP7_75t_SL g1945 ( 
.A1(n_1861),
.A2(n_1616),
.B(n_1735),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_SL g1946 ( 
.A1(n_1855),
.A2(n_1732),
.B(n_1739),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1781),
.B(n_1739),
.Y(n_1947)
);

AO21x2_ASAP7_75t_L g1948 ( 
.A1(n_1831),
.A2(n_1721),
.B(n_1642),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1810),
.B(n_458),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1818),
.B(n_128),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1766),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1866),
.A2(n_130),
.B(n_131),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1858),
.B(n_130),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1764),
.B(n_131),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1874),
.Y(n_1955)
);

OAI21x1_ASAP7_75t_L g1956 ( 
.A1(n_1865),
.A2(n_460),
.B(n_459),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1857),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1766),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1839),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1857),
.A2(n_132),
.B(n_133),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1870),
.A2(n_462),
.B(n_461),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1840),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1801),
.A2(n_464),
.B(n_463),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1795),
.B(n_133),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1789),
.A2(n_469),
.B(n_467),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1882),
.B(n_134),
.Y(n_1966)
);

OAI21x1_ASAP7_75t_L g1967 ( 
.A1(n_1767),
.A2(n_474),
.B(n_472),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1769),
.B(n_134),
.Y(n_1968)
);

OAI21x1_ASAP7_75t_L g1969 ( 
.A1(n_1786),
.A2(n_476),
.B(n_475),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1847),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1807),
.A2(n_135),
.B(n_136),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1833),
.A2(n_135),
.B(n_136),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1812),
.B(n_137),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1894),
.B(n_137),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_L g1975 ( 
.A(n_1792),
.B(n_1816),
.C(n_1825),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1778),
.B(n_138),
.Y(n_1976)
);

A2O1A1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1921),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1814),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1918),
.Y(n_1979)
);

NAND3xp33_ASAP7_75t_L g1980 ( 
.A(n_1845),
.B(n_139),
.C(n_141),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1773),
.B(n_142),
.Y(n_1981)
);

AND2x6_ASAP7_75t_L g1982 ( 
.A(n_1782),
.B(n_478),
.Y(n_1982)
);

A2O1A1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1822),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_1983)
);

AOI211x1_ASAP7_75t_L g1984 ( 
.A1(n_1868),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1800),
.A2(n_487),
.B(n_483),
.Y(n_1985)
);

NOR2xp67_ASAP7_75t_L g1986 ( 
.A(n_1837),
.B(n_145),
.Y(n_1986)
);

INVx2_ASAP7_75t_SL g1987 ( 
.A(n_1793),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1912),
.B(n_1869),
.Y(n_1988)
);

AND2x6_ASAP7_75t_L g1989 ( 
.A(n_1872),
.B(n_1920),
.Y(n_1989)
);

OAI21x1_ASAP7_75t_SL g1990 ( 
.A1(n_1799),
.A2(n_146),
.B(n_147),
.Y(n_1990)
);

OA21x2_ASAP7_75t_L g1991 ( 
.A1(n_1902),
.A2(n_148),
.B(n_149),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1775),
.A2(n_148),
.B(n_149),
.Y(n_1992)
);

OAI21x1_ASAP7_75t_SL g1993 ( 
.A1(n_1890),
.A2(n_150),
.B(n_151),
.Y(n_1993)
);

OAI21x1_ASAP7_75t_L g1994 ( 
.A1(n_1854),
.A2(n_490),
.B(n_488),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1849),
.A2(n_150),
.B(n_151),
.Y(n_1995)
);

NAND2x1_ASAP7_75t_L g1996 ( 
.A(n_1899),
.B(n_152),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1823),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1900),
.Y(n_1998)
);

NOR2x1_ASAP7_75t_L g1999 ( 
.A(n_1895),
.B(n_153),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1814),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1797),
.A2(n_492),
.B(n_491),
.Y(n_2001)
);

A2O1A1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1877),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_L g2003 ( 
.A1(n_1889),
.A2(n_494),
.B(n_493),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1785),
.B(n_1879),
.Y(n_2004)
);

OAI21xp33_ASAP7_75t_L g2005 ( 
.A1(n_1787),
.A2(n_155),
.B(n_156),
.Y(n_2005)
);

OAI22x1_ASAP7_75t_L g2006 ( 
.A1(n_1811),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1892),
.A2(n_1881),
.B(n_1875),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1898),
.A2(n_159),
.B(n_162),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1873),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1794),
.B(n_163),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_1905),
.B(n_164),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1843),
.Y(n_2012)
);

AO22x1_ASAP7_75t_L g2013 ( 
.A1(n_1899),
.A2(n_1793),
.B1(n_1896),
.B2(n_1911),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1909),
.B(n_165),
.Y(n_2014)
);

INVx4_ASAP7_75t_SL g2015 ( 
.A(n_1899),
.Y(n_2015)
);

AO32x2_ASAP7_75t_L g2016 ( 
.A1(n_1772),
.A2(n_168),
.A3(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1872),
.B(n_495),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1838),
.A2(n_166),
.B(n_170),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1901),
.A2(n_497),
.B(n_496),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1804),
.B(n_171),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1897),
.A2(n_502),
.B(n_500),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1820),
.B(n_172),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1887),
.Y(n_2023)
);

OAI21x1_ASAP7_75t_L g2024 ( 
.A1(n_1819),
.A2(n_504),
.B(n_503),
.Y(n_2024)
);

AOI21x1_ASAP7_75t_SL g2025 ( 
.A1(n_1884),
.A2(n_172),
.B(n_173),
.Y(n_2025)
);

OAI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1808),
.A2(n_173),
.B(n_174),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1796),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1806),
.B(n_175),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_2015),
.B(n_1903),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1926),
.Y(n_2030)
);

INVxp67_ASAP7_75t_L g2031 ( 
.A(n_1932),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1998),
.B(n_1820),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1923),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2027),
.B(n_1824),
.Y(n_2034)
);

NAND2xp33_ASAP7_75t_L g2035 ( 
.A(n_2005),
.B(n_1999),
.Y(n_2035)
);

O2A1O1Ixp5_ASAP7_75t_SL g2036 ( 
.A1(n_1979),
.A2(n_1951),
.B(n_1958),
.C(n_1927),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1936),
.A2(n_1790),
.B(n_1784),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1933),
.A2(n_1891),
.B(n_1903),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1923),
.B(n_1929),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1946),
.A2(n_1910),
.B(n_1907),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1988),
.B(n_1883),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1931),
.B(n_1830),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1959),
.Y(n_2043)
);

BUFx12f_ASAP7_75t_L g2044 ( 
.A(n_1998),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1941),
.B(n_1930),
.Y(n_2045)
);

BUFx12f_ASAP7_75t_L g2046 ( 
.A(n_1998),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1970),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1947),
.B(n_1832),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_2015),
.B(n_1768),
.Y(n_2049)
);

NOR2xp33_ASAP7_75t_L g2050 ( 
.A(n_1950),
.B(n_1813),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1954),
.B(n_1920),
.Y(n_2051)
);

INVx5_ASAP7_75t_L g2052 ( 
.A(n_1982),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1981),
.B(n_1987),
.Y(n_2053)
);

OAI21xp33_ASAP7_75t_L g2054 ( 
.A1(n_1952),
.A2(n_1826),
.B(n_1821),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1944),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_2004),
.B(n_1836),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1964),
.B(n_1973),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1978),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1976),
.B(n_1860),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1928),
.A2(n_1937),
.B(n_1975),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1959),
.B(n_1962),
.Y(n_2061)
);

BUFx10_ASAP7_75t_L g2062 ( 
.A(n_2022),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1984),
.A2(n_1856),
.B1(n_1917),
.B2(n_1886),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1966),
.Y(n_2064)
);

AOI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_1924),
.A2(n_1907),
.B(n_1835),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1962),
.Y(n_2066)
);

INVx5_ASAP7_75t_SL g2067 ( 
.A(n_2017),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1978),
.B(n_1805),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2012),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1938),
.A2(n_1907),
.B(n_1863),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1974),
.B(n_1922),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2012),
.B(n_1852),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_1957),
.B(n_1848),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1951),
.B(n_1913),
.Y(n_2074)
);

BUFx10_ASAP7_75t_L g2075 ( 
.A(n_1953),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1968),
.B(n_1878),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1934),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1939),
.Y(n_2078)
);

CKINVDCx20_ASAP7_75t_R g2079 ( 
.A(n_2014),
.Y(n_2079)
);

NAND2x1p5_ASAP7_75t_L g2080 ( 
.A(n_1996),
.B(n_1814),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_2000),
.Y(n_2081)
);

INVx5_ASAP7_75t_L g2082 ( 
.A(n_1982),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_2000),
.Y(n_2083)
);

BUFx2_ASAP7_75t_R g2084 ( 
.A(n_1948),
.Y(n_2084)
);

CKINVDCx8_ASAP7_75t_R g2085 ( 
.A(n_1989),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1989),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1983),
.A2(n_1851),
.B1(n_1841),
.B2(n_1867),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2011),
.B(n_1829),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1986),
.B(n_1829),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_1925),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1977),
.A2(n_1880),
.B(n_1916),
.C(n_1904),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_2013),
.Y(n_2092)
);

NOR2x1_ASAP7_75t_SL g2093 ( 
.A(n_1949),
.B(n_1906),
.Y(n_2093)
);

INVxp33_ASAP7_75t_L g2094 ( 
.A(n_2078),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2052),
.A2(n_1982),
.B1(n_1989),
.B2(n_1991),
.Y(n_2095)
);

INVx8_ASAP7_75t_L g2096 ( 
.A(n_2044),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2043),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2061),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2061),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2033),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_2052),
.Y(n_2101)
);

BUFx4f_ASAP7_75t_SL g2102 ( 
.A(n_2046),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2054),
.A2(n_1995),
.B1(n_2026),
.B2(n_1991),
.Y(n_2103)
);

INVx4_ASAP7_75t_L g2104 ( 
.A(n_2052),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2066),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_2047),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2054),
.A2(n_1980),
.B1(n_1982),
.B2(n_2018),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2035),
.A2(n_2008),
.B1(n_1971),
.B2(n_1972),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2039),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_SL g2110 ( 
.A1(n_2082),
.A2(n_1989),
.B1(n_1993),
.B2(n_2016),
.Y(n_2110)
);

CKINVDCx6p67_ASAP7_75t_R g2111 ( 
.A(n_2062),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_2076),
.Y(n_2112)
);

BUFx12f_ASAP7_75t_L g2113 ( 
.A(n_2062),
.Y(n_2113)
);

CKINVDCx6p67_ASAP7_75t_R g2114 ( 
.A(n_2075),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2069),
.Y(n_2115)
);

INVx6_ASAP7_75t_L g2116 ( 
.A(n_2082),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2045),
.B(n_2010),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_SL g2118 ( 
.A1(n_2082),
.A2(n_2016),
.B1(n_1842),
.B2(n_2009),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_2058),
.Y(n_2119)
);

AOI21xp33_ASAP7_75t_L g2120 ( 
.A1(n_2071),
.A2(n_2006),
.B(n_2020),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2072),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2057),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_2031),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2030),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2042),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2087),
.A2(n_1919),
.B1(n_1990),
.B2(n_1899),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2077),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2074),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2074),
.Y(n_2129)
);

CKINVDCx20_ASAP7_75t_R g2130 ( 
.A(n_2079),
.Y(n_2130)
);

CKINVDCx11_ASAP7_75t_R g2131 ( 
.A(n_2075),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_2087),
.A2(n_1942),
.B1(n_1955),
.B2(n_1940),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2128),
.B(n_2060),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2107),
.A2(n_2037),
.B1(n_2050),
.B2(n_2067),
.Y(n_2134)
);

A2O1A1Ixp33_ASAP7_75t_L g2135 ( 
.A1(n_2118),
.A2(n_2040),
.B(n_2070),
.C(n_2065),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_2103),
.A2(n_2038),
.B(n_2090),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2105),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_2101),
.B(n_2086),
.Y(n_2138)
);

AOI21x1_ASAP7_75t_SL g2139 ( 
.A1(n_2117),
.A2(n_2068),
.B(n_2088),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_2126),
.A2(n_2067),
.B1(n_1997),
.B2(n_2064),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2122),
.B(n_2041),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2105),
.Y(n_2142)
);

OAI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2095),
.A2(n_2110),
.B1(n_2108),
.B2(n_2111),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2128),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2115),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2111),
.A2(n_2085),
.B1(n_2092),
.B2(n_2063),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2101),
.B(n_2081),
.Y(n_2147)
);

OAI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_2114),
.A2(n_2063),
.B1(n_2002),
.B2(n_2053),
.Y(n_2148)
);

OA21x2_ASAP7_75t_L g2149 ( 
.A1(n_2129),
.A2(n_1958),
.B(n_2034),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2129),
.B(n_2056),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2123),
.B(n_2051),
.Y(n_2151)
);

O2A1O1Ixp5_ASAP7_75t_L g2152 ( 
.A1(n_2120),
.A2(n_2059),
.B(n_2089),
.C(n_2048),
.Y(n_2152)
);

O2A1O1Ixp5_ASAP7_75t_L g2153 ( 
.A1(n_2125),
.A2(n_2124),
.B(n_2121),
.C(n_2098),
.Y(n_2153)
);

A2O1A1Ixp33_ASAP7_75t_L g2154 ( 
.A1(n_2132),
.A2(n_2091),
.B(n_2078),
.C(n_1960),
.Y(n_2154)
);

INVxp33_ASAP7_75t_L g2155 ( 
.A(n_2131),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2149),
.Y(n_2156)
);

AND2x4_ASAP7_75t_SL g2157 ( 
.A(n_2138),
.B(n_2114),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2137),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_2138),
.B(n_2104),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_2144),
.B(n_2151),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2133),
.B(n_2123),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2150),
.B(n_2109),
.Y(n_2162)
);

CKINVDCx16_ASAP7_75t_R g2163 ( 
.A(n_2143),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2162),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2162),
.Y(n_2165)
);

OR2x6_ASAP7_75t_L g2166 ( 
.A(n_2159),
.B(n_2096),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2161),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2161),
.B(n_2136),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2160),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2168),
.A2(n_2163),
.B1(n_2156),
.B2(n_2140),
.Y(n_2170)
);

INVxp33_ASAP7_75t_SL g2171 ( 
.A(n_2167),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2165),
.A2(n_2156),
.B1(n_2149),
.B2(n_2134),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2166),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2166),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_2169),
.B(n_2160),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2164),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2164),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2167),
.B(n_2160),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2170),
.A2(n_2135),
.B1(n_2171),
.B2(n_2172),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2178),
.B(n_2175),
.Y(n_2180)
);

AOI33xp33_ASAP7_75t_L g2181 ( 
.A1(n_2174),
.A2(n_2157),
.A3(n_2135),
.B1(n_2158),
.B2(n_2159),
.B3(n_2141),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2178),
.B(n_2175),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2171),
.A2(n_2148),
.B1(n_2146),
.B2(n_2154),
.Y(n_2183)
);

AND2x6_ASAP7_75t_SL g2184 ( 
.A(n_2175),
.B(n_2032),
.Y(n_2184)
);

OAI31xp33_ASAP7_75t_SL g2185 ( 
.A1(n_2176),
.A2(n_2159),
.A3(n_2131),
.B(n_2113),
.Y(n_2185)
);

OR2x6_ASAP7_75t_L g2186 ( 
.A(n_2173),
.B(n_2096),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2176),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2175),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_2177),
.A2(n_2153),
.B(n_2158),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2188),
.B(n_2177),
.Y(n_2190)
);

INVxp67_ASAP7_75t_SL g2191 ( 
.A(n_2183),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2187),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2180),
.B(n_2173),
.Y(n_2193)
);

INVx1_ASAP7_75t_SL g2194 ( 
.A(n_2186),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_2182),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2186),
.B(n_2157),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2186),
.B(n_2155),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_2184),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2195),
.B(n_2130),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2196),
.B(n_2197),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2193),
.B(n_2179),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2194),
.B(n_2185),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2199),
.B(n_2198),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2199),
.B(n_2198),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2201),
.B(n_2191),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2200),
.B(n_2194),
.Y(n_2206)
);

HB1xp67_ASAP7_75t_L g2207 ( 
.A(n_2206),
.Y(n_2207)
);

OAI33xp33_ASAP7_75t_L g2208 ( 
.A1(n_2203),
.A2(n_2192),
.A3(n_2190),
.B1(n_2179),
.B2(n_2202),
.B3(n_2200),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_SL g2209 ( 
.A1(n_2204),
.A2(n_2102),
.B1(n_2155),
.B2(n_2130),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2205),
.A2(n_2189),
.B1(n_2113),
.B2(n_2181),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2203),
.B(n_2144),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2206),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2207),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2212),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2210),
.B(n_2185),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2211),
.B(n_2106),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2209),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_2208),
.A2(n_2149),
.B1(n_2078),
.B2(n_2094),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2207),
.B(n_2106),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2207),
.B(n_2096),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2212),
.B(n_2147),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2207),
.B(n_2096),
.Y(n_2222)
);

OAI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2213),
.A2(n_2152),
.B(n_2028),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2214),
.A2(n_2154),
.B1(n_2094),
.B2(n_2112),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2220),
.A2(n_1859),
.B(n_1853),
.Y(n_2225)
);

O2A1O1Ixp33_ASAP7_75t_L g2226 ( 
.A1(n_2217),
.A2(n_1876),
.B(n_1908),
.C(n_1888),
.Y(n_2226)
);

INVxp67_ASAP7_75t_L g2227 ( 
.A(n_2222),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2219),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2221),
.B(n_2099),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2221),
.B(n_2147),
.Y(n_2230)
);

OA21x2_ASAP7_75t_L g2231 ( 
.A1(n_2218),
.A2(n_1992),
.B(n_1915),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2216),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2216),
.B(n_2142),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2215),
.A2(n_2049),
.B1(n_2116),
.B2(n_2073),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2213),
.Y(n_2235)
);

AOI322xp5_ASAP7_75t_L g2236 ( 
.A1(n_2235),
.A2(n_2016),
.A3(n_1893),
.B1(n_1914),
.B2(n_2029),
.C1(n_2049),
.C2(n_2025),
.Y(n_2236)
);

OAI21xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2227),
.A2(n_1798),
.B(n_1871),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2230),
.B(n_2119),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2228),
.B(n_2119),
.Y(n_2239)
);

AOI21xp33_ASAP7_75t_L g2240 ( 
.A1(n_2232),
.A2(n_1908),
.B(n_1888),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2229),
.B(n_2100),
.Y(n_2241)
);

AOI221xp5_ASAP7_75t_L g2242 ( 
.A1(n_2223),
.A2(n_1943),
.B1(n_1945),
.B2(n_2145),
.C(n_2115),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2231),
.A2(n_2116),
.B1(n_2073),
.B2(n_2104),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2225),
.B(n_2036),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2233),
.B(n_175),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2226),
.B(n_176),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2234),
.A2(n_2116),
.B1(n_2080),
.B2(n_2104),
.Y(n_2247)
);

NOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2231),
.B(n_2224),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2235),
.A2(n_2116),
.B1(n_2084),
.B2(n_2083),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_2227),
.A2(n_1994),
.B(n_1956),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2243),
.A2(n_1834),
.B1(n_1864),
.B2(n_1803),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2248),
.B(n_177),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2239),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2245),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2241),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2246),
.B(n_1864),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2238),
.B(n_177),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2244),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2240),
.B(n_2237),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_2249),
.B(n_1864),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2242),
.A2(n_2017),
.B1(n_2127),
.B2(n_1803),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2247),
.B(n_178),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_2250),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2236),
.Y(n_2264)
);

AND3x4_ASAP7_75t_L g2265 ( 
.A(n_2253),
.B(n_2139),
.C(n_178),
.Y(n_2265)
);

NOR3xp33_ASAP7_75t_L g2266 ( 
.A(n_2252),
.B(n_2024),
.C(n_2019),
.Y(n_2266)
);

NOR3x1_ASAP7_75t_L g2267 ( 
.A(n_2257),
.B(n_179),
.C(n_180),
.Y(n_2267)
);

NOR2x1p5_ASAP7_75t_L g2268 ( 
.A(n_2264),
.B(n_1834),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2255),
.Y(n_2269)
);

OAI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2258),
.A2(n_1969),
.B(n_1965),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2254),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2263),
.B(n_179),
.Y(n_2272)
);

NOR3xp33_ASAP7_75t_L g2273 ( 
.A(n_2256),
.B(n_1963),
.C(n_2001),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2263),
.B(n_180),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2262),
.B(n_1885),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2259),
.Y(n_2276)
);

NOR2x1_ASAP7_75t_L g2277 ( 
.A(n_2260),
.B(n_181),
.Y(n_2277)
);

NOR3xp33_ASAP7_75t_L g2278 ( 
.A(n_2251),
.B(n_2021),
.C(n_2003),
.Y(n_2278)
);

CKINVDCx20_ASAP7_75t_R g2279 ( 
.A(n_2261),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_SL g2280 ( 
.A1(n_2264),
.A2(n_181),
.B(n_182),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2252),
.B(n_182),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_L g2282 ( 
.A(n_2252),
.B(n_184),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2257),
.A2(n_185),
.B(n_186),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2252),
.Y(n_2284)
);

NAND3xp33_ASAP7_75t_L g2285 ( 
.A(n_2252),
.B(n_1828),
.C(n_185),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2252),
.Y(n_2286)
);

AOI211xp5_ASAP7_75t_L g2287 ( 
.A1(n_2280),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2267),
.B(n_187),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_SL g2289 ( 
.A(n_2269),
.B(n_189),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2272),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2284),
.B(n_189),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_2276),
.A2(n_2127),
.B1(n_2097),
.B2(n_1961),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2282),
.B(n_190),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2283),
.B(n_191),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2274),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2286),
.B(n_191),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2271),
.A2(n_1985),
.B(n_1967),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2277),
.B(n_192),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2281),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2285),
.B(n_192),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2268),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2265),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2270),
.B(n_193),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2275),
.B(n_194),
.Y(n_2304)
);

AOI211xp5_ASAP7_75t_L g2305 ( 
.A1(n_2278),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2279),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2266),
.B(n_2273),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2269),
.B(n_196),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_2269),
.A2(n_197),
.B(n_198),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_L g2310 ( 
.A(n_2267),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2267),
.Y(n_2311)
);

NAND4xp25_ASAP7_75t_SL g2312 ( 
.A(n_2271),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2267),
.Y(n_2313)
);

INVx1_ASAP7_75t_SL g2314 ( 
.A(n_2281),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2267),
.B(n_204),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2267),
.Y(n_2316)
);

NAND5xp2_ASAP7_75t_L g2317 ( 
.A(n_2280),
.B(n_208),
.C(n_205),
.D(n_207),
.E(n_210),
.Y(n_2317)
);

O2A1O1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2280),
.A2(n_210),
.B(n_207),
.C(n_208),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2267),
.Y(n_2319)
);

NOR3xp33_ASAP7_75t_L g2320 ( 
.A(n_2276),
.B(n_211),
.C(n_212),
.Y(n_2320)
);

OAI22xp33_ASAP7_75t_SL g2321 ( 
.A1(n_2284),
.A2(n_2097),
.B1(n_1957),
.B2(n_2093),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_L g2322 ( 
.A(n_2280),
.B(n_211),
.C(n_212),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2269),
.Y(n_2323)
);

NOR3xp33_ASAP7_75t_L g2324 ( 
.A(n_2306),
.B(n_213),
.C(n_214),
.Y(n_2324)
);

NOR4xp75_ASAP7_75t_L g2325 ( 
.A(n_2288),
.B(n_215),
.C(n_213),
.D(n_214),
.Y(n_2325)
);

AOI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2323),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_2326)
);

NOR2x1_ASAP7_75t_L g2327 ( 
.A(n_2312),
.B(n_216),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2308),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_SL g2329 ( 
.A1(n_2315),
.A2(n_217),
.B(n_218),
.Y(n_2329)
);

AOI211xp5_ASAP7_75t_L g2330 ( 
.A1(n_2302),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_L g2331 ( 
.A(n_2310),
.B(n_222),
.C(n_219),
.D(n_221),
.Y(n_2331)
);

NAND3xp33_ASAP7_75t_L g2332 ( 
.A(n_2289),
.B(n_221),
.C(n_222),
.Y(n_2332)
);

NOR3xp33_ASAP7_75t_L g2333 ( 
.A(n_2290),
.B(n_223),
.C(n_224),
.Y(n_2333)
);

NAND3xp33_ASAP7_75t_L g2334 ( 
.A(n_2311),
.B(n_223),
.C(n_225),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2317),
.B(n_225),
.Y(n_2335)
);

NAND4xp25_ASAP7_75t_L g2336 ( 
.A(n_2313),
.B(n_228),
.C(n_226),
.D(n_227),
.Y(n_2336)
);

NOR3x1_ASAP7_75t_L g2337 ( 
.A(n_2322),
.B(n_226),
.C(n_227),
.Y(n_2337)
);

NAND3xp33_ASAP7_75t_L g2338 ( 
.A(n_2316),
.B(n_229),
.C(n_230),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2319),
.B(n_229),
.Y(n_2339)
);

AOI211xp5_ASAP7_75t_L g2340 ( 
.A1(n_2318),
.A2(n_233),
.B(n_230),
.C(n_232),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2303),
.A2(n_232),
.B(n_233),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2314),
.B(n_234),
.Y(n_2342)
);

NOR3xp33_ASAP7_75t_SL g2343 ( 
.A(n_2298),
.B(n_234),
.C(n_235),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2320),
.B(n_235),
.C(n_236),
.Y(n_2344)
);

NAND3xp33_ASAP7_75t_L g2345 ( 
.A(n_2287),
.B(n_236),
.C(n_237),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_SL g2346 ( 
.A(n_2291),
.B(n_238),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_SL g2347 ( 
.A(n_2293),
.B(n_238),
.Y(n_2347)
);

NAND3xp33_ASAP7_75t_L g2348 ( 
.A(n_2287),
.B(n_239),
.C(n_240),
.Y(n_2348)
);

NAND3xp33_ASAP7_75t_L g2349 ( 
.A(n_2299),
.B(n_239),
.C(n_241),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2304),
.B(n_242),
.Y(n_2350)
);

NAND3xp33_ASAP7_75t_SL g2351 ( 
.A(n_2309),
.B(n_243),
.C(n_244),
.Y(n_2351)
);

NOR3xp33_ASAP7_75t_L g2352 ( 
.A(n_2295),
.B(n_243),
.C(n_245),
.Y(n_2352)
);

AOI21xp33_ASAP7_75t_SL g2353 ( 
.A1(n_2294),
.A2(n_245),
.B(n_246),
.Y(n_2353)
);

OAI211xp5_ASAP7_75t_L g2354 ( 
.A1(n_2305),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2296),
.Y(n_2355)
);

AND4x1_ASAP7_75t_L g2356 ( 
.A(n_2301),
.B(n_250),
.C(n_248),
.D(n_249),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2331),
.B(n_2300),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2339),
.A2(n_2307),
.B(n_2297),
.Y(n_2358)
);

NAND3xp33_ASAP7_75t_L g2359 ( 
.A(n_2347),
.B(n_2292),
.C(n_2321),
.Y(n_2359)
);

NAND4xp25_ASAP7_75t_L g2360 ( 
.A(n_2337),
.B(n_251),
.C(n_249),
.D(n_250),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_L g2361 ( 
.A(n_2346),
.B(n_251),
.C(n_252),
.Y(n_2361)
);

NAND3x1_ASAP7_75t_L g2362 ( 
.A(n_2324),
.B(n_253),
.C(n_255),
.Y(n_2362)
);

AOI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_2335),
.A2(n_2007),
.B1(n_2055),
.B2(n_2023),
.Y(n_2363)
);

NOR2x1_ASAP7_75t_L g2364 ( 
.A(n_2336),
.B(n_253),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_L g2365 ( 
.A(n_2328),
.B(n_255),
.C(n_256),
.Y(n_2365)
);

OR3x1_ASAP7_75t_L g2366 ( 
.A(n_2351),
.B(n_256),
.C(n_258),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2356),
.B(n_258),
.Y(n_2367)
);

NAND4xp25_ASAP7_75t_L g2368 ( 
.A(n_2327),
.B(n_261),
.C(n_259),
.D(n_260),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2343),
.B(n_2350),
.Y(n_2369)
);

NOR2x1_ASAP7_75t_L g2370 ( 
.A(n_2334),
.B(n_260),
.Y(n_2370)
);

OAI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2338),
.A2(n_2055),
.B1(n_263),
.B2(n_261),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2353),
.B(n_262),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2329),
.B(n_262),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2355),
.A2(n_2055),
.B1(n_1935),
.B2(n_266),
.Y(n_2374)
);

NAND4xp25_ASAP7_75t_L g2375 ( 
.A(n_2340),
.B(n_2345),
.C(n_2348),
.D(n_2344),
.Y(n_2375)
);

OAI211xp5_ASAP7_75t_SL g2376 ( 
.A1(n_2341),
.A2(n_2342),
.B(n_2326),
.C(n_2330),
.Y(n_2376)
);

NOR3x1_ASAP7_75t_L g2377 ( 
.A(n_2349),
.B(n_264),
.C(n_265),
.Y(n_2377)
);

NAND4xp25_ASAP7_75t_L g2378 ( 
.A(n_2332),
.B(n_267),
.C(n_264),
.D(n_266),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2333),
.B(n_268),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2352),
.B(n_268),
.Y(n_2380)
);

NOR3xp33_ASAP7_75t_L g2381 ( 
.A(n_2354),
.B(n_2325),
.C(n_269),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2327),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2335),
.B(n_269),
.Y(n_2383)
);

OAI211xp5_ASAP7_75t_SL g2384 ( 
.A1(n_2329),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_2384)
);

AOI211xp5_ASAP7_75t_L g2385 ( 
.A1(n_2335),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2385)
);

NOR3x1_ASAP7_75t_L g2386 ( 
.A(n_2334),
.B(n_273),
.C(n_274),
.Y(n_2386)
);

O2A1O1Ixp33_ASAP7_75t_L g2387 ( 
.A1(n_2339),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2335),
.B(n_276),
.Y(n_2388)
);

OAI21xp33_ASAP7_75t_SL g2389 ( 
.A1(n_2327),
.A2(n_277),
.B(n_278),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_L g2390 ( 
.A(n_2347),
.B(n_277),
.C(n_279),
.Y(n_2390)
);

NAND4xp25_ASAP7_75t_L g2391 ( 
.A(n_2337),
.B(n_281),
.C(n_279),
.D(n_280),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2350),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2335),
.B(n_280),
.Y(n_2393)
);

NAND4xp25_ASAP7_75t_L g2394 ( 
.A(n_2337),
.B(n_284),
.C(n_282),
.D(n_283),
.Y(n_2394)
);

NOR2x1_ASAP7_75t_L g2395 ( 
.A(n_2336),
.B(n_282),
.Y(n_2395)
);

OAI22xp33_ASAP7_75t_L g2396 ( 
.A1(n_2339),
.A2(n_287),
.B1(n_284),
.B2(n_286),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2356),
.B(n_287),
.Y(n_2397)
);

OAI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2327),
.A2(n_288),
.B(n_289),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2335),
.B(n_289),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2339),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_2400)
);

AOI211xp5_ASAP7_75t_L g2401 ( 
.A1(n_2335),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_2401)
);

AOI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2331),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.C(n_296),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2327),
.Y(n_2403)
);

NAND4xp25_ASAP7_75t_SL g2404 ( 
.A(n_2340),
.B(n_297),
.C(n_293),
.D(n_296),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2356),
.B(n_298),
.Y(n_2405)
);

AOI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2339),
.A2(n_299),
.B(n_300),
.Y(n_2406)
);

AOI221x1_ASAP7_75t_L g2407 ( 
.A1(n_2339),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.C(n_303),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2382),
.B(n_301),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2366),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2392),
.B(n_302),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2369),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2403),
.Y(n_2412)
);

AOI222xp33_ASAP7_75t_L g2413 ( 
.A1(n_2389),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.C1(n_307),
.C2(n_308),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2383),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_2414)
);

AOI31xp33_ASAP7_75t_L g2415 ( 
.A1(n_2385),
.A2(n_2401),
.A3(n_2388),
.B(n_2399),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2364),
.B(n_2395),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2398),
.B(n_308),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2373),
.B(n_309),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2370),
.B(n_309),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2362),
.Y(n_2420)
);

OAI211xp5_ASAP7_75t_SL g2421 ( 
.A1(n_2358),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_2421)
);

A2O1A1Ixp33_ASAP7_75t_L g2422 ( 
.A1(n_2372),
.A2(n_314),
.B(n_310),
.C(n_313),
.Y(n_2422)
);

INVx1_ASAP7_75t_SL g2423 ( 
.A(n_2357),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2368),
.B(n_313),
.Y(n_2424)
);

OAI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2367),
.A2(n_314),
.B(n_316),
.Y(n_2425)
);

NOR2xp67_ASAP7_75t_L g2426 ( 
.A(n_2404),
.B(n_316),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_2381),
.B(n_317),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2397),
.Y(n_2428)
);

NAND4xp75_ASAP7_75t_L g2429 ( 
.A(n_2386),
.B(n_317),
.C(n_318),
.D(n_319),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_R g2430 ( 
.A(n_2393),
.B(n_318),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2405),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2387),
.A2(n_319),
.B(n_320),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2361),
.B(n_320),
.Y(n_2433)
);

NAND2xp33_ASAP7_75t_R g2434 ( 
.A(n_2379),
.B(n_321),
.Y(n_2434)
);

NOR2x1p5_ASAP7_75t_L g2435 ( 
.A(n_2360),
.B(n_321),
.Y(n_2435)
);

INVx2_ASAP7_75t_SL g2436 ( 
.A(n_2390),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2377),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2407),
.Y(n_2438)
);

CKINVDCx20_ASAP7_75t_R g2439 ( 
.A(n_2380),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2376),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_2440)
);

INVx1_ASAP7_75t_SL g2441 ( 
.A(n_2406),
.Y(n_2441)
);

OAI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2374),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_2442)
);

NOR2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2391),
.B(n_326),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2365),
.B(n_326),
.Y(n_2444)
);

CKINVDCx16_ASAP7_75t_R g2445 ( 
.A(n_2400),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2384),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_L g2447 ( 
.A(n_2394),
.Y(n_2447)
);

AOI221xp5_ASAP7_75t_L g2448 ( 
.A1(n_2371),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.C(n_330),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2378),
.Y(n_2449)
);

OAI22xp5_ASAP7_75t_L g2450 ( 
.A1(n_2359),
.A2(n_327),
.B1(n_328),
.B2(n_330),
.Y(n_2450)
);

OAI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2402),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_R g2452 ( 
.A(n_2396),
.B(n_331),
.Y(n_2452)
);

O2A1O1Ixp5_ASAP7_75t_SL g2453 ( 
.A1(n_2375),
.A2(n_332),
.B(n_334),
.C(n_335),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_2363),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2409),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2423),
.B(n_336),
.Y(n_2456)
);

AND2x2_ASAP7_75t_SL g2457 ( 
.A(n_2412),
.B(n_2420),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2438),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2419),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_2419),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2416),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2411),
.B(n_2437),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2408),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2408),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2428),
.B(n_336),
.Y(n_2465)
);

NOR2x1_ASAP7_75t_L g2466 ( 
.A(n_2410),
.B(n_337),
.Y(n_2466)
);

NAND4xp75_ASAP7_75t_L g2467 ( 
.A(n_2427),
.B(n_337),
.C(n_339),
.D(n_340),
.Y(n_2467)
);

NOR2x1_ASAP7_75t_L g2468 ( 
.A(n_2431),
.B(n_339),
.Y(n_2468)
);

NAND2x1_ASAP7_75t_SL g2469 ( 
.A(n_2447),
.B(n_340),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2429),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2435),
.Y(n_2471)
);

NAND2xp33_ASAP7_75t_L g2472 ( 
.A(n_2450),
.B(n_341),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2434),
.B(n_341),
.C(n_342),
.Y(n_2473)
);

OAI22x1_ASAP7_75t_L g2474 ( 
.A1(n_2414),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2441),
.B(n_343),
.Y(n_2475)
);

NOR2x1_ASAP7_75t_L g2476 ( 
.A(n_2418),
.B(n_345),
.Y(n_2476)
);

NAND4xp75_ASAP7_75t_L g2477 ( 
.A(n_2425),
.B(n_346),
.C(n_347),
.D(n_348),
.Y(n_2477)
);

NAND4xp75_ASAP7_75t_L g2478 ( 
.A(n_2426),
.B(n_347),
.C(n_348),
.D(n_349),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2443),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2446),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2417),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2424),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2445),
.B(n_350),
.Y(n_2483)
);

OR2x2_ASAP7_75t_L g2484 ( 
.A(n_2444),
.B(n_350),
.Y(n_2484)
);

NOR2x1_ASAP7_75t_L g2485 ( 
.A(n_2421),
.B(n_351),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2417),
.Y(n_2486)
);

XOR2xp5_ASAP7_75t_L g2487 ( 
.A(n_2439),
.B(n_351),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2430),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2433),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2449),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_2490)
);

HB1xp67_ASAP7_75t_L g2491 ( 
.A(n_2433),
.Y(n_2491)
);

NOR2x1_ASAP7_75t_L g2492 ( 
.A(n_2422),
.B(n_352),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2457),
.Y(n_2493)
);

NAND3x1_ASAP7_75t_L g2494 ( 
.A(n_2458),
.B(n_2440),
.C(n_2432),
.Y(n_2494)
);

NOR3xp33_ASAP7_75t_L g2495 ( 
.A(n_2461),
.B(n_2415),
.C(n_2436),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2462),
.B(n_2455),
.Y(n_2496)
);

NOR3xp33_ASAP7_75t_SL g2497 ( 
.A(n_2489),
.B(n_2454),
.C(n_2442),
.Y(n_2497)
);

OR2x2_ASAP7_75t_L g2498 ( 
.A(n_2460),
.B(n_2451),
.Y(n_2498)
);

NOR3xp33_ASAP7_75t_L g2499 ( 
.A(n_2464),
.B(n_2448),
.C(n_2452),
.Y(n_2499)
);

NOR5xp2_ASAP7_75t_L g2500 ( 
.A(n_2491),
.B(n_2413),
.C(n_2453),
.D(n_356),
.E(n_357),
.Y(n_2500)
);

OAI222xp33_ASAP7_75t_R g2501 ( 
.A1(n_2488),
.A2(n_2479),
.B1(n_2471),
.B2(n_2480),
.C1(n_2486),
.C2(n_2482),
.Y(n_2501)
);

OA22x2_ASAP7_75t_L g2502 ( 
.A1(n_2456),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.Y(n_2502)
);

AND5x1_ASAP7_75t_L g2503 ( 
.A(n_2490),
.B(n_355),
.C(n_357),
.D(n_358),
.E(n_359),
.Y(n_2503)
);

NOR4xp75_ASAP7_75t_L g2504 ( 
.A(n_2469),
.B(n_359),
.C(n_360),
.D(n_361),
.Y(n_2504)
);

NAND4xp25_ASAP7_75t_L g2505 ( 
.A(n_2473),
.B(n_360),
.C(n_361),
.D(n_362),
.Y(n_2505)
);

OAI211xp5_ASAP7_75t_L g2506 ( 
.A1(n_2483),
.A2(n_362),
.B(n_363),
.C(n_364),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2475),
.B(n_364),
.Y(n_2507)
);

NAND4xp75_ASAP7_75t_L g2508 ( 
.A(n_2476),
.B(n_365),
.C(n_366),
.D(n_367),
.Y(n_2508)
);

INVx5_ASAP7_75t_L g2509 ( 
.A(n_2463),
.Y(n_2509)
);

NOR2x1_ASAP7_75t_L g2510 ( 
.A(n_2478),
.B(n_366),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2459),
.B(n_368),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_L g2512 ( 
.A(n_2463),
.B(n_369),
.C(n_370),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_SL g2513 ( 
.A(n_2467),
.B(n_370),
.C(n_371),
.Y(n_2513)
);

NOR2x1p5_ASAP7_75t_L g2514 ( 
.A(n_2477),
.B(n_372),
.Y(n_2514)
);

NAND4xp25_ASAP7_75t_L g2515 ( 
.A(n_2468),
.B(n_372),
.C(n_373),
.D(n_374),
.Y(n_2515)
);

AND3x4_ASAP7_75t_L g2516 ( 
.A(n_2485),
.B(n_373),
.C(n_375),
.Y(n_2516)
);

XNOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2466),
.B(n_375),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2481),
.B(n_376),
.C(n_377),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2484),
.B(n_376),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_SL g2520 ( 
.A(n_2470),
.B(n_379),
.C(n_380),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2493),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_2509),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_2509),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2496),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2509),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2497),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2498),
.Y(n_2527)
);

OR2x2_ASAP7_75t_L g2528 ( 
.A(n_2519),
.B(n_2477),
.Y(n_2528)
);

INVx1_ASAP7_75t_SL g2529 ( 
.A(n_2517),
.Y(n_2529)
);

NAND2xp33_ASAP7_75t_L g2530 ( 
.A(n_2495),
.B(n_2487),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_2499),
.A2(n_2472),
.B(n_2474),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2507),
.B(n_2465),
.Y(n_2532)
);

HB1xp67_ASAP7_75t_L g2533 ( 
.A(n_2504),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2501),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2510),
.B(n_2492),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2511),
.B(n_379),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2516),
.Y(n_2537)
);

HB1xp67_ASAP7_75t_L g2538 ( 
.A(n_2514),
.Y(n_2538)
);

CKINVDCx20_ASAP7_75t_R g2539 ( 
.A(n_2513),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2502),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2523),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2534),
.Y(n_2542)
);

AOI32xp33_ASAP7_75t_L g2543 ( 
.A1(n_2522),
.A2(n_2500),
.A3(n_2494),
.B1(n_2503),
.B2(n_2505),
.Y(n_2543)
);

AOI322xp5_ASAP7_75t_L g2544 ( 
.A1(n_2521),
.A2(n_2520),
.A3(n_2518),
.B1(n_2515),
.B2(n_2508),
.C1(n_2506),
.C2(n_2512),
.Y(n_2544)
);

AOI221xp5_ASAP7_75t_L g2545 ( 
.A1(n_2524),
.A2(n_380),
.B1(n_381),
.B2(n_383),
.C(n_384),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2525),
.Y(n_2546)
);

OAI211xp5_ASAP7_75t_SL g2547 ( 
.A1(n_2530),
.A2(n_384),
.B(n_385),
.C(n_386),
.Y(n_2547)
);

OAI221xp5_ASAP7_75t_L g2548 ( 
.A1(n_2526),
.A2(n_385),
.B1(n_387),
.B2(n_388),
.C(n_389),
.Y(n_2548)
);

AOI322xp5_ASAP7_75t_L g2549 ( 
.A1(n_2529),
.A2(n_388),
.A3(n_389),
.B1(n_390),
.B2(n_391),
.C1(n_392),
.C2(n_393),
.Y(n_2549)
);

AOI322xp5_ASAP7_75t_L g2550 ( 
.A1(n_2538),
.A2(n_394),
.A3(n_395),
.B1(n_396),
.B2(n_397),
.C1(n_398),
.C2(n_399),
.Y(n_2550)
);

AOI221xp5_ASAP7_75t_L g2551 ( 
.A1(n_2527),
.A2(n_394),
.B1(n_396),
.B2(n_399),
.C(n_400),
.Y(n_2551)
);

AOI322xp5_ASAP7_75t_L g2552 ( 
.A1(n_2533),
.A2(n_400),
.A3(n_401),
.B1(n_402),
.B2(n_403),
.C1(n_404),
.C2(n_405),
.Y(n_2552)
);

NOR2x1_ASAP7_75t_L g2553 ( 
.A(n_2535),
.B(n_401),
.Y(n_2553)
);

OAI221xp5_ASAP7_75t_L g2554 ( 
.A1(n_2537),
.A2(n_402),
.B1(n_405),
.B2(n_406),
.C(n_407),
.Y(n_2554)
);

A2O1A1Ixp33_ASAP7_75t_L g2555 ( 
.A1(n_2531),
.A2(n_406),
.B(n_407),
.C(n_408),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2539),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_2556)
);

AO22x2_ASAP7_75t_L g2557 ( 
.A1(n_2541),
.A2(n_2531),
.B1(n_2532),
.B2(n_2528),
.Y(n_2557)
);

OAI22x1_ASAP7_75t_L g2558 ( 
.A1(n_2546),
.A2(n_2540),
.B1(n_2536),
.B2(n_412),
.Y(n_2558)
);

OAI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2542),
.A2(n_409),
.B1(n_411),
.B2(n_413),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2543),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.Y(n_2560)
);

AO22x2_ASAP7_75t_SL g2561 ( 
.A1(n_2553),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2548),
.Y(n_2562)
);

AO22x2_ASAP7_75t_L g2563 ( 
.A1(n_2544),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_2563)
);

NAND4xp25_ASAP7_75t_SL g2564 ( 
.A(n_2561),
.B(n_2555),
.C(n_2551),
.D(n_2545),
.Y(n_2564)
);

AND4x1_ASAP7_75t_L g2565 ( 
.A(n_2557),
.B(n_2556),
.C(n_2547),
.D(n_2554),
.Y(n_2565)
);

OAI21x1_ASAP7_75t_L g2566 ( 
.A1(n_2559),
.A2(n_2552),
.B(n_2549),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2558),
.Y(n_2567)
);

OAI222xp33_ASAP7_75t_L g2568 ( 
.A1(n_2562),
.A2(n_2550),
.B1(n_421),
.B2(n_422),
.C1(n_423),
.C2(n_425),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2567),
.A2(n_2563),
.B1(n_2564),
.B2(n_2566),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2565),
.A2(n_2560),
.B(n_421),
.Y(n_2570)
);

NOR3xp33_ASAP7_75t_L g2571 ( 
.A(n_2568),
.B(n_420),
.C(n_422),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2569),
.B(n_423),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2570),
.A2(n_425),
.B(n_427),
.Y(n_2573)
);

OAI22xp33_ASAP7_75t_L g2574 ( 
.A1(n_2571),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2572),
.B(n_428),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2573),
.B(n_430),
.Y(n_2576)
);

OAI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2575),
.A2(n_2574),
.B(n_431),
.Y(n_2577)
);

A2O1A1Ixp33_ASAP7_75t_L g2578 ( 
.A1(n_2576),
.A2(n_430),
.B(n_431),
.C(n_505),
.Y(n_2578)
);

AOI22xp5_ASAP7_75t_L g2579 ( 
.A1(n_2577),
.A2(n_506),
.B1(n_507),
.B2(n_509),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2578),
.A2(n_510),
.B1(n_512),
.B2(n_514),
.Y(n_2580)
);

OAI21xp33_ASAP7_75t_L g2581 ( 
.A1(n_2580),
.A2(n_515),
.B(n_518),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2581),
.B(n_2579),
.Y(n_2582)
);

AOI221x1_ASAP7_75t_L g2583 ( 
.A1(n_2582),
.A2(n_519),
.B1(n_522),
.B2(n_523),
.C(n_524),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2583),
.A2(n_525),
.B1(n_526),
.B2(n_527),
.Y(n_2584)
);

AOI211xp5_ASAP7_75t_L g2585 ( 
.A1(n_2584),
.A2(n_530),
.B(n_531),
.C(n_532),
.Y(n_2585)
);


endmodule