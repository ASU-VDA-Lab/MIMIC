module fake_ibex_1124_n_921 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_921);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_921;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_179;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_905;
wire n_410;
wire n_762;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_890;
wire n_816;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_11),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_87),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_78),
.Y(n_182)
);

INVxp33_ASAP7_75t_SL g183 ( 
.A(n_66),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_49),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_53),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_26),
.Y(n_191)
);

INVxp33_ASAP7_75t_SL g192 ( 
.A(n_62),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_35),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_15),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_13),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_17),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_39),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_37),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_168),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_14),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_85),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_52),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_54),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_139),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_84),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_89),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_97),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_48),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_31),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_79),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_60),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_71),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_169),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_110),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_105),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_121),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_115),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_129),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_81),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_122),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_20),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_67),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_42),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_73),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_132),
.B(n_46),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_36),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_98),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_4),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_59),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_151),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_92),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_36),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_108),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_111),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_76),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_96),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_86),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_175),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_154),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_16),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_61),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_114),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_65),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_0),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_0),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_210),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_193),
.B(n_1),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_2),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_44),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_215),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_2),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_3),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_178),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_199),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_185),
.B(n_7),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_203),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_185),
.B(n_9),
.Y(n_312)
);

XNOR2x2_ASAP7_75t_L g313 ( 
.A(n_214),
.B(n_10),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_245),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_242),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_189),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_245),
.B(n_266),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_195),
.Y(n_318)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_189),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_199),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_197),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g323 ( 
.A(n_188),
.B(n_47),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_184),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_195),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

BUFx8_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_15),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_186),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_187),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_18),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_176),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_190),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_194),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_19),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_195),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_196),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_234),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_198),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_183),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_202),
.B(n_21),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_204),
.B(n_23),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_180),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_234),
.B(n_23),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_206),
.Y(n_357)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_234),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_207),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_212),
.Y(n_360)
);

AOI22x1_ASAP7_75t_SL g361 ( 
.A1(n_197),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_216),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_182),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_349),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_301),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_304),
.B(n_205),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_306),
.A2(n_183),
.B1(n_192),
.B2(n_287),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_301),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_182),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_323),
.A2(n_218),
.B1(n_222),
.B2(n_250),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_191),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_345),
.Y(n_385)
);

AO22x1_ASAP7_75t_L g386 ( 
.A1(n_332),
.A2(n_192),
.B1(n_224),
.B2(n_284),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_310),
.B(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_R g394 ( 
.A(n_340),
.B(n_201),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_291),
.B(n_211),
.C(n_208),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_292),
.B(n_311),
.C(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_345),
.B(n_252),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_306),
.A2(n_289),
.B1(n_288),
.B2(n_228),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_254),
.Y(n_402)
);

CKINVDCx11_ASAP7_75t_R g403 ( 
.A(n_322),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_283),
.B1(n_255),
.B2(n_261),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_308),
.B(n_209),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_323),
.A2(n_209),
.B1(n_218),
.B2(n_262),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_319),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_324),
.B(n_223),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_317),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

OR2x6_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_222),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_264),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_293),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_293),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_319),
.B(n_227),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_354),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_294),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_334),
.B(n_225),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_298),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_334),
.B(n_226),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_229),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_298),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_303),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_303),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_305),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

AND2x6_ASAP7_75t_L g434 ( 
.A(n_299),
.B(n_230),
.Y(n_434)
);

BUFx4f_ASAP7_75t_L g435 ( 
.A(n_299),
.Y(n_435)
);

AND3x2_ASAP7_75t_L g436 ( 
.A(n_333),
.B(n_235),
.C(n_233),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_280),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_333),
.A2(n_243),
.B1(n_227),
.B2(n_247),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_295),
.A2(n_243),
.B1(n_247),
.B2(n_250),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_336),
.A2(n_282),
.B1(n_281),
.B2(n_236),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_335),
.A2(n_244),
.B1(n_276),
.B2(n_273),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_314),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_309),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_296),
.B(n_262),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_309),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_341),
.B(n_237),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_314),
.Y(n_451)
);

NAND3xp33_ASAP7_75t_L g452 ( 
.A(n_332),
.B(n_240),
.C(n_272),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_297),
.B(n_239),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_329),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_335),
.B(n_246),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_315),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_342),
.B(n_249),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_307),
.B(n_179),
.Y(n_458)
);

INVxp33_ASAP7_75t_SL g459 ( 
.A(n_361),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_346),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_325),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_322),
.B(n_270),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_357),
.A2(n_258),
.B1(n_260),
.B2(n_269),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_320),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_434),
.A2(n_332),
.B1(n_360),
.B2(n_270),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_357),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_359),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_411),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_369),
.B(n_377),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_367),
.B(n_356),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_411),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_366),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_328),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_362),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_388),
.B(n_348),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_350),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_414),
.B(n_353),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_373),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_434),
.A2(n_337),
.B1(n_361),
.B2(n_343),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_390),
.B(n_268),
.Y(n_488)
);

OAI221xp5_ASAP7_75t_L g489 ( 
.A1(n_371),
.A2(n_300),
.B1(n_339),
.B2(n_343),
.C(n_213),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_387),
.A2(n_339),
.B(n_338),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_363),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_390),
.B(n_234),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_379),
.B(n_181),
.Y(n_494)
);

O2A1O1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_338),
.B(n_327),
.C(n_320),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_395),
.B(n_385),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_370),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_452),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_382),
.B(n_313),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_435),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_375),
.B(n_219),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_376),
.B(n_220),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_450),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_383),
.B(n_221),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_383),
.B(n_238),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_435),
.B(n_313),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_456),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_454),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_241),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_374),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_374),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_454),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_418),
.B(n_278),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_389),
.B(n_251),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_365),
.B(n_409),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_439),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_436),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_397),
.B(n_267),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_401),
.B(n_256),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_401),
.B(n_24),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_419),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_454),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_444),
.B(n_463),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_422),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_381),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_365),
.B(n_409),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_31),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_463),
.B(n_445),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_394),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_449),
.B(n_55),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_394),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_537)
);

NOR3xp33_ASAP7_75t_L g538 ( 
.A(n_405),
.B(n_40),
.C(n_41),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_447),
.B(n_41),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_430),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_457),
.B(n_43),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_408),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_410),
.B(n_58),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_436),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_386),
.B(n_63),
.C(n_68),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_69),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_446),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_420),
.B(n_70),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_417),
.B(n_72),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_461),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_405),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_472),
.A2(n_455),
.B(n_440),
.Y(n_553)
);

OAI22x1_ASAP7_75t_L g554 ( 
.A1(n_476),
.A2(n_462),
.B1(n_438),
.B2(n_403),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_486),
.A2(n_459),
.B1(n_407),
.B2(n_413),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_485),
.A2(n_455),
.B(n_440),
.Y(n_556)
);

AO22x1_ASAP7_75t_L g557 ( 
.A1(n_517),
.A2(n_459),
.B1(n_417),
.B2(n_403),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_525),
.A2(n_447),
.B1(n_407),
.B2(n_413),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_468),
.A2(n_421),
.B(n_427),
.C(n_431),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_474),
.B(n_511),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

CKINVDCx8_ASAP7_75t_R g562 ( 
.A(n_549),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_517),
.A2(n_407),
.B1(n_413),
.B2(n_421),
.Y(n_563)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_493),
.A2(n_427),
.B(n_431),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_474),
.B(n_432),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_497),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_488),
.A2(n_364),
.B(n_368),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_549),
.A2(n_499),
.B1(n_465),
.B2(n_520),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g569 ( 
.A1(n_491),
.A2(n_464),
.B(n_443),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_477),
.B(n_469),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_549),
.A2(n_443),
.B1(n_441),
.B2(n_453),
.Y(n_572)
);

BUFx4_ASAP7_75t_SL g573 ( 
.A(n_539),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

AOI22x1_ASAP7_75t_L g575 ( 
.A1(n_490),
.A2(n_393),
.B1(n_378),
.B2(n_406),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

CKINVDCx11_ASAP7_75t_R g577 ( 
.A(n_529),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_498),
.A2(n_460),
.B1(n_433),
.B2(n_404),
.Y(n_579)
);

AO32x1_ASAP7_75t_L g580 ( 
.A1(n_546),
.A2(n_404),
.A3(n_400),
.B1(n_399),
.B2(n_396),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_487),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_547),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_480),
.A2(n_392),
.B(n_380),
.C(n_396),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_484),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_511),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_496),
.A2(n_393),
.B(n_384),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_496),
.A2(n_384),
.B(n_372),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_500),
.B(n_460),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_518),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_544),
.B(n_83),
.Y(n_590)
);

OR2x6_ASAP7_75t_SL g591 ( 
.A(n_521),
.B(n_90),
.Y(n_591)
);

O2A1O1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_489),
.A2(n_522),
.B(n_531),
.C(n_532),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_SL g593 ( 
.A(n_538),
.B(n_95),
.C(n_101),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_466),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_467),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_512),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_R g597 ( 
.A(n_519),
.B(n_103),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_507),
.B(n_104),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_526),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_475),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_174),
.Y(n_601)
);

O2A1O1Ixp33_ASAP7_75t_SL g602 ( 
.A1(n_536),
.A2(n_123),
.B(n_124),
.C(n_125),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_495),
.A2(n_127),
.B(n_128),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_471),
.Y(n_605)
);

OA22x2_ASAP7_75t_L g606 ( 
.A1(n_535),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_505),
.B(n_138),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_505),
.B(n_140),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_527),
.B(n_141),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_542),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_157),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_506),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_528),
.B(n_540),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_470),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_478),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_526),
.Y(n_616)
);

O2A1O1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_541),
.A2(n_538),
.B(n_533),
.C(n_534),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_551),
.A2(n_158),
.B1(n_159),
.B2(n_164),
.Y(n_618)
);

AOI21x1_ASAP7_75t_L g619 ( 
.A1(n_543),
.A2(n_166),
.B(n_167),
.Y(n_619)
);

NOR2x1_ASAP7_75t_L g620 ( 
.A(n_545),
.B(n_170),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_523),
.A2(n_537),
.B1(n_552),
.B2(n_550),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_508),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_501),
.A2(n_502),
.B(n_515),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_523),
.A2(n_473),
.B1(n_510),
.B2(n_508),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_509),
.A2(n_524),
.B(n_513),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_616),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_558),
.B(n_514),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_562),
.A2(n_504),
.B1(n_482),
.B2(n_492),
.Y(n_628)
);

CKINVDCx11_ASAP7_75t_R g629 ( 
.A(n_591),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_558),
.A2(n_514),
.B1(n_530),
.B2(n_516),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_595),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_616),
.Y(n_632)
);

AO32x2_ASAP7_75t_L g633 ( 
.A1(n_621),
.A2(n_516),
.A3(n_530),
.B1(n_548),
.B2(n_503),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

BUFx2_ASAP7_75t_R g635 ( 
.A(n_589),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_584),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_570),
.B(n_479),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_603),
.B(n_526),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_576),
.B(n_563),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_557),
.B(n_555),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_582),
.B(n_612),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_616),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_568),
.B(n_572),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_556),
.A2(n_592),
.B(n_625),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_586),
.A2(n_587),
.B(n_624),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_613),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_577),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_566),
.B(n_594),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_605),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

OAI22x1_ASAP7_75t_L g651 ( 
.A1(n_598),
.A2(n_554),
.B1(n_574),
.B2(n_573),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_596),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_574),
.B(n_581),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_585),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_599),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_601),
.B(n_596),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_606),
.B(n_614),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_600),
.B(n_622),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_606),
.A2(n_593),
.B1(n_610),
.B2(n_604),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_564),
.A2(n_575),
.B(n_619),
.Y(n_660)
);

INVx5_ASAP7_75t_SL g661 ( 
.A(n_588),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_588),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_569),
.B(n_560),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_609),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_579),
.Y(n_665)
);

BUFx8_ASAP7_75t_L g666 ( 
.A(n_561),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_590),
.B(n_571),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_567),
.A2(n_565),
.B(n_580),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_611),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_608),
.A2(n_571),
.B1(n_597),
.B2(n_620),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_602),
.B(n_618),
.Y(n_671)
);

AO31x2_ASAP7_75t_L g672 ( 
.A1(n_580),
.A2(n_559),
.A3(n_621),
.B(n_583),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_616),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_558),
.A2(n_381),
.B1(n_408),
.B2(n_439),
.Y(n_674)
);

AO21x1_ASAP7_75t_L g675 ( 
.A1(n_604),
.A2(n_610),
.B(n_536),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_578),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_578),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_595),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_616),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_558),
.B(n_447),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_570),
.B(n_578),
.Y(n_681)
);

OAI22x1_ASAP7_75t_L g682 ( 
.A1(n_562),
.A2(n_462),
.B1(n_438),
.B2(n_476),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_576),
.Y(n_683)
);

AO31x2_ASAP7_75t_L g684 ( 
.A1(n_559),
.A2(n_621),
.A3(n_583),
.B(n_610),
.Y(n_684)
);

OA21x2_ASAP7_75t_L g685 ( 
.A1(n_604),
.A2(n_583),
.B(n_559),
.Y(n_685)
);

AO31x2_ASAP7_75t_L g686 ( 
.A1(n_559),
.A2(n_621),
.A3(n_583),
.B(n_610),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_578),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_616),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_558),
.B(n_447),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_595),
.Y(n_690)
);

AO31x2_ASAP7_75t_L g691 ( 
.A1(n_559),
.A2(n_621),
.A3(n_583),
.B(n_610),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_582),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_570),
.B(n_578),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_595),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_617),
.A2(n_592),
.B(n_623),
.C(n_468),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_604),
.B(n_332),
.C(n_394),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_559),
.A2(n_553),
.B(n_556),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_576),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_570),
.B(n_578),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_570),
.A2(n_595),
.B1(n_584),
.B2(n_578),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_681),
.B(n_693),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_699),
.B(n_634),
.Y(n_702)
);

AO31x2_ASAP7_75t_L g703 ( 
.A1(n_695),
.A2(n_645),
.A3(n_675),
.B(n_644),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_629),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_631),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_636),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_678),
.Y(n_707)
);

AO21x2_ASAP7_75t_L g708 ( 
.A1(n_659),
.A2(n_660),
.B(n_697),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_687),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_634),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_700),
.A2(n_674),
.B1(n_680),
.B2(n_689),
.Y(n_711)
);

NOR2x1_ASAP7_75t_SL g712 ( 
.A(n_676),
.B(n_677),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_676),
.B(n_677),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_646),
.B(n_637),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_646),
.B(n_627),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_639),
.B(n_692),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_649),
.B(n_648),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_683),
.B(n_698),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_641),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_656),
.B(n_626),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_654),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_666),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

OAI21x1_ASAP7_75t_SL g724 ( 
.A1(n_690),
.A2(n_694),
.B(n_630),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_652),
.B(n_656),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_643),
.A2(n_682),
.B1(n_653),
.B2(n_628),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_658),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_640),
.B(n_661),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_666),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_665),
.B(n_657),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_696),
.A2(n_669),
.B(n_664),
.C(n_671),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_655),
.Y(n_732)
);

OAI21x1_ASAP7_75t_SL g733 ( 
.A1(n_652),
.A2(n_664),
.B(n_670),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_632),
.Y(n_734)
);

AO22x1_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_651),
.B1(n_647),
.B2(n_688),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_661),
.B(n_638),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_672),
.Y(n_739)
);

NOR2x1_ASAP7_75t_SL g740 ( 
.A(n_679),
.B(n_673),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_679),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_679),
.B(n_688),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_642),
.B(n_673),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_642),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_684),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_633),
.A2(n_667),
.B(n_686),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_691),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_666),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_681),
.B(n_693),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_681),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_681),
.Y(n_752)
);

AO31x2_ASAP7_75t_L g753 ( 
.A1(n_695),
.A2(n_645),
.A3(n_675),
.B(n_644),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_681),
.B(n_699),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_659),
.B(n_643),
.Y(n_755)
);

AO21x2_ASAP7_75t_L g756 ( 
.A1(n_668),
.A2(n_659),
.B(n_645),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_681),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_695),
.A2(n_645),
.A3(n_675),
.B(n_644),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_652),
.B(n_595),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_666),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_745),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_759),
.Y(n_762)
);

INVx6_ASAP7_75t_L g763 ( 
.A(n_754),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_754),
.B(n_701),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_750),
.B(n_711),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_751),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_752),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_710),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_713),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_759),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_705),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_741),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_755),
.B(n_735),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_757),
.B(n_702),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_705),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_760),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_707),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_727),
.B(n_712),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_741),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_717),
.B(n_715),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_730),
.B(n_723),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_706),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_714),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_729),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_721),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_709),
.Y(n_787)
);

HB1xp67_ASAP7_75t_SL g788 ( 
.A(n_760),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_755),
.B(n_724),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_737),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_725),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_746),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_719),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_729),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_718),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_716),
.B(n_732),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_734),
.Y(n_797)
);

INVx4_ASAP7_75t_SL g798 ( 
.A(n_703),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_736),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_742),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_726),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_753),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_753),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_731),
.A2(n_738),
.B1(n_725),
.B2(n_749),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_764),
.B(n_747),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_792),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_792),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_764),
.B(n_747),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_801),
.B(n_748),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_771),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_801),
.B(n_739),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_793),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_798),
.B(n_756),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_765),
.A2(n_728),
.B1(n_733),
.B2(n_749),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_761),
.Y(n_815)
);

CKINVDCx10_ASAP7_75t_R g816 ( 
.A(n_773),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_765),
.B(n_758),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_763),
.A2(n_722),
.B1(n_720),
.B2(n_744),
.Y(n_818)
);

INVx5_ASAP7_75t_L g819 ( 
.A(n_770),
.Y(n_819)
);

INVx5_ASAP7_75t_SL g820 ( 
.A(n_773),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_775),
.B(n_777),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_766),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_769),
.B(n_753),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_775),
.B(n_777),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_781),
.B(n_708),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_778),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_778),
.Y(n_827)
);

NOR2x1p5_ASAP7_75t_L g828 ( 
.A(n_770),
.B(n_722),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_806),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_819),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_810),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_812),
.B(n_794),
.C(n_795),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_805),
.B(n_802),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_806),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_807),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_813),
.B(n_798),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_807),
.Y(n_837)
);

AOI221xp5_ASAP7_75t_L g838 ( 
.A1(n_822),
.A2(n_784),
.B1(n_767),
.B2(n_790),
.C(n_781),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_805),
.B(n_803),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_819),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_826),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_821),
.B(n_790),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_815),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_821),
.B(n_783),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_824),
.B(n_783),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_808),
.B(n_803),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_808),
.B(n_798),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_840),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_833),
.B(n_839),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_829),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_833),
.B(n_809),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_839),
.B(n_809),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_843),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_846),
.B(n_825),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_834),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_835),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_846),
.B(n_823),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_835),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_847),
.B(n_811),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_847),
.B(n_811),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_837),
.B(n_823),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_842),
.B(n_826),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_844),
.B(n_827),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_837),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_849),
.B(n_841),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_849),
.B(n_854),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_861),
.B(n_845),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_862),
.A2(n_773),
.B1(n_763),
.B2(n_838),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_861),
.B(n_825),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_850),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_851),
.B(n_817),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_850),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_853),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_863),
.B(n_830),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_859),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_851),
.B(n_798),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_852),
.B(n_813),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_868),
.A2(n_773),
.B1(n_832),
.B2(n_785),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_866),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_871),
.B(n_852),
.Y(n_880)
);

OAI221xp5_ASAP7_75t_L g881 ( 
.A1(n_868),
.A2(n_814),
.B1(n_773),
.B2(n_804),
.C(n_786),
.Y(n_881)
);

NOR3xp33_ASAP7_75t_L g882 ( 
.A(n_865),
.B(n_797),
.C(n_776),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_876),
.A2(n_857),
.B1(n_860),
.B2(n_859),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_876),
.A2(n_874),
.B1(n_875),
.B2(n_877),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_873),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_869),
.B(n_854),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_870),
.Y(n_887)
);

OAI22xp33_ASAP7_75t_L g888 ( 
.A1(n_874),
.A2(n_830),
.B1(n_819),
.B2(n_831),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_867),
.B(n_872),
.Y(n_889)
);

AOI211xp5_ASAP7_75t_SL g890 ( 
.A1(n_881),
.A2(n_830),
.B(n_704),
.C(n_817),
.Y(n_890)
);

XNOR2xp5_ASAP7_75t_L g891 ( 
.A(n_882),
.B(n_704),
.Y(n_891)
);

NOR4xp25_ASAP7_75t_L g892 ( 
.A(n_879),
.B(n_787),
.C(n_796),
.D(n_799),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_884),
.B(n_819),
.Y(n_893)
);

AOI222xp33_ASAP7_75t_L g894 ( 
.A1(n_889),
.A2(n_877),
.B1(n_831),
.B2(n_796),
.C1(n_860),
.C2(n_864),
.Y(n_894)
);

OAI222xp33_ASAP7_75t_L g895 ( 
.A1(n_878),
.A2(n_874),
.B1(n_848),
.B2(n_788),
.C1(n_819),
.C2(n_810),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_894),
.A2(n_883),
.B1(n_874),
.B2(n_886),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_893),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_890),
.A2(n_828),
.B(n_885),
.C(n_880),
.Y(n_898)
);

OA21x2_ASAP7_75t_SL g899 ( 
.A1(n_896),
.A2(n_892),
.B(n_891),
.Y(n_899)
);

NAND4xp25_ASAP7_75t_SL g900 ( 
.A(n_898),
.B(n_895),
.C(n_893),
.D(n_816),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_900),
.B(n_828),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_899),
.B(n_897),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_901),
.B(n_887),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_902),
.A2(n_888),
.B(n_774),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_903),
.Y(n_905)
);

XNOR2x1_ASAP7_75t_L g906 ( 
.A(n_904),
.B(n_779),
.Y(n_906)
);

OA22x2_ASAP7_75t_L g907 ( 
.A1(n_905),
.A2(n_787),
.B1(n_799),
.B2(n_816),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_906),
.Y(n_908)
);

XNOR2xp5_ASAP7_75t_L g909 ( 
.A(n_905),
.B(n_818),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_SL g910 ( 
.A1(n_908),
.A2(n_819),
.B1(n_770),
.B2(n_791),
.Y(n_910)
);

OAI22x1_ASAP7_75t_L g911 ( 
.A1(n_909),
.A2(n_819),
.B1(n_720),
.B2(n_770),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_907),
.Y(n_912)
);

AOI221xp5_ASAP7_75t_L g913 ( 
.A1(n_908),
.A2(n_768),
.B1(n_779),
.B2(n_782),
.C(n_780),
.Y(n_913)
);

AOI222xp33_ASAP7_75t_L g914 ( 
.A1(n_910),
.A2(n_768),
.B1(n_820),
.B2(n_782),
.C1(n_780),
.C2(n_772),
.Y(n_914)
);

OAI222xp33_ASAP7_75t_L g915 ( 
.A1(n_912),
.A2(n_762),
.B1(n_772),
.B2(n_780),
.C1(n_789),
.C2(n_791),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_911),
.A2(n_740),
.B(n_743),
.Y(n_916)
);

AO22x2_ASAP7_75t_SL g917 ( 
.A1(n_913),
.A2(n_780),
.B1(n_772),
.B2(n_800),
.Y(n_917)
);

XNOR2xp5_ASAP7_75t_L g918 ( 
.A(n_917),
.B(n_791),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_SL g919 ( 
.A1(n_915),
.A2(n_742),
.B(n_836),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_SL g920 ( 
.A(n_918),
.B(n_916),
.C(n_914),
.Y(n_920)
);

AOI222xp33_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_919),
.B1(n_820),
.B2(n_858),
.C1(n_856),
.C2(n_855),
.Y(n_921)
);


endmodule