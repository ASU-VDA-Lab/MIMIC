module fake_netlist_1_1510_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NOR2xp33_ASAP7_75t_L g5 ( .A(n_2), .B(n_0), .Y(n_5) );
A2O1A1Ixp33_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
NOR2xp67_ASAP7_75t_SL g7 ( .A(n_3), .B(n_0), .Y(n_7) );
NOR2xp33_ASAP7_75t_R g8 ( .A(n_4), .B(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .Y(n_11) );
NOR2xp33_ASAP7_75t_SL g12 ( .A(n_9), .B(n_6), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_9), .Y(n_13) );
AOI32xp33_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_1), .A3(n_2), .B1(n_5), .B2(n_11), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
NAND4xp75_ASAP7_75t_L g16 ( .A(n_14), .B(n_12), .C(n_2), .D(n_1), .Y(n_16) );
AO21x2_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_1), .B(n_16), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_10), .Y(n_18) );
endmodule