module fake_jpeg_10934_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_46),
.B(n_49),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_57),
.Y(n_131)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_59),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_67),
.Y(n_150)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_72),
.Y(n_102)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_7),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_78),
.B(n_31),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_9),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_44),
.B(n_34),
.C(n_35),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_93),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_64),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_105),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_31),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_111),
.B(n_93),
.Y(n_199)
);

BUFx2_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_53),
.B(n_24),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_128),
.Y(n_161)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_43),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_149),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_45),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_52),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_147),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_47),
.B(n_37),
.C(n_40),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_91),
.Y(n_149)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_56),
.B1(n_70),
.B2(n_85),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_154),
.A2(n_164),
.B1(n_178),
.B2(n_100),
.Y(n_206)
);

CKINVDCx12_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_106),
.B(n_40),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_160),
.B(n_168),
.Y(n_207)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_145),
.A2(n_65),
.B1(n_88),
.B2(n_84),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_185),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_66),
.B1(n_83),
.B2(n_81),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_195),
.B1(n_77),
.B2(n_75),
.Y(n_205)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_105),
.A2(n_100),
.B1(n_16),
.B2(n_24),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_173),
.A2(n_175),
.B1(n_192),
.B2(n_196),
.Y(n_235)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_111),
.B1(n_123),
.B2(n_95),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_197),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_48),
.B1(n_69),
.B2(n_61),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_37),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_131),
.A2(n_150),
.B1(n_102),
.B2(n_104),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_38),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

AO22x2_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_86),
.B1(n_50),
.B2(n_62),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_35),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_11),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_193),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_194),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_97),
.A2(n_73),
.B1(n_71),
.B2(n_80),
.Y(n_195)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_200),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_134),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_109),
.C(n_134),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_210),
.B(n_157),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_182),
.B1(n_179),
.B2(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_118),
.B1(n_151),
.B2(n_136),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_217),
.B(n_158),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_168),
.A2(n_139),
.B(n_127),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_232),
.B(n_127),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_124),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_124),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_166),
.A2(n_144),
.B1(n_116),
.B2(n_137),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_233),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_144),
.B1(n_116),
.B2(n_136),
.Y(n_229)
);

AO21x1_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_182),
.B(n_175),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_174),
.B(n_175),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_112),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_267),
.B(n_183),
.Y(n_279)
);

CKINVDCx12_ASAP7_75t_R g239 ( 
.A(n_201),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_240),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_241),
.B(n_246),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_188),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_242),
.B(n_243),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_169),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_248),
.Y(n_272)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_184),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_253),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_254),
.B1(n_181),
.B2(n_192),
.Y(n_287)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_151),
.B1(n_118),
.B2(n_197),
.Y(n_254)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_256),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_257),
.B(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_153),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_266),
.B(n_211),
.Y(n_280)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_213),
.B1(n_115),
.B2(n_234),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_156),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_183),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_210),
.B(n_211),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_217),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_208),
.B(n_156),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_265),
.C(n_237),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_235),
.B(n_209),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_270),
.A2(n_241),
.B(n_266),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_215),
.B1(n_206),
.B2(n_224),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_285),
.B1(n_295),
.B2(n_299),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_278),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_292),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_205),
.B1(n_227),
.B2(n_196),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_263),
.B1(n_240),
.B2(n_245),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_292),
.B(n_252),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_234),
.B(n_213),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_262),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_297),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_251),
.A2(n_220),
.B1(n_170),
.B2(n_187),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_239),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_220),
.B1(n_190),
.B2(n_193),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_300),
.A2(n_326),
.B(n_274),
.Y(n_348)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_243),
.Y(n_302)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_287),
.B1(n_278),
.B2(n_282),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_304),
.A2(n_311),
.B1(n_316),
.B2(n_323),
.Y(n_354)
);

OR2x4_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_264),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_305),
.A2(n_317),
.B(n_321),
.C(n_252),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_255),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_307),
.B(n_308),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_244),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_269),
.C(n_297),
.Y(n_334)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_278),
.A2(n_282),
.B1(n_238),
.B2(n_291),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_272),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_315),
.Y(n_333)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_314),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_291),
.A2(n_247),
.B1(n_237),
.B2(n_293),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_276),
.B(n_293),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_274),
.B(n_281),
.Y(n_339)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_248),
.Y(n_328)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_328),
.Y(n_344)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_329),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_254),
.Y(n_330)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_254),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_271),
.B(n_242),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_271),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_337),
.C(n_353),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_320),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_343),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_324),
.A2(n_264),
.B1(n_250),
.B2(n_273),
.Y(n_336)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_336),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_295),
.Y(n_337)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_339),
.A2(n_348),
.B(n_362),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_317),
.A2(n_285),
.B1(n_250),
.B2(n_253),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_340),
.A2(n_357),
.B1(n_304),
.B2(n_300),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_320),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_311),
.B(n_277),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_328),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_310),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_299),
.B(n_256),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_349),
.B(n_351),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_268),
.C(n_225),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_317),
.A2(n_273),
.B1(n_284),
.B2(n_268),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_306),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_360),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_302),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_326),
.A2(n_284),
.B(n_256),
.Y(n_362)
);

O2A1O1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_301),
.B(n_319),
.C(n_318),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_167),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_326),
.C(n_327),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_373),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_367),
.B(n_162),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_368),
.A2(n_386),
.B1(n_389),
.B2(n_392),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_333),
.Y(n_369)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_324),
.B1(n_332),
.B2(n_322),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_322),
.B1(n_331),
.B2(n_330),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_374),
.A2(n_379),
.B1(n_380),
.B2(n_388),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_376),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_305),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_212),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_255),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_342),
.B(n_303),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_394),
.B(n_372),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_342),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_387),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_355),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_314),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_325),
.B1(n_323),
.B2(n_300),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_390),
.A2(n_393),
.B1(n_339),
.B2(n_350),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_SL g409 ( 
.A1(n_391),
.A2(n_357),
.B(n_356),
.C(n_363),
.Y(n_409)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_356),
.B1(n_350),
.B2(n_359),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_371),
.A2(n_365),
.B1(n_370),
.B2(n_388),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_414),
.A3(n_228),
.B1(n_230),
.B2(n_219),
.C1(n_172),
.C2(n_33),
.Y(n_432)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_404),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_345),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_353),
.C(n_364),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_412),
.C(n_413),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_372),
.A2(n_355),
.B(n_363),
.Y(n_407)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_348),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_411),
.Y(n_424)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_363),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_359),
.C(n_318),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_329),
.C(n_303),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_390),
.A2(n_284),
.B1(n_240),
.B2(n_245),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_366),
.B(n_394),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_416),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_301),
.C(n_236),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_381),
.C(n_392),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_419),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_236),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_109),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_397),
.Y(n_421)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_391),
.B1(n_389),
.B2(n_386),
.Y(n_422)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_393),
.B(n_204),
.Y(n_425)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_204),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

BUFx12f_ASAP7_75t_SL g429 ( 
.A(n_406),
.Y(n_429)
);

AOI21xp33_ASAP7_75t_L g458 ( 
.A1(n_429),
.A2(n_430),
.B(n_405),
.Y(n_458)
);

OA21x2_ASAP7_75t_SL g430 ( 
.A1(n_404),
.A2(n_216),
.B(n_219),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_432),
.A2(n_24),
.B1(n_16),
.B2(n_89),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_216),
.B(n_159),
.Y(n_434)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_230),
.B1(n_39),
.B2(n_33),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_435),
.A2(n_440),
.B1(n_39),
.B2(n_32),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g437 ( 
.A(n_409),
.B(n_115),
.CI(n_2),
.CON(n_437),
.SN(n_437)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_438),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_418),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_420),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_410),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_440)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_412),
.C(n_408),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_452),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_401),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_451),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_413),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_419),
.C(n_416),
.Y(n_452)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_409),
.C(n_417),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_456),
.A2(n_457),
.B(n_458),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_409),
.C(n_405),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_462),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_32),
.C(n_91),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_460),
.B(n_434),
.C(n_425),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_435),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_427),
.A2(n_16),
.B1(n_79),
.B2(n_3),
.Y(n_462)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_457),
.B(n_424),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_454),
.A2(n_441),
.B1(n_431),
.B2(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_470),
.B(n_476),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_443),
.C(n_426),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_472),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_421),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_447),
.A2(n_431),
.B(n_422),
.Y(n_475)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_475),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_439),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_437),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_477),
.B(n_478),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_445),
.B(n_437),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_444),
.B(n_456),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_480),
.A2(n_6),
.B(n_9),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_452),
.Y(n_486)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_486),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_475),
.Y(n_487)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_487),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g489 ( 
.A1(n_468),
.A2(n_449),
.B(n_455),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_491),
.B(n_5),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_460),
.C(n_42),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_5),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_10),
.B(n_2),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_465),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_494),
.Y(n_504)
);

AOI322xp5_ASAP7_75t_L g494 ( 
.A1(n_488),
.A2(n_475),
.A3(n_474),
.B1(n_463),
.B2(n_473),
.C1(n_10),
.C2(n_11),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_496),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_498),
.C(n_499),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_479),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_6),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_42),
.C(n_6),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_483),
.C(n_489),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_506),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_493),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_500),
.A2(n_484),
.B(n_481),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_12),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_494),
.A3(n_501),
.B1(n_12),
.B2(n_13),
.C1(n_9),
.C2(n_0),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_510),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_12),
.C(n_13),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_505),
.C(n_509),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_508),
.B(n_13),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_514),
.B(n_513),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_0),
.C(n_493),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_0),
.Y(n_517)
);


endmodule