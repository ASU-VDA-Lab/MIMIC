module real_jpeg_30273_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g140 ( 
.A(n_0),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_0),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g479 ( 
.A(n_0),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_1),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_1),
.B(n_50),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_1),
.B(n_107),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_1),
.B(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_1),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_1),
.B(n_342),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_3),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_3),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_272),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_3),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_3),
.B(n_292),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_3),
.B(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_3),
.B(n_342),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_13),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_5),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g352 ( 
.A(n_5),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_5),
.B(n_55),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_5),
.B(n_433),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_6),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_7),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_9),
.Y(n_482)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_10),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_233),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g276 ( 
.A(n_11),
.B(n_137),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_11),
.B(n_304),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_11),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_11),
.B(n_445),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g480 ( 
.A(n_11),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_11),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_12),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_12),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_12),
.B(n_50),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_12),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_12),
.B(n_166),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_12),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_12),
.B(n_502),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2x1_ASAP7_75t_SL g62 ( 
.A(n_14),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_14),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_139),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_15),
.Y(n_122)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_15),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

NAND2x1_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_16),
.B(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_18),
.B(n_185),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g218 ( 
.A(n_18),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_18),
.B(n_248),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_18),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_18),
.B(n_407),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_18),
.B(n_450),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_18),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_18),
.B(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_19),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_19),
.B(n_180),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_19),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_19),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_192),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_R g23 ( 
.A(n_24),
.B(n_190),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_146),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_25),
.B(n_146),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_111),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_72),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.C(n_57),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_28),
.B(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_30),
.A2(n_38),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_30),
.B(n_39),
.C(n_40),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_32),
.Y(n_167)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_32),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_33),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_129)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_37),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_48),
.C(n_53),
.Y(n_47)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_46),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_46),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_46),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_47),
.B(n_57),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_48),
.B(n_129),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_52),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_53),
.A2(n_54),
.B1(n_138),
.B2(n_183),
.Y(n_188)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_136),
.C(n_138),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_56),
.Y(n_430)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_56),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_66),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_66),
.B1(n_67),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_71),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_98),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_83),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_93),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_92),
.Y(n_304)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_96),
.Y(n_411)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_97),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_109),
.B2(n_110),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_130),
.B(n_145),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_128),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_116),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_123),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_120),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_122),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_125),
.B(n_279),
.Y(n_426)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g488 ( 
.A(n_127),
.Y(n_488)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_134),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.C(n_144),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_179),
.B1(n_183),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_144),
.Y(n_158)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_160),
.C(n_168),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_144),
.B(n_169),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_153),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_151),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_159),
.C(n_174),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_159),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_162),
.Y(n_229)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_187),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_176),
.B(n_178),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_182),
.Y(n_339)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_187),
.B(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_526),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_255),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_SL g527 ( 
.A(n_197),
.B(n_199),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_R g199 ( 
.A(n_200),
.B(n_203),
.C(n_206),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_203),
.Y(n_316)
);

XNOR2x2_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_207),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_230),
.C(n_252),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.C(n_228),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_213),
.C(n_228),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_213),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_226),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_218),
.B(n_227),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_221),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_253),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_241),
.B(n_251),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_309)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_247),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_247),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_242),
.B(n_247),
.Y(n_310)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_246),
.Y(n_355)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_246),
.Y(n_451)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_365),
.B(n_523),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_317),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_257),
.A2(n_524),
.B(n_525),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_314),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_258),
.B(n_314),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.C(n_312),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_260),
.B(n_312),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_263),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_287),
.C(n_305),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_321),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.C(n_281),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_266),
.B(n_268),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_269),
.A2(n_270),
.B1(n_281),
.B2(n_282),
.Y(n_392)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B(n_277),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_271),
.B(n_332),
.Y(n_331)
);

AOI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_278),
.B(n_280),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_274),
.A2(n_275),
.B1(n_280),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OA21x2_ASAP7_75t_SL g376 ( 
.A1(n_282),
.A2(n_283),
.B(n_286),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_306),
.B1(n_307),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_298),
.C(n_302),
.Y(n_288)
);

XOR2x1_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_362),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_293),
.Y(n_447)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_363),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_318),
.B(n_363),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_328),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_320),
.B(n_324),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_356),
.C(n_359),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_329),
.A2(n_330),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.C(n_345),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_334),
.A2(n_345),
.B1(n_346),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_340),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_335),
.A2(n_336),
.B1(n_340),
.B2(n_341),
.Y(n_412)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_344),
.Y(n_504)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.C(n_352),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_347),
.A2(n_348),
.B1(n_352),
.B2(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_351),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_360),
.B1(n_361),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_419),
.B(n_521),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_393),
.B(n_396),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_367),
.B(n_393),
.C(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.C(n_389),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.C(n_377),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_376),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_377),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_383),
.C(n_385),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_435),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_379),
.A2(n_380),
.B1(n_381),
.B2(n_382),
.Y(n_425)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_435)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_417),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_397),
.B(n_417),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.C(n_413),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_414),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.C(n_412),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_412),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.C(n_409),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_405),
.B(n_409),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_438),
.B(n_520),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_436),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g520 ( 
.A(n_421),
.B(n_436),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.C(n_434),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_422),
.B(n_518),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_424),
.B(n_434),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.C(n_427),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_426),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

AO22x1_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_460)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_515),
.B(n_519),
.Y(n_438)
);

OAI21x1_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_472),
.B(n_514),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_461),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_461),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_454),
.C(n_460),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_442),
.A2(n_443),
.B1(n_510),
.B2(n_512),
.Y(n_509)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_448),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_467),
.C(n_468),
.Y(n_466)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_454),
.A2(n_455),
.B1(n_460),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_459),
.Y(n_490)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_460),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_465),
.B2(n_471),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_462),
.B(n_466),
.C(n_469),
.Y(n_516)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_465),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_507),
.B(n_513),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_491),
.B(n_506),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_483),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_475),
.B(n_483),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_480),
.Y(n_499)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx8_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_480),
.B(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_490),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_489),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_485),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_489),
.C(n_490),
.Y(n_508)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_500),
.B(n_505),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_499),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_499),
.Y(n_505)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_SL g502 ( 
.A(n_503),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_509),
.Y(n_513)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_510),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);


endmodule