module fake_jpeg_19777_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_36),
.B1(n_30),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_50),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_24),
.B1(n_36),
.B2(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_38),
.B1(n_44),
.B2(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_60),
.B(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_33),
.B1(n_28),
.B2(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_91),
.B1(n_96),
.B2(n_67),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_41),
.B1(n_48),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_82),
.B1(n_97),
.B2(n_26),
.Y(n_123)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_40),
.B1(n_33),
.B2(n_28),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_98),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_58),
.B1(n_53),
.B2(n_25),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_18),
.B1(n_22),
.B2(n_35),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_51),
.A2(n_40),
.B(n_26),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_46),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_26),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_22),
.B1(n_35),
.B2(n_17),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_37),
.B1(n_17),
.B2(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_23),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_102),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_52),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_105),
.B(n_95),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_65),
.C(n_56),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_114),
.C(n_126),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_50),
.B1(n_58),
.B2(n_32),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_112),
.B1(n_123),
.B2(n_85),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_69),
.B1(n_88),
.B2(n_74),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_26),
.B1(n_13),
.B2(n_11),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_31),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_14),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_111),
.B1(n_131),
.B2(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_143),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_146),
.B(n_105),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_145),
.C(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_75),
.B1(n_81),
.B2(n_79),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_117),
.B1(n_127),
.B2(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_122),
.C(n_103),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_88),
.C(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_113),
.A2(n_131),
.B1(n_71),
.B2(n_121),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_132),
.B1(n_87),
.B2(n_77),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_68),
.B1(n_86),
.B2(n_90),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_104),
.B1(n_68),
.B2(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_104),
.B(n_103),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_163),
.A2(n_172),
.B(n_176),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_171),
.B(n_191),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_166),
.B1(n_147),
.B2(n_139),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_152),
.B1(n_156),
.B2(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_124),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_168),
.B(n_175),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_144),
.B(n_138),
.C(n_141),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_180),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_124),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_119),
.B(n_121),
.Y(n_176)
);

AO22x1_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_87),
.B1(n_119),
.B2(n_71),
.Y(n_180)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_133),
.B1(n_107),
.B2(n_129),
.Y(n_181)
);

AOI22x1_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_147),
.B1(n_115),
.B2(n_21),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_107),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_128),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_129),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_152),
.B1(n_148),
.B2(n_158),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_21),
.B1(n_29),
.B2(n_34),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_34),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_190),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_220),
.B1(n_223),
.B2(n_2),
.Y(n_238)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_197),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_173),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_199),
.B(n_202),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_180),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_159),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_159),
.C(n_139),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_216),
.C(n_164),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_21),
.C(n_29),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_166),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_212),
.A2(n_187),
.B1(n_172),
.B2(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_174),
.C(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_177),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_181),
.B(n_190),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_115),
.B1(n_29),
.B2(n_34),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_172),
.A2(n_115),
.B1(n_29),
.B2(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_167),
.B(n_15),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_198),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_233),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_245),
.C(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_248),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_171),
.B(n_180),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_191),
.B(n_189),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_194),
.A2(n_0),
.B(n_1),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_235),
.B(n_3),
.Y(n_264)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_200),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_8),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_247),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_212),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_2),
.B(n_3),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_8),
.C(n_12),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_9),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_9),
.B(n_12),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_252),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_196),
.B1(n_207),
.B2(n_194),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_265),
.B1(n_269),
.B2(n_197),
.Y(n_288)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVx2_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_270),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_208),
.C(n_196),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_229),
.C(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g270 ( 
.A(n_233),
.B(n_201),
.C(n_223),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_273),
.C(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_225),
.C(n_245),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_201),
.CI(n_247),
.CON(n_274),
.SN(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_230),
.C(n_228),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_234),
.B(n_248),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_227),
.B(n_218),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_260),
.C(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_279),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_243),
.B(n_244),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_230),
.C(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_195),
.C(n_237),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_257),
.C(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

XOR2x2_ASAP7_75t_SL g289 ( 
.A(n_266),
.B(n_210),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_235),
.C(n_218),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_257),
.B1(n_236),
.B2(n_268),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_294),
.B1(n_296),
.B2(n_304),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_258),
.B1(n_254),
.B2(n_220),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_221),
.B1(n_209),
.B2(n_250),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_238),
.B1(n_221),
.B2(n_271),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_305),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_262),
.B1(n_249),
.B2(n_5),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_276),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_272),
.C(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_286),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_277),
.C(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_285),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_281),
.C(n_274),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_295),
.A2(n_286),
.B(n_10),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_296),
.B(n_294),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_293),
.C(n_303),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_291),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_311),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_319),
.A2(n_316),
.B(n_317),
.C(n_301),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_331),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_322),
.A2(n_321),
.B(n_313),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_307),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_318),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_318),
.C(n_309),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_329),
.B(n_298),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_328),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_337),
.B(n_330),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_302),
.A3(n_326),
.B1(n_7),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_10),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_14),
.C(n_5),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_14),
.B(n_5),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_344),
.B(n_6),
.CI(n_337),
.CON(n_345),
.SN(n_345)
);


endmodule