module fake_jpeg_10168_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_2),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_56),
.B1(n_66),
.B2(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_33),
.B1(n_30),
.B2(n_24),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_63),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_0),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_16),
.B1(n_30),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_16),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_40),
.B1(n_44),
.B2(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_74),
.B1(n_81),
.B2(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_72),
.B1(n_78),
.B2(n_55),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_23),
.B(n_29),
.C(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_66),
.Y(n_98)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_27),
.B1(n_28),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_50),
.B1(n_45),
.B2(n_55),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_23),
.B1(n_31),
.B2(n_38),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_38),
.C(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_39),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_62),
.B(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_91),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_75),
.C(n_48),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_101),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_65),
.B1(n_38),
.B2(n_39),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_89),
.B1(n_52),
.B2(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_53),
.B1(n_55),
.B2(n_29),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_109),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_106),
.B1(n_112),
.B2(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_56),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_120),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_95),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_87),
.B1(n_69),
.B2(n_86),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_85),
.B1(n_68),
.B2(n_86),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_135),
.B1(n_98),
.B2(n_95),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_86),
.B(n_48),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_1),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_1),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_1),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_101),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_138),
.B1(n_60),
.B2(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_72),
.B1(n_78),
.B2(n_75),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_60),
.C(n_76),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_99),
.B1(n_112),
.B2(n_106),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_146),
.B1(n_155),
.B2(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_149),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_118),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_144),
.C(n_162),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_97),
.B(n_99),
.C(n_104),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_125),
.B(n_64),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_97),
.B1(n_105),
.B2(n_110),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_133),
.B1(n_125),
.B2(n_60),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_150),
.Y(n_180)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_9),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_78),
.B1(n_93),
.B2(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_156),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_100),
.B1(n_90),
.B2(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_79),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_137),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_137),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_176),
.C(n_181),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_133),
.B1(n_120),
.B2(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_177),
.A2(n_153),
.B1(n_145),
.B2(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_119),
.C(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_179),
.B1(n_152),
.B2(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_143),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_131),
.C(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_196),
.C(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_203),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_151),
.CI(n_3),
.CON(n_202),
.SN(n_202)
);

XOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_202),
.B(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_145),
.Y(n_205)
);

OAI31xp33_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_207),
.A3(n_168),
.B(n_180),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_141),
.B1(n_180),
.B2(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_2),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_221),
.C(n_222),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_220),
.B1(n_108),
.B2(n_76),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_165),
.B(n_172),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_176),
.B1(n_202),
.B2(n_197),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_184),
.C(n_141),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_201),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_196),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_201),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_190),
.B1(n_202),
.B2(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_191),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_207),
.B1(n_206),
.B2(n_189),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_236),
.B1(n_224),
.B2(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_189),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_235),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_214),
.Y(n_246)
);

XOR2x1_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_212),
.Y(n_247)
);

AOI21x1_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_233),
.B(n_208),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_232),
.C(n_230),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_216),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_239),
.B(n_243),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_253),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_228),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_208),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_261),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_243),
.B(n_215),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_258),
.B(n_7),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_251),
.B(n_252),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_7),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

OAI211xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_8),
.B(n_11),
.C(n_13),
.Y(n_267)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_8),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_270),
.A3(n_14),
.B1(n_266),
.B2(n_88),
.C(n_77),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_77),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_14),
.B(n_77),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_88),
.Y(n_273)
);


endmodule