module fake_netlist_1_11709_n_993 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_993);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_993;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_185;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_973;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_961;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_948;
wire n_898;
wire n_126;
wire n_989;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_962;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_947;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_967;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_43), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_41), .Y(n_113) );
CKINVDCx11_ASAP7_75t_R g114 ( .A(n_40), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_95), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_67), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_103), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_21), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_81), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_18), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_55), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_110), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_72), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_50), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_3), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_12), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_37), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_90), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_84), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_13), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_80), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_5), .Y(n_133) );
OR2x2_ASAP7_75t_L g134 ( .A(n_47), .B(n_12), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_15), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_79), .B(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_75), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_65), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_39), .Y(n_139) );
CKINVDCx14_ASAP7_75t_R g140 ( .A(n_107), .Y(n_140) );
OR2x2_ASAP7_75t_L g141 ( .A(n_22), .B(n_85), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_17), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_5), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_20), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_25), .Y(n_146) );
INVx1_ASAP7_75t_SL g147 ( .A(n_42), .Y(n_147) );
INVxp67_ASAP7_75t_SL g148 ( .A(n_104), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_21), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_49), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_31), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_7), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_138), .Y(n_153) );
AOI22x1_ASAP7_75t_SL g154 ( .A1(n_126), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_138), .Y(n_155) );
BUFx8_ASAP7_75t_SL g156 ( .A(n_133), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_114), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_131), .B(n_0), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
NOR2x1_ASAP7_75t_L g162 ( .A(n_136), .B(n_1), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_118), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g172 ( .A(n_113), .B(n_23), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_143), .A2(n_2), .B1(n_4), .B2(n_6), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_175), .B(n_120), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_165), .B(n_120), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_175), .B(n_113), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_165), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_177), .B(n_117), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_167), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_171), .B(n_177), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_167), .B(n_117), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_178), .B(n_119), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_178), .B(n_119), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_167), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_167), .B(n_121), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_167), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_163), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_176), .B(n_121), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_176), .B(n_132), .Y(n_208) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_168), .A2(n_132), .B(n_151), .Y(n_209) );
BUFx10_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
NOR2x1p5_ASAP7_75t_L g211 ( .A(n_157), .B(n_174), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_160), .B(n_151), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_168), .B(n_127), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_159), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
INVxp33_ASAP7_75t_SL g221 ( .A(n_172), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
BUFx10_ASAP7_75t_L g223 ( .A(n_160), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_160), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
INVxp33_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
BUFx10_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_154), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_169), .B(n_135), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_169), .B(n_112), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_173), .B(n_149), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_159), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_161), .B(n_152), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_173), .B(n_125), .Y(n_237) );
XNOR2xp5_ASAP7_75t_L g238 ( .A(n_154), .B(n_145), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_164), .B(n_128), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_200), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_210), .B(n_129), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_196), .B(n_164), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_200), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_210), .B(n_166), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_188), .B(n_166), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_210), .B(n_170), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_224), .A2(n_170), .B(n_162), .C(n_147), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_226), .B(n_162), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_210), .B(n_116), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_183), .B(n_130), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_200), .Y(n_251) );
NOR3xp33_ASAP7_75t_L g252 ( .A(n_228), .B(n_179), .C(n_150), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_223), .B(n_24), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_209), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_208), .B(n_8), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_196), .B(n_8), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_198), .B(n_26), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_214), .B(n_9), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_214), .B(n_9), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_234), .A2(n_197), .B1(n_214), .B2(n_209), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_214), .B(n_27), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_209), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_232), .B(n_10), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_182), .B(n_11), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_234), .B(n_14), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_182), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_207), .B(n_63), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_218), .Y(n_270) );
NOR2xp33_ASAP7_75t_SL g271 ( .A(n_221), .B(n_14), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_223), .B(n_64), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_223), .B(n_66), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_216), .B(n_15), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_231), .B(n_16), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_190), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_190), .B(n_212), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_181), .B(n_16), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_239), .B(n_236), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_224), .B(n_17), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_185), .B(n_211), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_223), .B(n_69), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_224), .B(n_18), .Y(n_284) );
INVx5_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_237), .B(n_19), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_227), .B(n_70), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_227), .B(n_68), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_227), .B(n_71), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_211), .B(n_19), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_227), .B(n_73), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_220), .B(n_20), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_222), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_229), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_235), .B(n_28), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_203), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_195), .B(n_29), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g298 ( .A(n_212), .B(n_30), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_235), .B(n_32), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_233), .B(n_33), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_233), .B(n_34), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_213), .B(n_35), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_233), .B(n_36), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_229), .B(n_38), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_213), .B(n_44), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_230), .B(n_45), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_202), .B(n_46), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_250), .B(n_180), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_244), .A2(n_204), .B(n_199), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_277), .A2(n_230), .B(n_225), .C(n_215), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_267), .Y(n_312) );
AO21x1_ASAP7_75t_L g313 ( .A1(n_303), .A2(n_201), .B(n_205), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_242), .B(n_219), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_246), .A2(n_199), .B(n_189), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_280), .A2(n_189), .B(n_204), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_247), .A2(n_201), .B(n_205), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_245), .B(n_219), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_245), .A2(n_191), .B(n_184), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_262), .B(n_222), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_268), .B(n_219), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_266), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_294), .A2(n_180), .B(n_225), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_248), .B(n_180), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_275), .A2(n_184), .B(n_191), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_259), .B(n_180), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_282), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_241), .A2(n_217), .B(n_215), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_257), .B(n_217), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_263), .A2(n_186), .B(n_203), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_253), .A2(n_186), .B(n_206), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_279), .B(n_222), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_260), .B(n_206), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_253), .A2(n_206), .B(n_194), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_258), .A2(n_206), .B(n_194), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_292), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_274), .B(n_276), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_254), .A2(n_194), .B1(n_238), .B2(n_193), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_255), .B(n_194), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_249), .B(n_238), .Y(n_343) );
OAI321xp33_ASAP7_75t_L g344 ( .A1(n_264), .A2(n_187), .A3(n_193), .B1(n_192), .B2(n_53), .C(n_54), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_286), .B(n_192), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_258), .A2(n_187), .B(n_51), .C(n_52), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_187), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_302), .A2(n_48), .B(n_56), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_295), .A2(n_57), .B(n_58), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_272), .A2(n_59), .B(n_60), .Y(n_350) );
AOI21x1_ASAP7_75t_L g351 ( .A1(n_273), .A2(n_61), .B(n_62), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_285), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g353 ( .A1(n_281), .A2(n_76), .B(n_77), .C(n_78), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_284), .B(n_111), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_283), .A2(n_82), .B(n_83), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_288), .A2(n_86), .B(n_87), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_285), .Y(n_357) );
AOI21x1_ASAP7_75t_L g358 ( .A1(n_291), .A2(n_89), .B(n_91), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_299), .A2(n_92), .B(n_93), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_287), .B(n_94), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_287), .A2(n_96), .B(n_97), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_348), .A2(n_303), .B(n_306), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_306), .B(n_305), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_312), .B(n_290), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_317), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_358), .A2(n_304), .B(n_301), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_325), .B(n_290), .Y(n_367) );
NOR2xp67_ASAP7_75t_L g368 ( .A(n_317), .B(n_285), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_340), .A2(n_289), .B(n_256), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_349), .A2(n_307), .B(n_308), .Y(n_370) );
INVx4_ASAP7_75t_L g371 ( .A(n_317), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_359), .A2(n_308), .B(n_297), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_317), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_324), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_323), .A2(n_289), .B(n_269), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_323), .A2(n_297), .B(n_269), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_325), .Y(n_377) );
INVx4_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_313), .A2(n_243), .B(n_296), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_316), .B(n_278), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_314), .B(n_252), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_354), .A2(n_353), .B(n_361), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_338), .A2(n_240), .B(n_296), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_347), .A2(n_256), .B(n_243), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_251), .B(n_240), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_321), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_357), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_335), .A2(n_251), .B(n_293), .Y(n_389) );
NOR2x1_ASAP7_75t_R g390 ( .A(n_330), .B(n_271), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_336), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_341), .A2(n_309), .B(n_322), .Y(n_393) );
NAND3xp33_ASAP7_75t_SL g394 ( .A(n_341), .B(n_298), .C(n_99), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_332), .B(n_300), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_392), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_392), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_382), .A2(n_356), .B(n_355), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_373), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_371), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_350), .B(n_360), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_366), .A2(n_334), .B(n_318), .Y(n_402) );
CKINVDCx11_ASAP7_75t_R g403 ( .A(n_371), .Y(n_403) );
AOI21x1_ASAP7_75t_L g404 ( .A1(n_366), .A2(n_333), .B(n_337), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_393), .A2(n_311), .B(n_309), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_387), .Y(n_407) );
AOI21x1_ASAP7_75t_L g408 ( .A1(n_363), .A2(n_320), .B(n_342), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_363), .A2(n_331), .B(n_328), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_391), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_362), .A2(n_344), .B(n_346), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
OAI21x1_ASAP7_75t_L g413 ( .A1(n_362), .A2(n_315), .B(n_310), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_329), .B(n_326), .Y(n_416) );
OAI21x1_ASAP7_75t_L g417 ( .A1(n_370), .A2(n_329), .B(n_327), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_370), .A2(n_327), .B(n_343), .Y(n_418) );
AO21x2_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_332), .B(n_343), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_383), .Y(n_420) );
OAI21x1_ASAP7_75t_SL g421 ( .A1(n_380), .A2(n_98), .B(n_100), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
OAI21x1_ASAP7_75t_L g423 ( .A1(n_376), .A2(n_300), .B(n_293), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_365), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_365), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_374), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_394), .B(n_101), .Y(n_427) );
INVx6_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_415), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_419), .A2(n_364), .B1(n_381), .B2(n_377), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_410), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_415), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_410), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_420), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_381), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_420), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_419), .A2(n_364), .B1(n_393), .B2(n_367), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_422), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_414), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_422), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_422), .B(n_368), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_414), .A2(n_374), .B1(n_390), .B2(n_378), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_412), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_407), .B(n_368), .Y(n_451) );
INVx5_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_403), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_426), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_426), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_400), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_419), .A2(n_378), .B1(n_388), .B2(n_395), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
CKINVDCx11_ASAP7_75t_R g460 ( .A(n_424), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_399), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
OAI21x1_ASAP7_75t_L g463 ( .A1(n_423), .A2(n_379), .B(n_376), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_419), .B(n_378), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_425), .Y(n_466) );
INVxp33_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_399), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_423), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
OAI21x1_ASAP7_75t_L g472 ( .A1(n_404), .A2(n_379), .B(n_384), .Y(n_472) );
INVx6_ASAP7_75t_L g473 ( .A(n_428), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_400), .B(n_395), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_421), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_404), .Y(n_476) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_408), .A2(n_372), .B(n_369), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_408), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_428), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
OR2x2_ASAP7_75t_SL g484 ( .A(n_454), .B(n_390), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_449), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_441), .B(n_416), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_416), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_432), .B(n_416), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_433), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_435), .B(n_416), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_450), .B(n_417), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_435), .B(n_417), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_437), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_452), .A2(n_428), .B1(n_427), .B2(n_395), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_437), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_434), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_443), .B(n_428), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_452), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_430), .A2(n_428), .B1(n_427), .B2(n_388), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_444), .B(n_388), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_436), .A2(n_405), .B1(n_411), .B2(n_372), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_452), .A2(n_411), .B1(n_385), .B2(n_389), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_434), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_436), .A2(n_411), .B1(n_413), .B2(n_398), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_444), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_439), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_439), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_453), .B(n_102), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_438), .A2(n_411), .B1(n_413), .B2(n_398), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_446), .B(n_409), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_447), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_448), .B(n_409), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_448), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_450), .B(n_409), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_476), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_476), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_455), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_455), .B(n_413), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_442), .B(n_402), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_461), .B(n_402), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_440), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
BUFx6f_ASAP7_75t_SL g532 ( .A(n_457), .Y(n_532) );
AO31x2_ASAP7_75t_L g533 ( .A1(n_459), .A2(n_386), .A3(n_402), .B(n_401), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_452), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_468), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_481), .Y(n_540) );
NOR2xp33_ASAP7_75t_R g541 ( .A(n_453), .B(n_105), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_465), .Y(n_542) );
CKINVDCx11_ASAP7_75t_R g543 ( .A(n_460), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_465), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_440), .B(n_398), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_442), .B(n_401), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_442), .B(n_401), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_481), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_442), .B(n_106), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_475), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_475), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_108), .Y(n_554) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_463), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_469), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_478), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_457), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_482), .B(n_109), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_440), .B(n_293), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_469), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_452), .B(n_293), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_480), .B(n_300), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_462), .B(n_300), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_462), .B(n_471), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_466), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_466), .B(n_470), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_478), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_471), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_472), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_528), .B(n_470), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_522), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_528), .B(n_470), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_531), .B(n_466), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_522), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_558), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_539), .B(n_458), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_537), .A2(n_445), .B1(n_473), .B2(n_474), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_486), .B(n_474), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_451), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_504), .B(n_467), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_504), .B(n_474), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_536), .B(n_451), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_535), .Y(n_584) );
BUFx2_ASAP7_75t_R g585 ( .A(n_490), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_485), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_485), .B(n_474), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_489), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_558), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_493), .B(n_495), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_545), .B(n_480), .Y(n_591) );
BUFx4f_ASAP7_75t_SL g592 ( .A(n_490), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_545), .B(n_451), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_535), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_489), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_530), .B(n_477), .C(n_473), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_524), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_493), .B(n_477), .Y(n_598) );
BUFx12f_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_524), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_525), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_491), .B(n_473), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_505), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_536), .B(n_477), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_491), .B(n_473), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_495), .B(n_472), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_527), .B(n_498), .Y(n_609) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_505), .B(n_566), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_499), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_499), .Y(n_612) );
INVx3_ASAP7_75t_R g613 ( .A(n_541), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_483), .B(n_488), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_527), .B(n_498), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_483), .B(n_502), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_501), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_518), .B(n_521), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_547), .B(n_548), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_518), .B(n_521), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_488), .B(n_515), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_534), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_562), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_501), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_567), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_503), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_494), .B(n_510), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_567), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_525), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_532), .A2(n_550), .B1(n_566), .B2(n_500), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_487), .B(n_492), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_512), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_532), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_512), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_487), .B(n_492), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_565), .B(n_548), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_513), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_513), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_519), .B(n_520), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_565), .B(n_547), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_552), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_519), .B(n_520), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_526), .B(n_551), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_532), .A2(n_550), .B1(n_484), .B2(n_559), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_569), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_551), .B(n_553), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_569), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_526), .B(n_553), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_557), .B(n_568), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_516), .B(n_508), .C(n_511), .D(n_546), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_559), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_557), .A2(n_568), .B1(n_507), .B2(n_496), .Y(n_653) );
AND2x4_ASAP7_75t_SL g654 ( .A(n_507), .B(n_502), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_538), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_538), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_540), .B(n_549), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_542), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_494), .B(n_497), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_484), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_540), .B(n_549), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_497), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_523), .B(n_515), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_510), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_542), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_514), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_529), .B(n_523), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_514), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_529), .B(n_496), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_554), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_560), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_554), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_506), .A2(n_517), .B1(n_570), .B2(n_564), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_570), .B(n_561), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_544), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_544), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_564), .A2(n_509), .B1(n_556), .B2(n_561), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_556), .B(n_533), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_533), .B(n_552), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_533), .B(n_563), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_533), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_533), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_552), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_637), .B(n_552), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_590), .B(n_552), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_644), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_644), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_637), .B(n_555), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_646), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_590), .B(n_555), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_649), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_632), .B(n_555), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_632), .B(n_555), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_636), .B(n_555), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_662), .Y(n_696) );
AND2x4_ASAP7_75t_L g697 ( .A(n_619), .B(n_571), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_666), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_649), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_572), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_619), .B(n_571), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_641), .B(n_609), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_641), .B(n_609), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_575), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_666), .Y(n_705) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_634), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_619), .B(n_571), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_586), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_648), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_615), .B(n_636), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_645), .B(n_631), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_588), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_648), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_610), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_655), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_595), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_611), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_615), .B(n_618), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_618), .B(n_620), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_620), .B(n_669), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_617), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_624), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_581), .B(n_582), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_660), .A2(n_651), .B1(n_578), .B2(n_599), .Y(n_725) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_604), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_654), .B(n_669), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_625), .B(n_629), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_654), .B(n_591), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_625), .B(n_667), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_589), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_650), .B(n_657), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_623), .B(n_573), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_626), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_655), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_623), .B(n_573), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_573), .B(n_593), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_627), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_650), .B(n_657), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_608), .B(n_598), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_667), .B(n_574), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_633), .Y(n_742) );
INVx5_ASAP7_75t_L g743 ( .A(n_605), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_656), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_667), .B(n_577), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_608), .B(n_598), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_574), .B(n_589), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_635), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_661), .B(n_652), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_661), .B(n_638), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_574), .B(n_622), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_639), .B(n_663), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_663), .B(n_579), .Y(n_753) );
OR2x2_ASAP7_75t_L g754 ( .A(n_671), .B(n_587), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_640), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_647), .B(n_602), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_592), .Y(n_757) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_682), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_576), .B(n_580), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_643), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_647), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_583), .B(n_672), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_647), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_656), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_653), .B(n_607), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_603), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_584), .Y(n_767) );
BUFx2_ASAP7_75t_L g768 ( .A(n_592), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_614), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_678), .B(n_653), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_670), .B(n_668), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_616), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_678), .B(n_679), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_613), .B(n_578), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_606), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_621), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_628), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_664), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_679), .B(n_674), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_659), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_675), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_602), .B(n_673), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_676), .B(n_584), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_594), .B(n_630), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_594), .B(n_630), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_602), .B(n_673), .Y(n_786) );
BUFx2_ASAP7_75t_L g787 ( .A(n_599), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_585), .B(n_597), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_597), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_600), .B(n_601), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_600), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_601), .B(n_681), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_658), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_642), .B(n_674), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_658), .B(n_665), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_719), .B(n_680), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_696), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_696), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_726), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_721), .B(n_665), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_752), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_749), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_686), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_726), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_710), .B(n_674), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_687), .Y(n_806) );
NOR2x1p5_ASAP7_75t_L g807 ( .A(n_714), .B(n_596), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_710), .B(n_682), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_702), .B(n_677), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_702), .B(n_677), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_768), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_692), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_698), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_714), .Y(n_814) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_714), .B(n_642), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_703), .B(n_642), .Y(n_816) );
NAND2x1p5_ASAP7_75t_L g817 ( .A(n_757), .B(n_683), .Y(n_817) );
AND2x4_ASAP7_75t_L g818 ( .A(n_697), .B(n_683), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_699), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_703), .B(n_770), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_750), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_780), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_697), .B(n_701), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_698), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_787), .B(n_706), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_700), .Y(n_826) );
OR2x6_ASAP7_75t_L g827 ( .A(n_705), .B(n_711), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_704), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_770), .B(n_720), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_775), .B(n_755), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_775), .B(n_760), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_708), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_774), .B(n_724), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_740), .B(n_746), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_697), .B(n_701), .Y(n_835) );
AND2x2_ASAP7_75t_SL g836 ( .A(n_701), .B(n_707), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_712), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_740), .B(n_746), .Y(n_838) );
AO22x1_ASAP7_75t_L g839 ( .A1(n_743), .A2(n_774), .B1(n_707), .B2(n_788), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_753), .B(n_732), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_725), .A2(n_711), .B1(n_743), .B2(n_705), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_725), .B(n_731), .C(n_782), .Y(n_842) );
INVx2_ASAP7_75t_SL g843 ( .A(n_727), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_716), .Y(n_844) );
BUFx2_ASAP7_75t_L g845 ( .A(n_707), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_769), .B(n_772), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_717), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_741), .B(n_737), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_731), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_718), .Y(n_850) );
BUFx2_ASAP7_75t_L g851 ( .A(n_743), .Y(n_851) );
AND2x4_ASAP7_75t_L g852 ( .A(n_756), .B(n_763), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_776), .B(n_777), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_786), .B(n_739), .Y(n_854) );
NOR2x1_ASAP7_75t_L g855 ( .A(n_756), .B(n_778), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_733), .B(n_736), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_722), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_751), .B(n_779), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_785), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_723), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_779), .B(n_773), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_734), .B(n_748), .Y(n_862) );
AND2x2_ASAP7_75t_SL g863 ( .A(n_756), .B(n_729), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_766), .B(n_765), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_773), .B(n_745), .Y(n_865) );
INVxp33_ASAP7_75t_L g866 ( .A(n_759), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_743), .Y(n_867) );
OAI21xp33_ASAP7_75t_SL g868 ( .A1(n_747), .A2(n_730), .B(n_728), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_684), .B(n_688), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_689), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_762), .B(n_761), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_794), .B(n_754), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_771), .B(n_738), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_794), .B(n_685), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_742), .A2(n_690), .B1(n_695), .B2(n_693), .Y(n_875) );
AND2x4_ASAP7_75t_L g876 ( .A(n_794), .B(n_694), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_781), .B(n_790), .Y(n_877) );
INVx1_ASAP7_75t_SL g878 ( .A(n_825), .Y(n_878) );
NAND2x1p5_ASAP7_75t_L g879 ( .A(n_851), .B(n_744), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_823), .Y(n_880) );
INVx1_ASAP7_75t_SL g881 ( .A(n_811), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_862), .Y(n_882) );
AOI32xp33_ASAP7_75t_L g883 ( .A1(n_868), .A2(n_758), .A3(n_764), .B1(n_791), .B2(n_789), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_870), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_862), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_800), .B(n_792), .Y(n_886) );
NAND3xp33_ASAP7_75t_SL g887 ( .A(n_841), .B(n_783), .C(n_784), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_830), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_830), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_831), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_842), .A2(n_758), .B1(n_735), .B2(n_744), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_845), .B(n_715), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_831), .Y(n_893) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_799), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_810), .B(n_793), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_797), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_868), .B(n_715), .Y(n_897) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_849), .Y(n_898) );
INVxp67_ASAP7_75t_L g899 ( .A(n_798), .Y(n_899) );
INVx1_ASAP7_75t_SL g900 ( .A(n_863), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_872), .B(n_735), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_804), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_854), .B(n_689), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_822), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_813), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_872), .B(n_691), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_846), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_836), .B(n_691), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_846), .Y(n_909) );
AOI33xp33_ASAP7_75t_L g910 ( .A1(n_802), .A2(n_709), .A3(n_713), .B1(n_767), .B2(n_795), .B3(n_821), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_853), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_834), .B(n_709), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_796), .B(n_713), .Y(n_913) );
AND2x4_ASAP7_75t_L g914 ( .A(n_823), .B(n_767), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_853), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_824), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_826), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_827), .A2(n_841), .B1(n_842), .B2(n_866), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_828), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_838), .B(n_835), .Y(n_920) );
XNOR2xp5_ASAP7_75t_L g921 ( .A(n_827), .B(n_843), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_835), .Y(n_922) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_827), .A2(n_809), .B1(n_855), .B2(n_867), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_832), .Y(n_924) );
INVx3_ASAP7_75t_L g925 ( .A(n_814), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_900), .A2(n_855), .B1(n_814), .B2(n_817), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_879), .Y(n_927) );
OA22x2_ASAP7_75t_L g928 ( .A1(n_918), .A2(n_852), .B1(n_801), .B2(n_864), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_882), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g930 ( .A(n_878), .B(n_833), .Y(n_930) );
INVx2_ASAP7_75t_SL g931 ( .A(n_881), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_910), .B(n_854), .Y(n_932) );
OAI21xp33_ASAP7_75t_SL g933 ( .A1(n_883), .A2(n_807), .B(n_861), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_885), .Y(n_934) );
O2A1O1Ixp33_ASAP7_75t_L g935 ( .A1(n_923), .A2(n_873), .B(n_820), .C(n_844), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_907), .B(n_829), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_909), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_891), .B(n_839), .C(n_875), .Y(n_938) );
OAI222xp33_ASAP7_75t_L g939 ( .A1(n_923), .A2(n_875), .B1(n_840), .B2(n_815), .C1(n_865), .C2(n_808), .Y(n_939) );
AOI31xp33_ASAP7_75t_L g940 ( .A1(n_921), .A2(n_856), .A3(n_805), .B(n_816), .Y(n_940) );
OAI322xp33_ASAP7_75t_L g941 ( .A1(n_897), .A2(n_877), .A3(n_806), .B1(n_812), .B2(n_803), .C1(n_819), .C2(n_837), .Y(n_941) );
AOI211xp5_ASAP7_75t_L g942 ( .A1(n_887), .A2(n_818), .B(n_852), .C(n_860), .Y(n_942) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_894), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_894), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_879), .Y(n_945) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_880), .B(n_858), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_911), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_898), .A2(n_818), .B(n_876), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_884), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_898), .A2(n_876), .B(n_874), .Y(n_950) );
OAI21xp33_ASAP7_75t_L g951 ( .A1(n_891), .A2(n_874), .B(n_859), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_933), .A2(n_880), .B1(n_922), .B2(n_925), .C(n_893), .Y(n_952) );
AOI221x1_ASAP7_75t_L g953 ( .A1(n_938), .A2(n_925), .B1(n_889), .B2(n_888), .C(n_890), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_932), .B(n_910), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_935), .A2(n_922), .B1(n_925), .B2(n_915), .C(n_899), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_939), .A2(n_899), .B1(n_904), .B2(n_917), .C(n_919), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_939), .A2(n_924), .B1(n_896), .B2(n_895), .C(n_903), .Y(n_957) );
NOR2xp67_ASAP7_75t_L g958 ( .A(n_943), .B(n_916), .Y(n_958) );
OAI32xp33_ASAP7_75t_L g959 ( .A1(n_928), .A2(n_916), .A3(n_920), .B1(n_886), .B2(n_913), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_943), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_944), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_936), .B(n_847), .Y(n_962) );
OAI21xp5_ASAP7_75t_L g963 ( .A1(n_928), .A2(n_914), .B(n_908), .Y(n_963) );
AOI222xp33_ASAP7_75t_L g964 ( .A1(n_944), .A2(n_850), .B1(n_857), .B2(n_902), .C1(n_905), .C2(n_892), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_931), .B(n_901), .Y(n_965) );
NAND2xp33_ASAP7_75t_L g966 ( .A(n_963), .B(n_951), .Y(n_966) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_959), .A2(n_941), .B1(n_926), .B2(n_930), .C(n_940), .Y(n_967) );
NAND2x1_ASAP7_75t_L g968 ( .A(n_958), .B(n_950), .Y(n_968) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_956), .A2(n_942), .B1(n_930), .B2(n_948), .C(n_927), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_954), .B(n_937), .Y(n_970) );
NAND4xp75_ASAP7_75t_L g971 ( .A(n_953), .B(n_945), .C(n_947), .D(n_934), .Y(n_971) );
NOR4xp25_ASAP7_75t_L g972 ( .A(n_952), .B(n_926), .C(n_929), .D(n_949), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_960), .Y(n_973) );
NOR2x1_ASAP7_75t_SL g974 ( .A(n_971), .B(n_961), .Y(n_974) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_967), .B(n_957), .C(n_955), .Y(n_975) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_972), .A2(n_964), .B(n_965), .C(n_962), .Y(n_976) );
NOR2xp67_ASAP7_75t_L g977 ( .A(n_969), .B(n_902), .Y(n_977) );
AOI21x1_ASAP7_75t_L g978 ( .A1(n_977), .A2(n_968), .B(n_973), .Y(n_978) );
NOR2x1_ASAP7_75t_L g979 ( .A(n_975), .B(n_966), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_976), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_979), .B(n_974), .Y(n_981) );
NOR2x1p5_ASAP7_75t_L g982 ( .A(n_980), .B(n_970), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_981), .B(n_964), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_982), .A2(n_946), .B1(n_978), .B2(n_914), .Y(n_984) );
XNOR2x1_ASAP7_75t_L g985 ( .A(n_983), .B(n_914), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_984), .B(n_905), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_986), .Y(n_987) );
AOI21xp33_ASAP7_75t_L g988 ( .A1(n_987), .A2(n_985), .B(n_884), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_988), .Y(n_989) );
XNOR2xp5_ASAP7_75t_L g990 ( .A(n_989), .B(n_906), .Y(n_990) );
OR2x6_ASAP7_75t_L g991 ( .A(n_990), .B(n_912), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_991), .B(n_848), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_992), .A2(n_871), .B(n_869), .Y(n_993) );
endmodule