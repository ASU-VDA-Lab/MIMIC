module fake_jpeg_21400_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_30),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_5),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_0),
.B(n_1),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_54),
.B(n_45),
.C(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_36),
.B1(n_43),
.B2(n_35),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_28),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_24),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_56),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_68),
.Y(n_102)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_15),
.B1(n_2),
.B2(n_9),
.Y(n_111)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_81),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_89),
.B(n_1),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_21),
.B(n_18),
.C(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_76),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_15),
.B1(n_16),
.B2(n_3),
.Y(n_105)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_26),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_91),
.B1(n_44),
.B2(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_17),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_24),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_24),
.C(n_16),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_21),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_111),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_16),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_107),
.B(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_66),
.B1(n_90),
.B2(n_77),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_79),
.B1(n_7),
.B2(n_77),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_2),
.B(n_4),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_83),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_2),
.B(n_4),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_74),
.B1(n_80),
.B2(n_75),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_87),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_71),
.C(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_125),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_129),
.B1(n_105),
.B2(n_99),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_126),
.Y(n_133)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_131),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_111),
.B(n_109),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_128),
.A2(n_114),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_146),
.B(n_120),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_111),
.B1(n_128),
.B2(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_72),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_120),
.B1(n_123),
.B2(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_92),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_99),
.B(n_111),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_117),
.B1(n_114),
.B2(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_151),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_157),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_153),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_121),
.B(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_97),
.B1(n_94),
.B2(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_162),
.Y(n_168)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

XNOR2x2_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_164),
.A2(n_153),
.B1(n_141),
.B2(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_143),
.C(n_151),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_141),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_167),
.C(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_173),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_160),
.C(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_161),
.B(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_182),
.B1(n_174),
.B2(n_97),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_150),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_183),
.B(n_180),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_186),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_7),
.Y(n_189)
);


endmodule