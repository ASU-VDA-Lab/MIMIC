module real_jpeg_3847_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_178;
wire n_67;
wire n_79;
wire n_76;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_1),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_1),
.A2(n_88),
.B1(n_103),
.B2(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_3),
.A2(n_42),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_42),
.B1(n_95),
.B2(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_4),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_94),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_94),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_177),
.B1(n_178),
.B2(n_182),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_5),
.Y(n_182)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_9),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_9),
.A2(n_132),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_205),
.C(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_9),
.B(n_121),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_9),
.B(n_152),
.Y(n_244)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_12),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_189),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_187),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_142),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_16),
.B(n_142),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_69),
.C(n_104),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_17),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_47),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_18),
.B(n_47),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_28),
.B(n_31),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_20),
.A2(n_32),
.B1(n_176),
.B2(n_183),
.Y(n_175)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_22),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_30),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_31),
.A2(n_237),
.B(n_243),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_32),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_32),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_34),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_37),
.B(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_44),
.Y(n_177)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.A3(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_50),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_50),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_54),
.Y(n_199)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_69),
.A2(n_104),
.B1(n_105),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_69),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_82),
.B1(n_91),
.B2(n_98),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_98),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_70),
.A2(n_146),
.B(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_71),
.B(n_147),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_82),
.A2(n_91),
.B(n_224),
.Y(n_223)
);

AOI22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_88),
.B(n_231),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_128),
.B(n_134),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_121),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_121),
.Y(n_141)
);

AO22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_132),
.B(n_133),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_132),
.A2(n_217),
.B(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_156),
.B(n_162),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_154),
.B2(n_186),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_175),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_255),
.B(n_260),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_227),
.B(n_254),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_209),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_193),
.A2(n_200),
.B1(n_201),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_221),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_210),
.B(n_222),
.C(n_226),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_217),
.B(n_218),
.Y(n_210)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_246),
.B(n_253),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_235),
.B(n_245),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_244),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_251),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);


endmodule