module fake_jpeg_15456_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_5),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_46),
.C(n_58),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_69),
.C(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_47),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_65),
.B(n_48),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_60),
.B(n_63),
.Y(n_74)
);

OAI31xp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_75),
.A3(n_66),
.B(n_64),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_66),
.B(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_77),
.B(n_43),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_61),
.A3(n_63),
.B1(n_62),
.B2(n_37),
.C1(n_58),
.C2(n_23),
.Y(n_78)
);

OAI221xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_42),
.B1(n_20),
.B2(n_21),
.C(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_81),
.A3(n_62),
.B1(n_37),
.B2(n_40),
.C1(n_35),
.C2(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_39),
.B1(n_34),
.B2(n_50),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_39),
.Y(n_86)
);


endmodule