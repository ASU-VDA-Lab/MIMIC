module fake_jpeg_11305_n_185 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_86),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_65),
.B1(n_57),
.B2(n_53),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_97),
.B1(n_72),
.B2(n_67),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_65),
.B1(n_57),
.B2(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_64),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_125),
.B1(n_24),
.B2(n_45),
.Y(n_137)
);

AOI22x1_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_76),
.B1(n_75),
.B2(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_117),
.B1(n_62),
.B2(n_54),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

CKINVDCx10_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_76),
.B1(n_63),
.B2(n_67),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_51),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_68),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_2),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_52),
.B1(n_69),
.B2(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_1),
.B(n_2),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_12),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_1),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_140),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_23),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_28),
.CI(n_37),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_3),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_4),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_30),
.C(n_44),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_48),
.C(n_16),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_33),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_147),
.B(n_11),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_148),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_155),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_18),
.B(n_19),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_161),
.B(n_162),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_20),
.C(n_27),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_38),
.C(n_42),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_137),
.B1(n_139),
.B2(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_173),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_177),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_133),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_170),
.C(n_167),
.Y(n_179)
);

AO221x1_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_142),
.B1(n_152),
.B2(n_150),
.C(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_170),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_178),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_181),
.B(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_158),
.B1(n_174),
.B2(n_157),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_146),
.B(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_162),
.Y(n_185)
);


endmodule