module fake_jpeg_9706_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_29),
.B1(n_18),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_59),
.B1(n_39),
.B2(n_20),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_29),
.B1(n_43),
.B2(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_29),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_24),
.B1(n_20),
.B2(n_34),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_0),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_62),
.C(n_48),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_77),
.C(n_78),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_90),
.B1(n_92),
.B2(n_26),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_53),
.B1(n_66),
.B2(n_45),
.Y(n_97)
);

XOR2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_37),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_85),
.B1(n_30),
.B2(n_25),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_87),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_41),
.B1(n_38),
.B2(n_18),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_104),
.B1(n_112),
.B2(n_121),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_111),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_46),
.A3(n_37),
.B1(n_35),
.B2(n_27),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_78),
.B(n_21),
.C(n_35),
.D(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_115),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_113),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_79),
.B1(n_89),
.B2(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_30),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_22),
.B1(n_50),
.B2(n_25),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_71),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_84),
.B1(n_22),
.B2(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_35),
.B(n_37),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_131),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_78),
.C(n_86),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_96),
.C(n_106),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_15),
.C(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_146),
.B1(n_41),
.B2(n_38),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_87),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_82),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_41),
.B1(n_38),
.B2(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_52),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_99),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_120),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_159),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_113),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_155),
.C(n_180),
.Y(n_191)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_106),
.B1(n_99),
.B2(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_167),
.B1(n_143),
.B2(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_21),
.B(n_31),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_170),
.B(n_132),
.Y(n_190)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_152),
.B1(n_179),
.B2(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_38),
.B1(n_31),
.B2(n_28),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_100),
.B(n_116),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_137),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

BUFx4f_ASAP7_75t_SL g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_173),
.B(n_176),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_31),
.C(n_28),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_188),
.B1(n_207),
.B2(n_167),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_194),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_163),
.B(n_157),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_130),
.C(n_135),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_196),
.C(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_133),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_124),
.A3(n_138),
.B1(n_128),
.B2(n_131),
.C1(n_125),
.C2(n_31),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_159),
.Y(n_218)
);

OR2x2_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_124),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_178),
.B(n_172),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_124),
.C(n_100),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_100),
.C(n_15),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_207),
.C(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_217),
.B(n_195),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_180),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_212),
.C(n_156),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_215),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_224),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_165),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_176),
.B1(n_168),
.B2(n_161),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_221),
.B1(n_160),
.B2(n_6),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_161),
.B(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

HAxp5_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_190),
.CON(n_221),
.SN(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_172),
.A3(n_177),
.B1(n_5),
.B2(n_6),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_196),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_2),
.CI(n_4),
.CON(n_224),
.SN(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_227),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_4),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_7),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_199),
.B1(n_193),
.B2(n_186),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_246),
.B1(n_224),
.B2(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_217),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_205),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_241),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_198),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_249),
.C(n_227),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_223),
.B(n_231),
.C(n_229),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_7),
.C(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_259),
.C(n_260),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_261),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_230),
.C(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_262),
.C(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_213),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_208),
.C(n_220),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_221),
.CI(n_224),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_239),
.C(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_247),
.C(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_256),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_259),
.B(n_11),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_235),
.B1(n_242),
.B2(n_244),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_12),
.C(n_13),
.Y(n_292)
);

OAI211xp5_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_285),
.B(n_286),
.C(n_275),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_251),
.B1(n_255),
.B2(n_252),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_284),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_270),
.B(n_268),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_10),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_12),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_267),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_272),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_292),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_282),
.A2(n_13),
.B(n_14),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_283),
.B(n_284),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_295),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_299),
.B(n_300),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_294),
.C(n_298),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_297),
.Y(n_304)
);


endmodule