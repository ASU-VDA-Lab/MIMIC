module fake_jpeg_20736_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_22),
.B(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_68),
.B1(n_34),
.B2(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_34),
.B1(n_19),
.B2(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_17),
.B(n_35),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_75),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_86),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_43),
.B1(n_47),
.B2(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NAND2x1_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_38),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_31),
.B1(n_23),
.B2(n_24),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_32),
.B1(n_24),
.B2(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_26),
.B1(n_35),
.B2(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_90),
.B1(n_36),
.B2(n_21),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_26),
.B1(n_35),
.B2(n_27),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_44),
.B1(n_36),
.B2(n_30),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_92),
.Y(n_131)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_95),
.Y(n_122)
);

AND2x4_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_22),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_50),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_50),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_98),
.B1(n_92),
.B2(n_80),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_46),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_128),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_126),
.B1(n_80),
.B2(n_117),
.Y(n_154)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_85),
.B1(n_78),
.B2(n_36),
.Y(n_159)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_133),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_36),
.B1(n_30),
.B2(n_28),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_116),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_80),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_138),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_81),
.B(n_75),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_75),
.B(n_81),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_94),
.B(n_75),
.C(n_86),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_131),
.B1(n_134),
.B2(n_123),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_94),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_91),
.B1(n_89),
.B2(n_100),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_105),
.B1(n_115),
.B2(n_106),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_79),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_79),
.B(n_88),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_163),
.B1(n_105),
.B2(n_123),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_159),
.B1(n_133),
.B2(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_104),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_192),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_106),
.B1(n_134),
.B2(n_131),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_111),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_194),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_185),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_107),
.B1(n_135),
.B2(n_110),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_124),
.B(n_13),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_163),
.B(n_138),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_108),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_139),
.B(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_110),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_111),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_201),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_206),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_215),
.B1(n_218),
.B2(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_137),
.B1(n_146),
.B2(n_141),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_207),
.B1(n_226),
.B2(n_185),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_161),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_173),
.C(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_211),
.C(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_166),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_137),
.B1(n_141),
.B2(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_145),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_186),
.C(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_203),
.B1(n_168),
.B2(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_141),
.B1(n_156),
.B2(n_148),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_174),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_153),
.B(n_113),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_111),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_108),
.C(n_110),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_21),
.B(n_28),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_176),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_175),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_233),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_211),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_179),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_241),
.B1(n_243),
.B2(n_207),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_215),
.B(n_209),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_168),
.B1(n_178),
.B2(n_177),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_188),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_247),
.C(n_217),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_188),
.C(n_177),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_195),
.A2(n_107),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_206),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_253),
.B(n_258),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_234),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_268),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_263),
.B1(n_264),
.B2(n_270),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_200),
.B1(n_224),
.B2(n_223),
.Y(n_264)
);

NOR4xp25_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_210),
.C(n_219),
.D(n_204),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_251),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_208),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_240),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_219),
.B1(n_210),
.B2(n_208),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_227),
.A2(n_225),
.B(n_202),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_263),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_202),
.B(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_236),
.C(n_230),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_277),
.C(n_280),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_236),
.C(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_246),
.C(n_229),
.Y(n_280)
);

AOI22x1_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_242),
.B1(n_261),
.B2(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_239),
.B1(n_235),
.B2(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_285)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_28),
.C(n_8),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_292),
.C(n_254),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_0),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_15),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_14),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_13),
.C(n_12),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_267),
.B1(n_265),
.B2(n_262),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_304),
.B1(n_283),
.B2(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_270),
.C(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_291),
.C(n_277),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_290),
.A2(n_282),
.B(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_273),
.B(n_14),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_0),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_0),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_289),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_319),
.C(n_306),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_292),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_312),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_318),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_291),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_297),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_0),
.C(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_324),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_307),
.B1(n_299),
.B2(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_294),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_308),
.C(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_298),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_315),
.B1(n_305),
.B2(n_310),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_335),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_323),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_334),
.C(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

NOR2x1_ASAP7_75t_R g337 ( 
.A(n_330),
.B(n_325),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.C(n_338),
.Y(n_341)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_326),
.B(n_329),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_321),
.A3(n_314),
.B1(n_293),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_2),
.Y(n_344)
);

OAI321xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_345)
);

OAI31xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_3),
.A3(n_4),
.B(n_6),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_3),
.Y(n_347)
);


endmodule