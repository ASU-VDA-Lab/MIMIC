module fake_netlist_6_4349_n_1858 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1858);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1858;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_139),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_70),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_74),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_57),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_68),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_9),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_66),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_59),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_28),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_77),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_92),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_55),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_125),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_149),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_86),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_67),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_18),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_103),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_55),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_89),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_21),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_130),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_41),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_45),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_33),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_107),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_152),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_3),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_23),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_60),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_188),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_109),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_98),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_114),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_113),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_10),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_20),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_30),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_138),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_169),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_166),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_54),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_116),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_75),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_111),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_148),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_117),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_53),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_45),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_83),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_105),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_24),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_165),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_61),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_164),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_62),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_140),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_104),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_51),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_37),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_156),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_157),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_168),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_34),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_187),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_163),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_155),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_11),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_43),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_64),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_172),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_44),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_53),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_58),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_120),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_112),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_123),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_41),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_141),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_9),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_177),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_158),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_96),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_16),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_27),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_22),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_29),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_108),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_69),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_16),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_54),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_189),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_0),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_49),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_174),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_178),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_161),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_39),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_71),
.Y(n_338)
);

BUFx8_ASAP7_75t_SL g339 ( 
.A(n_170),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_183),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_12),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_91),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_94),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_100),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_162),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_133),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_76),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_37),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_21),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_26),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_40),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_124),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_31),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_40),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_57),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_59),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_38),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_151),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_176),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_46),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_42),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_136),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_36),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_46),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_144),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_58),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_118),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_93),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_42),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_102),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_8),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_15),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_43),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_185),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_154),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_192),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_88),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_119),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_179),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_126),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_4),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_44),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_28),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_101),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_203),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_219),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_210),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_337),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_322),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_278),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_241),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_260),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_240),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_294),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_260),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_260),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_260),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_198),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_260),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_290),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_290),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_299),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_242),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_290),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_290),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_245),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_308),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_246),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_246),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_237),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_290),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_310),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_353),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_310),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_348),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_310),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_310),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_310),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_205),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_339),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_225),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_234),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_211),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_234),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_226),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_238),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_250),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_223),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g449 ( 
.A(n_321),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_207),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_253),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_207),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_255),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_214),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_212),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_280),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_283),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_256),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_236),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_266),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_204),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_236),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_271),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_204),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_217),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_212),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_204),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_211),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_257),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_211),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_361),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_257),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_261),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_199),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_288),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_195),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_293),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_196),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_273),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_208),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_297),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_231),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_306),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_321),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_439),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_392),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_411),
.B(n_217),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_398),
.A2(n_386),
.B1(n_374),
.B2(n_230),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_251),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_389),
.B(n_223),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_389),
.B(n_223),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_391),
.B(n_251),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_429),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_465),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_388),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_461),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_197),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_476),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_465),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_403),
.A2(n_259),
.B1(n_292),
.B2(n_384),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_441),
.B(n_197),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_418),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_397),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_461),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_200),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_399),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_478),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_401),
.Y(n_537)
);

CKINVDCx6p67_ASAP7_75t_R g538 ( 
.A(n_473),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_402),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_436),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_443),
.B(n_218),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_482),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_436),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_468),
.B(n_287),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_464),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_402),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_404),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_470),
.B(n_200),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_405),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_405),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_467),
.A2(n_324),
.B(n_312),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_432),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_435),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_423),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_449),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_556),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_556),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_417),
.C(n_404),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_488),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_496),
.A2(n_431),
.B1(n_400),
.B2(n_395),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_417),
.Y(n_569)
);

NAND2x1_ASAP7_75t_L g570 ( 
.A(n_556),
.B(n_287),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_531),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_420),
.Y(n_573)
);

AO22x2_ASAP7_75t_L g574 ( 
.A1(n_493),
.A2(n_311),
.B1(n_372),
.B2(n_243),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_490),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_563),
.B(n_412),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_563),
.B(n_458),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_485),
.A2(n_422),
.B1(n_311),
.B2(n_372),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_525),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_560),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_520),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_510),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_563),
.B(n_458),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_531),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_517),
.B(n_460),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_488),
.Y(n_589)
);

AND3x1_ASAP7_75t_L g590 ( 
.A(n_523),
.B(n_243),
.C(n_341),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_490),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_489),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_547),
.B(n_495),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_529),
.Y(n_596)
);

BUFx6f_ASAP7_75t_SL g597 ( 
.A(n_560),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_485),
.B(n_460),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_529),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_515),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_485),
.A2(n_425),
.B1(n_455),
.B2(n_452),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_497),
.Y(n_602)
);

INVx8_ASAP7_75t_L g603 ( 
.A(n_504),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_497),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_515),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_534),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_495),
.A2(n_466),
.B1(n_358),
.B2(n_375),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_517),
.B(n_463),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_495),
.B(n_463),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_552),
.B(n_479),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_496),
.A2(n_390),
.B1(n_394),
.B2(n_479),
.Y(n_612)
);

AOI21x1_ASAP7_75t_L g613 ( 
.A1(n_492),
.A2(n_537),
.B(n_534),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_499),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_499),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_534),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_449),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_537),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_523),
.A2(n_501),
.B1(n_385),
.B2(n_367),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_526),
.Y(n_623)
);

OAI22xp33_ASAP7_75t_L g624 ( 
.A1(n_501),
.A2(n_295),
.B1(n_296),
.B2(n_279),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_503),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_490),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_526),
.B(n_449),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_532),
.B(n_484),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_537),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_490),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_545),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_490),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_424),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_484),
.B(n_394),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_510),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_539),
.B(n_448),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_549),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_503),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_549),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_505),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_493),
.B(n_448),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_553),
.B(n_221),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_535),
.B(n_454),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_502),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_505),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_492),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_502),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_492),
.A2(n_387),
.B(n_344),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_504),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_525),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_561),
.B(n_471),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_502),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_553),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_554),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_554),
.B(n_224),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_492),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_492),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_525),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_558),
.B(n_426),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_535),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_562),
.B(n_270),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_525),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_562),
.B(n_270),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_525),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_525),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_562),
.B(n_270),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_506),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_504),
.A2(n_359),
.B1(n_387),
.B2(n_344),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_538),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_512),
.Y(n_682)
);

BUFx6f_ASAP7_75t_SL g683 ( 
.A(n_504),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_512),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_504),
.A2(n_451),
.B1(n_438),
.B2(n_440),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_558),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_538),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_538),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_528),
.B(n_248),
.Y(n_689)
);

INVxp33_ASAP7_75t_SL g690 ( 
.A(n_487),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_528),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_562),
.B(n_281),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_486),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_528),
.B(n_533),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_502),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_486),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_512),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_491),
.Y(n_698)
);

AND3x1_ASAP7_75t_L g699 ( 
.A(n_491),
.B(n_428),
.C(n_445),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_498),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_494),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_498),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_500),
.B(n_303),
.C(n_272),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_528),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_500),
.Y(n_705)
);

AO21x2_ASAP7_75t_L g706 ( 
.A1(n_508),
.A2(n_228),
.B(n_227),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_562),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_494),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_508),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_509),
.B(n_447),
.C(n_446),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_504),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_509),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_600),
.B(n_201),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_711),
.B(n_229),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_594),
.A2(n_408),
.B1(n_416),
.B2(n_407),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_600),
.B(n_528),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_652),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_666),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_606),
.B(n_201),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_567),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_606),
.B(n_528),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_623),
.B(n_533),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_623),
.B(n_569),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_666),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_594),
.B(n_533),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_611),
.B(n_202),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_598),
.B(n_533),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_636),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_594),
.B(n_533),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_594),
.B(n_541),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_712),
.B(n_541),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_608),
.A2(n_453),
.B1(n_456),
.B2(n_457),
.C(n_265),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_667),
.B(n_541),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_652),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_686),
.B(n_541),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_709),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_667),
.B(n_541),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_637),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_686),
.B(n_541),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_589),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_589),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_592),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_634),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_572),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_620),
.B(n_555),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_628),
.A2(n_421),
.B1(n_427),
.B2(n_433),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_689),
.A2(n_522),
.B(n_507),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_564),
.B(n_555),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_634),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_573),
.B(n_475),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_564),
.B(n_555),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_622),
.B(n_555),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_593),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_565),
.B(n_555),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_481),
.C(n_477),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_612),
.B(n_481),
.C(n_477),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_206),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_593),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_669),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_565),
.B(n_555),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_576),
.A2(n_483),
.B(n_334),
.C(n_232),
.Y(n_764)
);

O2A1O1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_576),
.A2(n_540),
.B(n_511),
.C(n_514),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_572),
.B(n_434),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_624),
.B(n_483),
.C(n_301),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_659),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_627),
.B(n_513),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_571),
.A2(n_504),
.B1(n_204),
.B2(n_378),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_669),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_577),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_711),
.B(n_204),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_613),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_647),
.B(n_513),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_628),
.A2(n_320),
.B1(n_286),
.B2(n_282),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_665),
.B(n_513),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_587),
.B(n_206),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_693),
.B(n_513),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_696),
.B(n_513),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_595),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_696),
.B(n_698),
.Y(n_782)
);

OAI22x1_ASAP7_75t_L g783 ( 
.A1(n_646),
.A2(n_292),
.B1(n_349),
.B2(n_350),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_587),
.A2(n_574),
.B1(n_590),
.B2(n_648),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_698),
.B(n_530),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_595),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_262),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_700),
.B(n_530),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_568),
.B(n_204),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_674),
.B(n_268),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_616),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_628),
.A2(n_384),
.B1(n_357),
.B2(n_356),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_702),
.B(n_530),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_616),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_613),
.B(n_204),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_702),
.B(n_530),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_588),
.B(n_609),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_628),
.B(n_209),
.Y(n_799)
);

AND3x4_ASAP7_75t_L g800 ( 
.A(n_703),
.B(n_350),
.C(n_349),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_699),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_578),
.A2(n_331),
.B1(n_314),
.B2(n_276),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_601),
.B(n_616),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_705),
.B(n_530),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_638),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_586),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_602),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_602),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_583),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_585),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_675),
.B(n_548),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_574),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_586),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_574),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_597),
.A2(n_291),
.B1(n_275),
.B2(n_269),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_694),
.B(n_204),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_596),
.B(n_378),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_706),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_597),
.B(n_209),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_677),
.B(n_548),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_603),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_681),
.B(n_691),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_605),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_605),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_596),
.B(n_548),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_599),
.B(n_378),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_597),
.B(n_580),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_604),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_583),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_599),
.B(n_548),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_570),
.A2(n_655),
.B(n_707),
.C(n_673),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_607),
.B(n_378),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_607),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_604),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_639),
.B(n_548),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_642),
.B(n_551),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_642),
.B(n_551),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_643),
.B(n_551),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_643),
.B(n_551),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_644),
.B(n_378),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_644),
.B(n_662),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_662),
.B(n_378),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_614),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_663),
.B(n_551),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_663),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_664),
.B(n_494),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_664),
.B(n_668),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_668),
.B(n_494),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_SL g849 ( 
.A(n_690),
.B(n_281),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_581),
.A2(n_522),
.B(n_507),
.Y(n_850)
);

OAI22xp33_ASAP7_75t_L g851 ( 
.A1(n_570),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_701),
.B(n_378),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_701),
.B(n_378),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_615),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_690),
.B(n_281),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_704),
.B(n_494),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_704),
.B(n_511),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_603),
.B(n_233),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_618),
.B(n_514),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_621),
.B(n_516),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_629),
.B(n_516),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_631),
.B(n_518),
.Y(n_863)
);

NOR2x1p5_ASAP7_75t_L g864 ( 
.A(n_687),
.B(n_352),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_671),
.A2(n_335),
.B1(n_239),
.B2(n_235),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_615),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_676),
.B(n_692),
.Y(n_867)
);

AO221x1_ASAP7_75t_L g868 ( 
.A1(n_574),
.A2(n_289),
.B1(n_284),
.B2(n_285),
.C(n_298),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_723),
.B(n_635),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_718),
.Y(n_870)
);

NOR2x1p5_ASAP7_75t_L g871 ( 
.A(n_791),
.B(n_687),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_SL g872 ( 
.A(n_793),
.B(n_357),
.C(n_355),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_747),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_774),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_812),
.A2(n_706),
.B1(n_679),
.B2(n_683),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_724),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_723),
.B(n_706),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_766),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_805),
.B(n_575),
.Y(n_879)
);

OAI22xp33_ASAP7_75t_L g880 ( 
.A1(n_812),
.A2(n_632),
.B1(n_670),
.B2(n_680),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_737),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_768),
.B(n_632),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_798),
.B(n_688),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_728),
.B(n_670),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_823),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_717),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_740),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_717),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_772),
.B(n_814),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_868),
.A2(n_683),
.B1(n_504),
.B2(n_381),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_809),
.B(n_710),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_823),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_774),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_821),
.B(n_657),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_805),
.B(n_575),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_829),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_726),
.B(n_575),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_726),
.B(n_626),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_824),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_829),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_824),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_821),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_774),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_792),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_821),
.Y(n_905)
);

OR2x4_ASAP7_75t_L g906 ( 
.A(n_827),
.B(n_274),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_806),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_720),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_760),
.B(n_630),
.Y(n_909)
);

HB1xp67_ASAP7_75t_SL g910 ( 
.A(n_791),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_713),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_855),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_801),
.B(n_658),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_818),
.A2(n_683),
.B1(n_504),
.B2(n_346),
.Y(n_914)
);

AND3x2_ASAP7_75t_SL g915 ( 
.A(n_793),
.B(n_584),
.C(n_0),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_762),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_813),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_760),
.B(n_713),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_774),
.B(n_581),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_719),
.B(n_782),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_821),
.B(n_657),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_719),
.B(n_630),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_833),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_716),
.B(n_721),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_722),
.B(n_630),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_795),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_798),
.B(n_581),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_735),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_810),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_867),
.A2(n_685),
.B1(n_316),
.B2(n_370),
.Y(n_930)
);

AO22x1_ASAP7_75t_L g931 ( 
.A1(n_800),
.A2(n_323),
.B1(n_313),
.B2(n_307),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_753),
.B(n_633),
.Y(n_932)
);

BUFx4_ASAP7_75t_L g933 ( 
.A(n_771),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_778),
.B(n_746),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_739),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_778),
.B(n_827),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_795),
.B(n_603),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_752),
.B(n_658),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_745),
.B(n_769),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_725),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_845),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_729),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_727),
.B(n_633),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_867),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_787),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_727),
.B(n_649),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_803),
.A2(n_783),
.B1(n_799),
.B2(n_819),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_742),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_799),
.B(n_442),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_789),
.A2(n_658),
.B1(n_708),
.B2(n_603),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_715),
.B(n_444),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_755),
.A2(n_504),
.B1(n_340),
.B2(n_327),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_714),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_784),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_755),
.A2(n_315),
.B1(n_318),
.B2(n_684),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_730),
.B(n_657),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_784),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_789),
.A2(n_708),
.B1(n_649),
.B2(n_695),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_748),
.B(n_649),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_849),
.B(n_213),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_731),
.A2(n_619),
.B(n_591),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_751),
.B(n_653),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_743),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_784),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_864),
.B(n_444),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_754),
.B(n_653),
.Y(n_966)
);

NOR3xp33_ASAP7_75t_SL g967 ( 
.A(n_851),
.B(n_317),
.C(n_305),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_749),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_757),
.A2(n_619),
.B(n_591),
.Y(n_969)
);

NOR2x1_ASAP7_75t_R g970 ( 
.A(n_773),
.B(n_213),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_763),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_744),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_759),
.B(n_459),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_819),
.B(n_215),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_776),
.B(n_851),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_733),
.B(n_326),
.C(n_325),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_854),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_764),
.A2(n_518),
.B(n_521),
.C(n_524),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_802),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_714),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_775),
.B(n_653),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_787),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_773),
.A2(n_695),
.B1(n_244),
.B2(n_247),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_815),
.Y(n_984)
);

CKINVDCx8_ASAP7_75t_R g985 ( 
.A(n_787),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_787),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_841),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_816),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_865),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_767),
.B(n_462),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_777),
.B(n_695),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_736),
.B(n_591),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_741),
.B(n_657),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_732),
.B(n_591),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_841),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_SL g996 ( 
.A(n_764),
.B(n_330),
.C(n_329),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_SL g997 ( 
.A(n_770),
.B(n_215),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_734),
.A2(n_365),
.B1(n_249),
.B2(n_252),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_756),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_817),
.B(n_826),
.Y(n_1000)
);

AO21x1_ASAP7_75t_L g1001 ( 
.A1(n_796),
.A2(n_655),
.B(n_524),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_817),
.B(n_462),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_787),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_761),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_779),
.B(n_619),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_780),
.B(n_657),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_790),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_785),
.B(n_619),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_788),
.B(n_619),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_790),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_790),
.Y(n_1011)
);

AND2x6_ASAP7_75t_SL g1012 ( 
.A(n_860),
.B(n_469),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_758),
.B(n_216),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_826),
.B(n_469),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_794),
.B(n_333),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_781),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_797),
.B(n_363),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_786),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_847),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_816),
.B(n_832),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_804),
.B(n_216),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_807),
.B(n_640),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_808),
.B(n_640),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_828),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_834),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_843),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_866),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_831),
.B(n_640),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_770),
.A2(n_697),
.B1(n_684),
.B2(n_682),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_832),
.B(n_472),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_734),
.A2(n_258),
.B1(n_254),
.B2(n_263),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_738),
.A2(n_347),
.B1(n_222),
.B2(n_277),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_861),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_840),
.B(n_472),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_862),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_858),
.B(n_640),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_738),
.A2(n_222),
.B1(n_220),
.B2(n_277),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_822),
.B(n_640),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_848),
.B(n_656),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_863),
.B(n_656),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_765),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_825),
.B(n_656),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_840),
.B(n_656),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_790),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_918),
.A2(n_796),
.B(n_857),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_900),
.B(n_790),
.Y(n_1046)
);

BUFx2_ASAP7_75t_SL g1047 ( 
.A(n_896),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_920),
.B(n_830),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_936),
.A2(n_842),
.B(n_820),
.C(n_811),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_969),
.A2(n_750),
.B(n_835),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_874),
.A2(n_859),
.B(n_661),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_SL g1052 ( 
.A1(n_975),
.A2(n_842),
.B(n_852),
.C(n_853),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_936),
.B(n_836),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_934),
.B(n_852),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_SL g1055 ( 
.A1(n_968),
.A2(n_364),
.B1(n_366),
.B2(n_369),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_911),
.B(n_837),
.Y(n_1056)
);

INVx3_ASAP7_75t_SL g1057 ( 
.A(n_910),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_990),
.A2(n_853),
.B1(n_846),
.B2(n_844),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_887),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_926),
.B(n_838),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_911),
.B(n_220),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_874),
.A2(n_656),
.B(n_661),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_944),
.B(n_342),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_916),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_924),
.A2(n_661),
.B(n_839),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_944),
.B(n_376),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_878),
.B(n_661),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1033),
.A2(n_342),
.B(n_343),
.C(n_347),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_979),
.B(n_343),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_912),
.B(n_354),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_916),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_971),
.A2(n_354),
.B1(n_382),
.B2(n_383),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_870),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_989),
.B(n_929),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_919),
.A2(n_661),
.B(n_850),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_971),
.B(n_625),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_65),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1035),
.B(n_625),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_889),
.A2(n_521),
.B(n_527),
.C(n_536),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1019),
.B(n_641),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1019),
.B(n_641),
.Y(n_1081)
);

AO32x2_ASAP7_75t_L g1082 ( 
.A1(n_930),
.A2(n_1),
.A3(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_902),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_949),
.B(n_645),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_929),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_884),
.B(n_383),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_871),
.B(n_73),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_884),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_869),
.B(n_645),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_947),
.A2(n_264),
.B(n_267),
.C(n_300),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_927),
.A2(n_697),
.B(n_682),
.C(n_678),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_913),
.A2(n_1015),
.B(n_1017),
.C(n_877),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_893),
.A2(n_302),
.B1(n_304),
.B2(n_328),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_902),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_933),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_893),
.A2(n_336),
.B1(n_380),
.B2(n_379),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_876),
.B(n_650),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_919),
.A2(n_522),
.B(n_519),
.Y(n_1098)
);

AO21x1_ASAP7_75t_L g1099 ( 
.A1(n_1041),
.A2(n_546),
.B(n_536),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_903),
.A2(n_338),
.B1(n_373),
.B2(n_368),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_980),
.B(n_377),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_913),
.B(n_678),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_904),
.B(n_660),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_980),
.B(n_502),
.Y(n_1104)
);

AO32x1_ASAP7_75t_L g1105 ( 
.A1(n_951),
.A2(n_546),
.A3(n_540),
.B1(n_542),
.B2(n_543),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1028),
.A2(n_522),
.B(n_507),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_939),
.B(n_660),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1015),
.A2(n_654),
.B(n_651),
.C(n_650),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_902),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1017),
.B(n_654),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_889),
.A2(n_542),
.B1(n_527),
.B2(n_543),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_L g1112 ( 
.A(n_953),
.B(n_79),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_885),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_883),
.A2(n_651),
.B(n_6),
.C(n_7),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_957),
.A2(n_562),
.B1(n_559),
.B2(n_557),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_980),
.B(n_519),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_SL g1117 ( 
.A1(n_991),
.A2(n_519),
.B(n_507),
.C(n_502),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_905),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_892),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_907),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_882),
.B(n_562),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_984),
.B(n_519),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1028),
.A2(n_522),
.B(n_519),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_899),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_965),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_991),
.A2(n_522),
.B(n_519),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_980),
.B(n_519),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_905),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_903),
.A2(n_507),
.B1(n_559),
.B2(n_557),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_935),
.B(n_559),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_974),
.A2(n_2),
.B(n_10),
.C(n_11),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_905),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_873),
.B(n_78),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_970),
.A2(n_13),
.B(n_14),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_935),
.B(n_559),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_906),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_917),
.B(n_559),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_923),
.B(n_559),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_901),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_965),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_SL g1141 ( 
.A1(n_957),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1036),
.A2(n_557),
.B(n_81),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_886),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_906),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_956),
.A2(n_82),
.B(n_173),
.C(n_153),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_941),
.B(n_557),
.Y(n_1146)
);

CKINVDCx16_ASAP7_75t_R g1147 ( 
.A(n_965),
.Y(n_1147)
);

BUFx4f_ASAP7_75t_L g1148 ( 
.A(n_937),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_1012),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1000),
.A2(n_557),
.B(n_19),
.C(n_22),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_897),
.A2(n_143),
.B(n_142),
.C(n_137),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_977),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_937),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_932),
.B(n_557),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_964),
.A2(n_135),
.B1(n_134),
.B2(n_131),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_988),
.A2(n_17),
.B(n_23),
.C(n_25),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_880),
.B(n_960),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_937),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_987),
.B(n_17),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_973),
.B(n_26),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_880),
.B(n_31),
.Y(n_1161)
);

OAI22x1_ASAP7_75t_L g1162 ( 
.A1(n_954),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_964),
.B(n_38),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1038),
.A2(n_84),
.B(n_127),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_990),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_SL g1166 ( 
.A1(n_915),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_961),
.A2(n_85),
.B(n_97),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_908),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_940),
.B(n_47),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_976),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_940),
.B(n_50),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_891),
.B(n_52),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1038),
.A2(n_87),
.B(n_90),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_982),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_953),
.B(n_95),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_995),
.B(n_52),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_SL g1177 ( 
.A1(n_915),
.A2(n_56),
.B1(n_129),
.B2(n_875),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_940),
.A2(n_56),
.B1(n_938),
.B2(n_875),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_973),
.B(n_938),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_982),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_962),
.A2(n_966),
.B(n_1040),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_982),
.B(n_940),
.Y(n_1182)
);

AO22x1_ASAP7_75t_L g1183 ( 
.A1(n_928),
.A2(n_1011),
.B1(n_986),
.B2(n_1003),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_879),
.B(n_895),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_982),
.B(n_1010),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_942),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_872),
.B(n_967),
.C(n_976),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_928),
.B(n_886),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_888),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_948),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1053),
.B(n_888),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1048),
.B(n_1034),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1182),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1075),
.A2(n_1039),
.B(n_943),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1050),
.A2(n_1123),
.B(n_1106),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1157),
.A2(n_967),
.B(n_996),
.C(n_872),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_L g1197 ( 
.A(n_1086),
.B(n_996),
.C(n_931),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1099),
.A2(n_1001),
.A3(n_909),
.B(n_898),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1182),
.B(n_1007),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1092),
.A2(n_955),
.B(n_997),
.C(n_922),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1108),
.A2(n_959),
.A3(n_981),
.B(n_1005),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1057),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1187),
.A2(n_955),
.B(n_1020),
.C(n_1013),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1177),
.A2(n_914),
.B1(n_952),
.B2(n_985),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1049),
.A2(n_1045),
.B(n_1065),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1178),
.A2(n_1008),
.A3(n_1009),
.B(n_992),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1177),
.A2(n_914),
.B1(n_952),
.B2(n_945),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1088),
.B(n_1030),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1120),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_SL g1210 ( 
.A1(n_1134),
.A2(n_1104),
.B(n_1116),
.C(n_1127),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1182),
.Y(n_1211)
);

OAI22x1_ASAP7_75t_L g1212 ( 
.A1(n_1161),
.A2(n_1021),
.B1(n_1039),
.B2(n_1030),
.Y(n_1212)
);

INVxp67_ASAP7_75t_SL g1213 ( 
.A(n_1064),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1110),
.A2(n_945),
.B(n_994),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1152),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1056),
.B(n_1004),
.Y(n_1216)
);

NOR2x1_ASAP7_75t_L g1217 ( 
.A(n_1074),
.B(n_999),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1122),
.A2(n_945),
.B(n_1042),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1185),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1179),
.B(n_972),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1166),
.A2(n_1029),
.B1(n_1010),
.B2(n_890),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1054),
.B(n_1018),
.Y(n_1222)
);

BUFx8_ASAP7_75t_SL g1223 ( 
.A(n_1059),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1076),
.A2(n_925),
.B(n_956),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1165),
.B(n_1014),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1071),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1090),
.A2(n_946),
.A3(n_1022),
.B(n_1023),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1168),
.Y(n_1228)
);

AO22x2_ASAP7_75t_L g1229 ( 
.A1(n_1166),
.A2(n_1037),
.B1(n_1032),
.B2(n_1006),
.Y(n_1229)
);

OA22x2_ASAP7_75t_L g1230 ( 
.A1(n_1055),
.A2(n_1031),
.B1(n_998),
.B2(n_1014),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1136),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1109),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1160),
.A2(n_1014),
.B1(n_1002),
.B2(n_1027),
.Y(n_1233)
);

AOI221x1_ASAP7_75t_L g1234 ( 
.A1(n_1170),
.A2(n_1024),
.B1(n_1016),
.B2(n_1044),
.C(n_1043),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1084),
.A2(n_894),
.B(n_921),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1151),
.A2(n_958),
.B(n_978),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1184),
.B(n_1026),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1115),
.A2(n_1029),
.B1(n_890),
.B2(n_1044),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1066),
.B(n_1025),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1080),
.B(n_1081),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1185),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1131),
.A2(n_983),
.B(n_963),
.C(n_1043),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1107),
.B(n_1002),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1115),
.A2(n_950),
.B1(n_1002),
.B2(n_1006),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1147),
.B(n_1046),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1114),
.A2(n_993),
.B(n_894),
.C(n_921),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1186),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1169),
.B(n_993),
.Y(n_1248)
);

NAND2x1_ASAP7_75t_L g1249 ( 
.A(n_1094),
.B(n_1189),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1154),
.A2(n_1102),
.B(n_1089),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1183),
.A2(n_1126),
.B(n_1138),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_SL g1252 ( 
.A(n_1144),
.B(n_1155),
.C(n_1069),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1125),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1159),
.C(n_1068),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1078),
.B(n_1163),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1109),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1098),
.A2(n_1167),
.B(n_1062),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1047),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1148),
.B(n_1094),
.Y(n_1259)
);

OA21x2_ASAP7_75t_L g1260 ( 
.A1(n_1142),
.A2(n_1146),
.B(n_1137),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1109),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1164),
.A2(n_1173),
.B(n_1129),
.Y(n_1262)
);

AOI21xp33_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1162),
.B(n_1072),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1052),
.A2(n_1185),
.B(n_1117),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1155),
.A2(n_1135),
.B(n_1130),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1150),
.A2(n_1156),
.A3(n_1105),
.B(n_1188),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1058),
.A2(n_1148),
.B(n_1097),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1103),
.A2(n_1143),
.B(n_1175),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1190),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1063),
.B(n_1061),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1087),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1077),
.B(n_1121),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1111),
.A2(n_1141),
.B(n_1091),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1095),
.Y(n_1274)
);

AOI221x1_ASAP7_75t_L g1275 ( 
.A1(n_1055),
.A2(n_1100),
.B1(n_1096),
.B2(n_1093),
.C(n_1087),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1101),
.A2(n_1112),
.B(n_1139),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1172),
.A2(n_1070),
.B(n_1077),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1111),
.A2(n_1112),
.B(n_1124),
.Y(n_1278)
);

AOI221x1_ASAP7_75t_L g1279 ( 
.A1(n_1105),
.A2(n_1082),
.B1(n_1158),
.B2(n_1153),
.C(n_1133),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1083),
.A2(n_1119),
.B(n_1113),
.Y(n_1280)
);

AO21x1_ASAP7_75t_L g1281 ( 
.A1(n_1189),
.A2(n_1082),
.B(n_1067),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1105),
.A2(n_1067),
.B(n_1145),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1060),
.B(n_1140),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1153),
.A2(n_1158),
.B(n_1180),
.Y(n_1284)
);

AND3x2_ASAP7_75t_L g1285 ( 
.A(n_1082),
.B(n_1149),
.C(n_1172),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1060),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1060),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1174),
.A2(n_1180),
.B(n_1153),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1158),
.A2(n_1174),
.B1(n_1180),
.B2(n_1132),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1149),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1174),
.B(n_1118),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1132),
.B(n_1118),
.Y(n_1292)
);

AO22x2_ASAP7_75t_L g1293 ( 
.A1(n_1118),
.A2(n_1178),
.B1(n_975),
.B2(n_1187),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1128),
.A2(n_1075),
.B(n_1050),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1128),
.A2(n_1092),
.B(n_918),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1087),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1181),
.A2(n_874),
.B(n_1092),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1088),
.B(n_766),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1053),
.B(n_936),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1064),
.Y(n_1300)
);

AOI31xp67_ASAP7_75t_L g1301 ( 
.A1(n_1110),
.A2(n_877),
.A3(n_927),
.B(n_1028),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1088),
.B(n_768),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_SL g1303 ( 
.A(n_1086),
.B(n_856),
.C(n_849),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1088),
.B(n_768),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1099),
.A2(n_1092),
.A3(n_764),
.B(n_1181),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1053),
.B(n_936),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1181),
.A2(n_1028),
.B(n_1051),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1088),
.B(n_766),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1177),
.B(n_1057),
.Y(n_1309)
);

AOI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1181),
.A2(n_1028),
.B(n_1051),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1057),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_SL g1312 ( 
.A(n_1125),
.B(n_829),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_R g1313 ( 
.A(n_1057),
.B(n_809),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1053),
.B(n_936),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1057),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1165),
.B(n_936),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1073),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1182),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1157),
.A2(n_936),
.B(n_918),
.C(n_1092),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1126),
.A2(n_1099),
.B(n_1181),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1117),
.A2(n_1092),
.B(n_1126),
.Y(n_1321)
);

NOR4xp25_ASAP7_75t_L g1322 ( 
.A(n_1161),
.B(n_918),
.C(n_1131),
.D(n_1170),
.Y(n_1322)
);

O2A1O1Ixp5_ASAP7_75t_L g1323 ( 
.A1(n_1122),
.A2(n_918),
.B(n_936),
.C(n_975),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1092),
.A2(n_918),
.B(n_1181),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1165),
.B(n_1085),
.Y(n_1325)
);

AO32x2_ASAP7_75t_L g1326 ( 
.A1(n_1177),
.A2(n_1178),
.A3(n_1166),
.B1(n_818),
.B2(n_930),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1232),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1319),
.A2(n_1323),
.B(n_1324),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1299),
.A2(n_1314),
.B(n_1306),
.C(n_1197),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1194),
.A2(n_1310),
.B(n_1307),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_SL g1331 ( 
.A(n_1322),
.B(n_1196),
.C(n_1309),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1316),
.B(n_1225),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1240),
.B(n_1192),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1204),
.A2(n_1207),
.B1(n_1221),
.B2(n_1229),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_SL g1335 ( 
.A(n_1202),
.B(n_1290),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1303),
.A2(n_1263),
.B(n_1252),
.C(n_1254),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1262),
.A2(n_1264),
.B(n_1268),
.Y(n_1337)
);

AND2x2_ASAP7_75t_SL g1338 ( 
.A(n_1309),
.B(n_1322),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1205),
.A2(n_1234),
.B(n_1236),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1267),
.B(n_1293),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1197),
.A2(n_1263),
.B(n_1207),
.C(n_1204),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1298),
.A2(n_1308),
.B(n_1255),
.C(n_1203),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1251),
.A2(n_1214),
.B(n_1282),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1280),
.A2(n_1224),
.B(n_1218),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1313),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1236),
.A2(n_1295),
.B(n_1250),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1221),
.A2(n_1229),
.B1(n_1233),
.B2(n_1277),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1295),
.Y(n_1348)
);

NOR2x1_ASAP7_75t_L g1349 ( 
.A(n_1217),
.B(n_1311),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1200),
.A2(n_1278),
.B(n_1250),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1210),
.A2(n_1244),
.B(n_1242),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1230),
.A2(n_1277),
.B1(n_1285),
.B2(n_1293),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1239),
.A2(n_1222),
.B1(n_1212),
.B2(n_1281),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1315),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1275),
.A2(n_1279),
.B1(n_1233),
.B2(n_1222),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1215),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1260),
.A2(n_1278),
.B(n_1244),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1260),
.A2(n_1273),
.B(n_1320),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1226),
.B(n_1300),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1302),
.B(n_1304),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1232),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1247),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1208),
.B(n_1272),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1265),
.A2(n_1220),
.B1(n_1248),
.B2(n_1216),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1273),
.A2(n_1246),
.B(n_1191),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1317),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1320),
.A2(n_1238),
.B(n_1286),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1238),
.A2(n_1289),
.B(n_1284),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1271),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1219),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1301),
.A2(n_1191),
.B(n_1243),
.Y(n_1371)
);

BUFx4f_ASAP7_75t_SL g1372 ( 
.A(n_1271),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1289),
.A2(n_1287),
.B(n_1241),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1199),
.B(n_1259),
.Y(n_1374)
);

AOI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1321),
.A2(n_1270),
.B(n_1237),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1253),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1223),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1228),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1258),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1206),
.B(n_1193),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1219),
.A2(n_1241),
.B(n_1288),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1231),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1269),
.A2(n_1305),
.B(n_1321),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1283),
.A2(n_1292),
.B(n_1318),
.C(n_1193),
.Y(n_1384)
);

OAI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1213),
.A2(n_1258),
.B1(n_1245),
.B2(n_1312),
.C(n_1274),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1211),
.A2(n_1318),
.B(n_1259),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1232),
.Y(n_1387)
);

AO22x2_ASAP7_75t_L g1388 ( 
.A1(n_1326),
.A2(n_1206),
.B1(n_1305),
.B2(n_1261),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1199),
.A2(n_1249),
.B(n_1305),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1199),
.A2(n_1201),
.B(n_1291),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1206),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1326),
.A2(n_1296),
.B1(n_1256),
.B2(n_1266),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1201),
.A2(n_1227),
.B(n_1198),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1296),
.B(n_1256),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1256),
.A2(n_1326),
.B1(n_1227),
.B2(n_1266),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1198),
.B(n_1266),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1201),
.A2(n_1227),
.B(n_1198),
.Y(n_1397)
);

NOR2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1252),
.B(n_1303),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1232),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1252),
.A2(n_1177),
.B1(n_1166),
.B2(n_936),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1252),
.A2(n_1177),
.B1(n_1166),
.B2(n_936),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1309),
.A2(n_1299),
.B1(n_1314),
.B2(n_1306),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1232),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1319),
.A2(n_936),
.B(n_918),
.C(n_1157),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1319),
.A2(n_918),
.B(n_936),
.C(n_1299),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1319),
.A2(n_936),
.B(n_918),
.C(n_1157),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1223),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1209),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1267),
.B(n_1293),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1199),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1279),
.A2(n_1099),
.A3(n_1281),
.B(n_1319),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1325),
.B(n_1199),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1311),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1209),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1299),
.A2(n_1314),
.B1(n_1306),
.B2(n_1177),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1252),
.A2(n_1177),
.B1(n_1166),
.B2(n_936),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1205),
.A2(n_1324),
.B(n_1297),
.Y(n_1422)
);

AOI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1299),
.A2(n_622),
.B1(n_936),
.B2(n_1314),
.C(n_1306),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1219),
.B(n_1241),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1325),
.B(n_1199),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1232),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1319),
.A2(n_936),
.B(n_918),
.C(n_1157),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1319),
.A2(n_1323),
.B(n_1092),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1311),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1219),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1319),
.A2(n_1323),
.B(n_1092),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1434)
);

AND2x2_ASAP7_75t_SL g1435 ( 
.A(n_1309),
.B(n_1322),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1313),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1313),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1311),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1319),
.B(n_768),
.C(n_936),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1209),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1209),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1309),
.A2(n_1299),
.B1(n_1314),
.B2(n_1306),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1195),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1406),
.A2(n_1428),
.B(n_1408),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1400),
.A2(n_1401),
.B1(n_1421),
.B2(n_1420),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1359),
.B(n_1347),
.Y(n_1449)
);

O2A1O1Ixp5_ASAP7_75t_L g1450 ( 
.A1(n_1351),
.A2(n_1420),
.B(n_1433),
.C(n_1429),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1380),
.A2(n_1396),
.B(n_1391),
.Y(n_1451)
);

O2A1O1Ixp5_ASAP7_75t_L g1452 ( 
.A1(n_1351),
.A2(n_1429),
.B(n_1433),
.C(n_1328),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1334),
.B(n_1331),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1376),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1430),
.Y(n_1456)
);

INVxp33_ASAP7_75t_L g1457 ( 
.A(n_1360),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1363),
.B(n_1415),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1380),
.A2(n_1396),
.B(n_1391),
.Y(n_1459)
);

AOI211xp5_ASAP7_75t_L g1460 ( 
.A1(n_1336),
.A2(n_1331),
.B(n_1445),
.C(n_1402),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1415),
.B(n_1426),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1400),
.A2(n_1421),
.B1(n_1401),
.B2(n_1352),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1382),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1407),
.A2(n_1336),
.B(n_1342),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1352),
.A2(n_1341),
.B1(n_1398),
.B2(n_1435),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1345),
.Y(n_1466)
);

INVx8_ASAP7_75t_L g1467 ( 
.A(n_1374),
.Y(n_1467)
);

NOR2xp67_ASAP7_75t_L g1468 ( 
.A(n_1437),
.B(n_1354),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1407),
.A2(n_1342),
.B(n_1439),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1416),
.B(n_1385),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1338),
.A2(n_1435),
.B1(n_1440),
.B2(n_1403),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1366),
.B(n_1356),
.Y(n_1472)
);

O2A1O1Ixp5_ASAP7_75t_L g1473 ( 
.A1(n_1328),
.A2(n_1350),
.B(n_1355),
.C(n_1343),
.Y(n_1473)
);

O2A1O1Ixp5_ASAP7_75t_L g1474 ( 
.A1(n_1350),
.A2(n_1355),
.B(n_1375),
.C(n_1402),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1338),
.A2(n_1434),
.B1(n_1418),
.B2(n_1403),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1417),
.A2(n_1440),
.B1(n_1434),
.B2(n_1418),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1417),
.A2(n_1423),
.B1(n_1385),
.B2(n_1445),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1438),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1423),
.A2(n_1374),
.B(n_1422),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1379),
.B(n_1378),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1364),
.A2(n_1353),
.B1(n_1349),
.B2(n_1412),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1357),
.A2(n_1358),
.B(n_1397),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1364),
.A2(n_1353),
.B1(n_1412),
.B2(n_1340),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1441),
.B(n_1442),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1370),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1340),
.A2(n_1412),
.B1(n_1372),
.B2(n_1369),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1367),
.Y(n_1488)
);

BUFx2_ASAP7_75t_R g1489 ( 
.A(n_1431),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1413),
.B(n_1386),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1377),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1340),
.A2(n_1372),
.B1(n_1369),
.B2(n_1392),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1362),
.Y(n_1493)
);

O2A1O1Ixp5_ASAP7_75t_L g1494 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1389),
.C(n_1390),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1393),
.A2(n_1330),
.B(n_1348),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1411),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1409),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1419),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1373),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1436),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1369),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1392),
.A2(n_1395),
.B1(n_1339),
.B2(n_1346),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1388),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1381),
.B(n_1327),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1383),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1337),
.A2(n_1344),
.B(n_1368),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1388),
.Y(n_1509)
);

O2A1O1Ixp5_ASAP7_75t_L g1510 ( 
.A1(n_1414),
.A2(n_1387),
.B(n_1361),
.C(n_1388),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1365),
.A2(n_1387),
.B(n_1361),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1365),
.A2(n_1427),
.B1(n_1399),
.B2(n_1404),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1414),
.B(n_1427),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1405),
.A2(n_1446),
.B(n_1425),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1384),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1384),
.B(n_1427),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1399),
.A2(n_1404),
.B(n_1335),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1414),
.B(n_1410),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1432),
.A2(n_1443),
.B(n_1444),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1351),
.A2(n_1357),
.B(n_1358),
.Y(n_1520)
);

INVx8_ASAP7_75t_L g1521 ( 
.A(n_1374),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1406),
.A2(n_1324),
.B(n_1297),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1377),
.Y(n_1523)
);

INVxp33_ASAP7_75t_SL g1524 ( 
.A(n_1335),
.Y(n_1524)
);

OAI31xp33_ASAP7_75t_L g1525 ( 
.A1(n_1398),
.A2(n_622),
.A3(n_1408),
.B(n_1406),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1406),
.A2(n_1319),
.B(n_1207),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_L g1528 ( 
.A(n_1345),
.B(n_1437),
.Y(n_1528)
);

AND2x4_ASAP7_75t_SL g1529 ( 
.A(n_1377),
.B(n_1271),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1377),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1406),
.A2(n_1324),
.B(n_1297),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1351),
.A2(n_1357),
.B(n_1358),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_R g1535 ( 
.A(n_1345),
.B(n_809),
.Y(n_1535)
);

INVxp33_ASAP7_75t_L g1536 ( 
.A(n_1332),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1400),
.A2(n_1421),
.B1(n_1401),
.B2(n_1420),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1406),
.A2(n_1319),
.B(n_1207),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1406),
.A2(n_1324),
.B(n_1297),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1500),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_R g1543 ( 
.A(n_1455),
.B(n_1535),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1504),
.B(n_1509),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1484),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1457),
.B(n_1536),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1449),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1475),
.B(n_1453),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1513),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1490),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1499),
.B(n_1488),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1527),
.B(n_1530),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1463),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1522),
.A2(n_1533),
.B(n_1539),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1479),
.B(n_1522),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1498),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1472),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1506),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1482),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1473),
.A2(n_1494),
.B(n_1474),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1482),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1473),
.A2(n_1494),
.B(n_1474),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1506),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1454),
.B(n_1458),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1488),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1452),
.B(n_1496),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1507),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1452),
.B(n_1496),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1514),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1515),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1483),
.B(n_1520),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1533),
.A2(n_1539),
.B(n_1447),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1510),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1480),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1510),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1450),
.A2(n_1532),
.B(n_1481),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1467),
.Y(n_1579)
);

AO21x2_ASAP7_75t_L g1580 ( 
.A1(n_1519),
.A2(n_1469),
.B(n_1464),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1490),
.B(n_1450),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1534),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1526),
.A2(n_1538),
.B(n_1511),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1512),
.A2(n_1487),
.B(n_1477),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1456),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1534),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1493),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1492),
.B(n_1495),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1555),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1575),
.B(n_1495),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1460),
.Y(n_1592)
);

NOR4xp25_ASAP7_75t_SL g1593 ( 
.A(n_1543),
.B(n_1497),
.C(n_1489),
.D(n_1525),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1581),
.B(n_1544),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1560),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1508),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1544),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1581),
.B(n_1508),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1577),
.B(n_1514),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1577),
.B(n_1465),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1542),
.A2(n_1448),
.B1(n_1537),
.B2(n_1462),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1568),
.B(n_1485),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1563),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1560),
.B(n_1516),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1570),
.B(n_1470),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1546),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1569),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1565),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1553),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1570),
.B(n_1486),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1551),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1540),
.B(n_1461),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1540),
.B(n_1478),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_L g1618 ( 
.A(n_1602),
.B(n_1574),
.C(n_1556),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1595),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1602),
.A2(n_1583),
.B1(n_1550),
.B2(n_1557),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1547),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1606),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1612),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1608),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1612),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1606),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1608),
.B(n_1552),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1589),
.B(n_1541),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1592),
.A2(n_1583),
.B1(n_1557),
.B2(n_1580),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1593),
.A2(n_1557),
.B1(n_1489),
.B2(n_1554),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1593),
.A2(n_1557),
.B1(n_1601),
.B2(n_1578),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1467),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1601),
.A2(n_1578),
.B1(n_1576),
.B2(n_1549),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1601),
.A2(n_1548),
.B1(n_1578),
.B2(n_1573),
.C(n_1549),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1610),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1594),
.B(n_1552),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1614),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1612),
.B(n_1545),
.Y(n_1641)
);

NOR2x2_ASAP7_75t_L g1642 ( 
.A(n_1611),
.B(n_1558),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1580),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1613),
.B(n_1578),
.C(n_1564),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1616),
.A2(n_1583),
.B1(n_1580),
.B2(n_1584),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1604),
.A2(n_1586),
.B(n_1582),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1589),
.A2(n_1585),
.B1(n_1521),
.B2(n_1579),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1590),
.B(n_1566),
.Y(n_1650)
);

AOI221x1_ASAP7_75t_L g1651 ( 
.A1(n_1609),
.A2(n_1572),
.B1(n_1517),
.B2(n_1567),
.C(n_1587),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1597),
.A2(n_1451),
.B(n_1459),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1618),
.A2(n_1524),
.B(n_1529),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

INVx4_ASAP7_75t_SL g1655 ( 
.A(n_1635),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1652),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_SL g1657 ( 
.A(n_1618),
.B(n_1588),
.C(n_1605),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1624),
.B(n_1628),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1640),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1645),
.A2(n_1607),
.B(n_1599),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1623),
.B(n_1615),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1644),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1640),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1620),
.B(n_1617),
.Y(n_1666)
);

OA21x2_ASAP7_75t_L g1667 ( 
.A1(n_1651),
.A2(n_1607),
.B(n_1596),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1642),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1619),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1620),
.B(n_1562),
.C(n_1564),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1619),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1629),
.B(n_1591),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1664),
.B(n_1629),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1669),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1664),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1659),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1668),
.B(n_1630),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1653),
.B(n_1466),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1659),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1675),
.B(n_1636),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1670),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1621),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1665),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1661),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1665),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1671),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1669),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1653),
.B(n_1631),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1671),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1655),
.B(n_1648),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1491),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_SL g1696 ( 
.A1(n_1658),
.A2(n_1637),
.B(n_1646),
.C(n_1632),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1654),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1656),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1656),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1671),
.B(n_1621),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1670),
.B(n_1649),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1661),
.B(n_1660),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1638),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.B(n_1622),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1660),
.B(n_1639),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_L g1707 ( 
.A(n_1666),
.B(n_1633),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1674),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1674),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1656),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1662),
.B(n_1648),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1662),
.B(n_1650),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1654),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1709),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1690),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1679),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1692),
.B(n_1663),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1696),
.B(n_1650),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1681),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1690),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1677),
.B(n_1675),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1655),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1523),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1693),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1710),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1676),
.B(n_1666),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1707),
.A2(n_1657),
.B1(n_1672),
.B2(n_1634),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1681),
.B(n_1655),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1681),
.B(n_1655),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1710),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1676),
.B(n_1705),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1677),
.B(n_1675),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1676),
.B(n_1641),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1680),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1531),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1698),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1686),
.B(n_1657),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1698),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1678),
.A2(n_1672),
.B1(n_1667),
.B2(n_1670),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1641),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1683),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1683),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1655),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1711),
.B(n_1625),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1655),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1697),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1687),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1684),
.B(n_1700),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1693),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1730),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1720),
.B(n_1711),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1720),
.B(n_1711),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1715),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1744),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1728),
.A2(n_1701),
.B1(n_1656),
.B2(n_1584),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1715),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1721),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1712),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1712),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1737),
.B(n_1688),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1732),
.B(n_1712),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1723),
.B(n_1705),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1730),
.B(n_1678),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1719),
.A2(n_1584),
.B1(n_1685),
.B2(n_1667),
.Y(n_1765)
);

AO21x1_ASAP7_75t_L g1766 ( 
.A1(n_1740),
.A2(n_1691),
.B(n_1702),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1718),
.A2(n_1727),
.B1(n_1729),
.B2(n_1691),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1726),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1723),
.B(n_1706),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1721),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1714),
.B(n_1726),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1725),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1731),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1750),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1724),
.B(n_1736),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1744),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1763),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1768),
.Y(n_1779)
);

AOI221x1_ASAP7_75t_L g1780 ( 
.A1(n_1768),
.A2(n_1739),
.B1(n_1737),
.B2(n_1731),
.C(n_1744),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1766),
.B(n_1730),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1729),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1755),
.B(n_1739),
.Y(n_1783)
);

O2A1O1Ixp5_ASAP7_75t_L g1784 ( 
.A1(n_1766),
.A2(n_1738),
.B(n_1746),
.C(n_1688),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_L g1785 ( 
.A(n_1767),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1756),
.B(n_1738),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1769),
.B(n_1746),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1776),
.B(n_1734),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1764),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1755),
.B(n_1749),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1765),
.A2(n_1699),
.B(n_1685),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1751),
.B(n_1685),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1777),
.B(n_1749),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1751),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1777),
.A2(n_1699),
.B1(n_1673),
.B2(n_1703),
.C(n_1702),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_L g1797 ( 
.A(n_1764),
.B(n_1688),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1761),
.A2(n_1772),
.B(n_1751),
.C(n_1764),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1778),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1795),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1795),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1782),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1788),
.B(n_1772),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1779),
.Y(n_1804)
);

NAND2x1_ASAP7_75t_L g1805 ( 
.A(n_1793),
.B(n_1751),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1791),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1787),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1790),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1789),
.B(n_1769),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1788),
.B(n_1764),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1803),
.A2(n_1781),
.B(n_1786),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1802),
.B(n_1783),
.Y(n_1812)
);

AOI221x1_ASAP7_75t_L g1813 ( 
.A1(n_1800),
.A2(n_1798),
.B1(n_1774),
.B2(n_1793),
.C(n_1792),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_SL g1814 ( 
.A(n_1803),
.B(n_1784),
.C(n_1785),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1805),
.A2(n_1786),
.B(n_1781),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1808),
.A2(n_1798),
.B1(n_1796),
.B2(n_1794),
.C(n_1774),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1807),
.A2(n_1760),
.B1(n_1793),
.B2(n_1752),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1810),
.B(n_1752),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1799),
.A2(n_1774),
.B(n_1771),
.C(n_1754),
.Y(n_1819)
);

OAI211xp5_ASAP7_75t_L g1820 ( 
.A1(n_1809),
.A2(n_1780),
.B(n_1761),
.C(n_1797),
.Y(n_1820)
);

AOI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1801),
.A2(n_1775),
.B(n_1773),
.C(n_1758),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1811),
.A2(n_1804),
.B(n_1806),
.C(n_1754),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1814),
.A2(n_1775),
.B1(n_1773),
.B2(n_1771),
.C(n_1757),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1815),
.A2(n_1813),
.B1(n_1817),
.B2(n_1816),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1812),
.A2(n_1753),
.B1(n_1684),
.B2(n_1762),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1818),
.B(n_1753),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1819),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1821),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1820),
.A2(n_1762),
.B1(n_1759),
.B2(n_1722),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1824),
.B(n_1759),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1826),
.B(n_1722),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1827),
.B(n_1757),
.Y(n_1832)
);

NAND2xp33_ASAP7_75t_SL g1833 ( 
.A(n_1829),
.B(n_1758),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1828),
.B(n_1770),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1825),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1822),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1830),
.B(n_1831),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1733),
.Y(n_1838)
);

AOI322xp5_ASAP7_75t_L g1839 ( 
.A1(n_1833),
.A2(n_1823),
.A3(n_1770),
.B1(n_1688),
.B2(n_1702),
.C1(n_1703),
.C2(n_1673),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1832),
.Y(n_1840)
);

XOR2x2_ASAP7_75t_L g1841 ( 
.A(n_1835),
.B(n_1834),
.Y(n_1841)
);

NAND2xp33_ASAP7_75t_R g1842 ( 
.A(n_1837),
.B(n_1673),
.Y(n_1842)
);

NAND5xp2_ASAP7_75t_L g1843 ( 
.A(n_1839),
.B(n_1717),
.C(n_1743),
.D(n_1742),
.E(n_1735),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1838),
.B(n_1748),
.Y(n_1844)
);

XOR2x2_ASAP7_75t_L g1845 ( 
.A(n_1844),
.B(n_1841),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1843),
.B1(n_1840),
.B2(n_1842),
.C(n_1747),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1846),
.Y(n_1847)
);

OAI21xp33_ASAP7_75t_L g1848 ( 
.A1(n_1846),
.A2(n_1747),
.B(n_1750),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

AND3x2_ASAP7_75t_L g1850 ( 
.A(n_1847),
.B(n_1528),
.C(n_1468),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1849),
.Y(n_1851)
);

OAI22x1_ASAP7_75t_L g1852 ( 
.A1(n_1850),
.A2(n_1733),
.B1(n_1697),
.B2(n_1713),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1851),
.A2(n_1713),
.B(n_1697),
.C(n_1708),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1852),
.B(n_1713),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1854),
.A2(n_1741),
.B(n_1745),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1855),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1708),
.B1(n_1689),
.B2(n_1687),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1689),
.B(n_1700),
.C(n_1704),
.Y(n_1858)
);


endmodule