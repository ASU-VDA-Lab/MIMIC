module fake_jpeg_15564_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_64),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_45),
.B(n_38),
.C(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_50),
.B1(n_43),
.B2(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_37),
.C(n_39),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_63),
.C(n_5),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_0),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_64),
.B(n_61),
.C(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_4),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_3),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_93),
.B(n_94),
.Y(n_98)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_72),
.B1(n_85),
.B2(n_90),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_73),
.C(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_87),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_103),
.B(n_105),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_94),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_104),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_72),
.C(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_88),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_99),
.B(n_19),
.C(n_21),
.D(n_22),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_16),
.C(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_110),
.B1(n_106),
.B2(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_26),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_27),
.C(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_34),
.Y(n_119)
);


endmodule