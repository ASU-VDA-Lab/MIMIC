module fake_jpeg_4389_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp33_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_39),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_40),
.B(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_16),
.B1(n_31),
.B2(n_12),
.Y(n_71)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_61),
.Y(n_84)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_51),
.B(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_59),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_14),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_2),
.B(n_4),
.Y(n_112)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_69),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_68),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_83),
.B1(n_98),
.B2(n_8),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_64),
.B1(n_44),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_82),
.B1(n_2),
.B2(n_4),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_103),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_29),
.C(n_18),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_74),
.C(n_98),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_91),
.B1(n_101),
.B2(n_109),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_88),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_87),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_5),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_57),
.B1(n_52),
.B2(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_23),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_100),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_1),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_122),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_65),
.B1(n_69),
.B2(n_100),
.Y(n_164)
);

OR2x4_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_5),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_117),
.A2(n_121),
.B(n_75),
.Y(n_178)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_137),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_6),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_82),
.B1(n_86),
.B2(n_81),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_71),
.B1(n_77),
.B2(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_131),
.B1(n_125),
.B2(n_133),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_147),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_86),
.B1(n_110),
.B2(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_81),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_156),
.B1(n_170),
.B2(n_116),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_157),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_159),
.Y(n_213)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_160),
.B(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_182),
.B1(n_140),
.B2(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_166),
.B(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_66),
.B1(n_97),
.B2(n_79),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_175),
.B1(n_180),
.B2(n_145),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_119),
.A2(n_75),
.B1(n_107),
.B2(n_97),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_181),
.B(n_129),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_130),
.A2(n_66),
.B(n_107),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_107),
.B1(n_142),
.B2(n_113),
.Y(n_182)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_205),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_156),
.C(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_171),
.C(n_107),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_190),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_189),
.A2(n_197),
.B1(n_208),
.B2(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_191),
.B(n_193),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_197),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_135),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_126),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_157),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_215),
.B(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_126),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_135),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_135),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_210),
.A2(n_216),
.B1(n_219),
.B2(n_159),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_137),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_137),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_198),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_127),
.Y(n_214)
);

NAND2x1p5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_118),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_229),
.B(n_231),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_246),
.B(n_218),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_232),
.C(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_150),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_118),
.B1(n_165),
.B2(n_143),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_129),
.B(n_154),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_209),
.B1(n_214),
.B2(n_201),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_240),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_160),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_244),
.C(n_215),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_115),
.B1(n_134),
.B2(n_183),
.C(n_177),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_213),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_115),
.C(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_189),
.A2(n_149),
.B1(n_162),
.B2(n_205),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_149),
.Y(n_267)
);

AO22x2_ASAP7_75t_SL g246 ( 
.A1(n_199),
.A2(n_149),
.B1(n_162),
.B2(n_185),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_253),
.B1(n_267),
.B2(n_237),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_223),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_218),
.B1(n_214),
.B2(n_187),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_261),
.C(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_221),
.B(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_191),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_225),
.B(n_199),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_266),
.B(n_231),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_194),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_217),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_265),
.C(n_261),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_190),
.C(n_216),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_233),
.B(n_204),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_246),
.B1(n_235),
.B2(n_229),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_272),
.A2(n_278),
.B(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_256),
.A2(n_234),
.B1(n_268),
.B2(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_259),
.B1(n_245),
.B2(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_247),
.C(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_289),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_256),
.B1(n_279),
.B2(n_299),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_260),
.B1(n_266),
.B2(n_220),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_260),
.B(n_252),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_296),
.C(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_273),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_247),
.C(n_263),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_297),
.A2(n_249),
.B1(n_200),
.B2(n_280),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_248),
.B1(n_276),
.B2(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_270),
.B1(n_274),
.B2(n_266),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_264),
.C(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_305),
.C(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_309),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_275),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_260),
.B1(n_243),
.B2(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_292),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_282),
.B(n_228),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_308),
.C(n_305),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_287),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_298),
.B(n_290),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_223),
.Y(n_326)
);

NAND4xp25_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_289),
.C(n_298),
.D(n_202),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_244),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_303),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_326),
.B(n_327),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_325),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_315),
.B(n_320),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_324),
.Y(n_333)
);

AOI31xp67_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_326),
.A3(n_323),
.B(n_314),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);

AOI221xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_330),
.B1(n_317),
.B2(n_308),
.C(n_302),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_300),
.Y(n_336)
);


endmodule