module fake_jpeg_3654_n_84 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_21),
.C(n_19),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_26),
.B(n_28),
.C(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_33),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_23),
.B1(n_31),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_37),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_27),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_53),
.B(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_10),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_13),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_61),
.B1(n_6),
.B2(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_48),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_5),
.B(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_67),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_49),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_46),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_71),
.C(n_7),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_14),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_15),
.B(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_68),
.C(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_76),
.B1(n_66),
.B2(n_74),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_63),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_71),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_78),
.C(n_73),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_8),
.Y(n_84)
);


endmodule