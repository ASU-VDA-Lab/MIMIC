module fake_jpeg_20905_n_85 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_SL g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_19),
.B1(n_18),
.B2(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_10),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_12),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_40),
.B(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_27),
.C(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_27),
.B1(n_8),
.B2(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_27),
.B2(n_8),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_27),
.B(n_23),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_59),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_0),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_53),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_66),
.C(n_57),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_67),
.C(n_1),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_55),
.A3(n_11),
.B1(n_13),
.B2(n_6),
.C(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_13),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_0),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_80),
.B1(n_67),
.B2(n_3),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_2),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_2),
.Y(n_85)
);


endmodule