module fake_jpeg_10011_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_38),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_20),
.C(n_31),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_39),
.B1(n_38),
.B2(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_20),
.C(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_71),
.B1(n_78),
.B2(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_64),
.Y(n_95)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_41),
.B1(n_17),
.B2(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_41),
.B1(n_17),
.B2(n_18),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_35),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_55),
.C(n_40),
.Y(n_105)
);

NOR4xp25_ASAP7_75t_SL g80 ( 
.A(n_42),
.B(n_58),
.C(n_35),
.D(n_3),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_25),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_1),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_28),
.C(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_24),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g99 ( 
.A(n_88),
.Y(n_99)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_34),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_21),
.B1(n_19),
.B2(n_33),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_21),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_112),
.B(n_76),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_110),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_107),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_109),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_65),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_52),
.C(n_40),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_40),
.B1(n_28),
.B2(n_3),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_21),
.B(n_19),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_67),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_94),
.B1(n_89),
.B2(n_60),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_59),
.B1(n_69),
.B2(n_63),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_133),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_21),
.Y(n_170)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_80),
.B1(n_75),
.B2(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_112),
.B1(n_105),
.B2(n_104),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_74),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_90),
.C(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_87),
.B(n_72),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_114),
.B(n_33),
.Y(n_167)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_72),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_90),
.B(n_81),
.C(n_63),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_104),
.B1(n_66),
.B2(n_64),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_149),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_68),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_147),
.B1(n_126),
.B2(n_132),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_99),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_163),
.C(n_176),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_160),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_114),
.C(n_92),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_59),
.B1(n_97),
.B2(n_116),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_97),
.B1(n_120),
.B2(n_122),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_173),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_148),
.B(n_138),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_133),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_127),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_62),
.C(n_110),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_178),
.C(n_136),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_33),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_187),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_190),
.C(n_191),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_148),
.B(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_131),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_123),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_143),
.B1(n_172),
.B2(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_146),
.C(n_143),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_200),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_126),
.B1(n_19),
.B2(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_160),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_1),
.B(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_168),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_144),
.C(n_110),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_177),
.C(n_180),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_62),
.B1(n_33),
.B2(n_5),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_219),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_217),
.C(n_184),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_153),
.B1(n_189),
.B2(n_195),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_222),
.B1(n_199),
.B2(n_200),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_171),
.C(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_223),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_187),
.B(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_183),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_235),
.C(n_236),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_154),
.C(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_229),
.B(n_234),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_215),
.B1(n_62),
.B2(n_110),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_212),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_168),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_184),
.C(n_191),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_217),
.C(n_213),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_239),
.C(n_14),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_169),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_241),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_249),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_15),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_236),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_13),
.B1(n_3),
.B2(n_5),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_230),
.B1(n_228),
.B2(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_231),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_247),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_241),
.C(n_248),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_2),
.C(n_7),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_2),
.B(n_8),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_265),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_243),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_254),
.B(n_259),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_240),
.B(n_9),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_271),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_263),
.C(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_274),
.A2(n_275),
.B(n_276),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_10),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_11),
.B(n_12),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_277),
.B1(n_11),
.B2(n_12),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_12),
.Y(n_281)
);


endmodule