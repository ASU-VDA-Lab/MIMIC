module real_jpeg_31286_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_556;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_1),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_1),
.A2(n_346),
.B1(n_471),
.B2(n_473),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_1),
.A2(n_346),
.B1(n_525),
.B2(n_527),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_2),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_2),
.A2(n_159),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_2),
.A2(n_159),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_2),
.A2(n_159),
.B1(n_334),
.B2(n_500),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_3),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_4),
.A2(n_198),
.B1(n_203),
.B2(n_204),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_4),
.A2(n_203),
.B1(n_380),
.B2(n_382),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_4),
.A2(n_203),
.B1(n_455),
.B2(n_458),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_4),
.A2(n_203),
.B1(n_446),
.B2(n_543),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

INVx2_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_5),
.A2(n_72),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_5),
.A2(n_72),
.B1(n_277),
.B2(n_281),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g425 ( 
.A1(n_5),
.A2(n_72),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_5),
.A2(n_72),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_6),
.A2(n_33),
.B1(n_37),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_41),
.B1(n_118),
.B2(n_124),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_6),
.A2(n_41),
.B1(n_248),
.B2(n_252),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_6),
.A2(n_41),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_7),
.A2(n_101),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_143),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_7),
.A2(n_143),
.B1(n_389),
.B2(n_391),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_7),
.A2(n_143),
.B1(n_444),
.B2(n_446),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_8),
.A2(n_410),
.B1(n_412),
.B2(n_415),
.Y(n_409)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_8),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_8),
.A2(n_382),
.B1(n_415),
.B2(n_492),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_8),
.A2(n_415),
.B1(n_577),
.B2(n_579),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_9),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_9),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_9),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_10),
.Y(n_184)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_12),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_12),
.A2(n_289),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_12),
.A2(n_289),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g566 ( 
.A1(n_12),
.A2(n_289),
.B1(n_543),
.B2(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g464 ( 
.A1(n_14),
.A2(n_412),
.B1(n_465),
.B2(n_468),
.Y(n_464)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_14),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_14),
.A2(n_215),
.B1(n_468),
.B2(n_533),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_588),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_15),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_16),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_17),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_18),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_19),
.A2(n_32),
.B1(n_42),
.B2(n_47),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_19),
.B(n_174),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_19),
.A2(n_207),
.A3(n_209),
.B1(n_214),
.B2(n_219),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_19),
.A2(n_55),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_19),
.B(n_334),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_19),
.A2(n_333),
.B(n_357),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_556),
.B2(n_587),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_395),
.B(n_551),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_308),
.B(n_394),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_257),
.B(n_307),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_186),
.B(n_256),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_149),
.Y(n_27)
);

AOI21x1_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_85),
.B(n_146),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_62),
.B(n_84),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_53),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_32),
.A2(n_47),
.B1(n_64),
.B2(n_73),
.Y(n_63)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_36),
.Y(n_345)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_36),
.Y(n_414)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_36),
.Y(n_467)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_42),
.A2(n_47),
.B1(n_409),
.B2(n_463),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_46),
.Y(n_153)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_46),
.Y(n_419)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_47),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_47),
.A2(n_141),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_47),
.A2(n_342),
.B1(n_409),
.B2(n_416),
.Y(n_408)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_47),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_50),
.Y(n_196)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_50),
.Y(n_340)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_52),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_97),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_55),
.A2(n_96),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_55),
.B(n_215),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_R g293 ( 
.A(n_55),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_58),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_75),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_68),
.Y(n_291)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_76),
.A2(n_134),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_76),
.A2(n_134),
.B1(n_264),
.B2(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_76),
.A2(n_134),
.B1(n_379),
.B2(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_76),
.A2(n_134),
.B1(n_403),
.B2(n_470),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_76),
.A2(n_134),
.B1(n_470),
.B2(n_491),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g572 ( 
.A1(n_76),
.A2(n_134),
.B(n_532),
.Y(n_572)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AO21x2_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_106),
.B(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_139),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_114),
.B1(n_115),
.B2(n_138),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_87),
.B(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B1(n_100),
.B2(n_105),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_110),
.Y(n_386)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_138),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_129),
.B2(n_133),
.Y(n_115)
);

NAND2x1_ASAP7_75t_SL g165 ( 
.A(n_116),
.B(n_166),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g228 ( 
.A1(n_116),
.A2(n_133),
.B1(n_166),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_116),
.A2(n_133),
.B1(n_531),
.B2(n_536),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_133),
.Y(n_164)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_128),
.Y(n_268)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_155),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_144),
.A2(n_197),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_144),
.A2(n_288),
.B1(n_338),
.B2(n_341),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_163),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_173),
.C(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B(n_173),
.C(n_185),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.C(n_173),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_R g190 ( 
.A(n_164),
.B(n_165),
.Y(n_190)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_169),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_172),
.Y(n_407)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

AOI22x1_ASAP7_75t_L g503 ( 
.A1(n_174),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_174),
.A2(n_504),
.B1(n_506),
.B2(n_524),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AO21x2_ASAP7_75t_L g234 ( 
.A1(n_175),
.A2(n_219),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_182),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_176),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_176),
.Y(n_493)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2x1_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_189),
.B(n_191),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_226),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_192),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_206),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_193),
.B(n_206),
.Y(n_261)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_211),
.Y(n_245)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_212),
.Y(n_434)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_221),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_228),
.B(n_232),
.C(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_234),
.A2(n_246),
.B1(n_247),
.B2(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_234),
.A2(n_246),
.B1(n_276),
.B2(n_388),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g432 ( 
.A1(n_234),
.A2(n_246),
.B1(n_388),
.B2(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_234),
.A2(n_246),
.B1(n_433),
.B2(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_234),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_234),
.A2(n_246),
.B1(n_575),
.B2(n_576),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_236),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_248),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_250),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_255),
.Y(n_511)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_255),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_305),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_273),
.B2(n_274),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_271),
.B2(n_272),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_262),
.B(n_272),
.C(n_273),
.Y(n_393)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_268),
.Y(n_475)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_268),
.Y(n_535)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_293),
.C(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_280),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

BUFx4f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_356),
.B1(n_360),
.B2(n_371),
.Y(n_355)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_294),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_294),
.A2(n_360),
.B1(n_443),
.B2(n_450),
.Y(n_442)
);

OAI22x1_ASAP7_75t_SL g497 ( 
.A1(n_294),
.A2(n_360),
.B1(n_443),
.B2(n_498),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_300),
.Y(n_526)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_301),
.Y(n_578)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_301),
.Y(n_580)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_393),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_393),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_353),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_351),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_311),
.B(n_351),
.C(n_353),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_337),
.B1(n_349),
.B2(n_350),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_312),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_312),
.B(n_350),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_312),
.B(n_350),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.A3(n_318),
.B1(n_325),
.B2(n_332),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_323),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_345),
.Y(n_348)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_377),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_SL g400 ( 
.A(n_355),
.B(n_378),
.C(n_387),
.Y(n_400)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_361),
.A2(n_424),
.B1(n_425),
.B2(n_431),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_361),
.A2(n_424),
.B1(n_499),
.B2(n_542),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_361),
.A2(n_424),
.B1(n_542),
.B2(n_566),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_366),
.B2(n_368),
.Y(n_362)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_363),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_370),
.Y(n_373)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_370),
.Y(n_545)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_376),
.Y(n_449)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_376),
.Y(n_502)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_376),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND4xp25_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_436),
.C(n_514),
.D(n_546),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_397),
.B(n_398),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_420),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_400),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_401),
.B(n_420),
.C(n_548),
.Y(n_547)
);

XOR2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_408),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_408),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_432),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_432),
.C(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

A2O1A1O1Ixp25_ASAP7_75t_L g551 ( 
.A1(n_436),
.A2(n_514),
.B(n_552),
.C(n_554),
.D(n_555),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_476),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_437),
.B(n_476),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_459),
.C(n_461),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_439),
.B(n_461),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_478),
.C(n_480),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_453),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_453),
.Y(n_480)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_454),
.Y(n_505)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_459),
.B(n_550),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_469),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_485),
.B(n_487),
.Y(n_484)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

BUFx4f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_481),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_482),
.C(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_494),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_484),
.B1(n_488),
.B2(n_489),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_484),
.B(n_490),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_484),
.A2(n_541),
.B(n_583),
.Y(n_582)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_495),
.A2(n_496),
.B1(n_512),
.B2(n_513),
.Y(n_494)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_495),
.Y(n_513)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_503),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_497),
.Y(n_520)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_503),
.Y(n_519)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_519),
.C(n_520),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_517),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_517),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_518),
.B(n_560),
.C(n_561),
.Y(n_559)
);

XOR2x1_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_538),
.Y(n_521)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_522),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_530),
.B(n_537),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_530),
.Y(n_537)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_524),
.Y(n_575)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_535),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_538),
.Y(n_560)
);

XNOR2x1_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_539),
.Y(n_583)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_547),
.B(n_549),
.C(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_556),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_585),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_562),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_562),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_581),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_570),
.Y(n_564)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_571),
.A2(n_572),
.B1(n_573),
.B2(n_574),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_584),
.Y(n_581)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_591),
.Y(n_588)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);


endmodule