module fake_netlist_1_8799_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
BUFx4f_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
OR2x6_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_4), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
OAI33xp33_ASAP7_75t_L g11 ( .A1(n_8), .A2(n_7), .A3(n_4), .B1(n_3), .B2(n_2), .B3(n_1), .Y(n_11) );
AOI221xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_4), .B1(n_3), .B2(n_7), .C(n_0), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_13), .B(n_10), .Y(n_14) );
AOI222xp33_ASAP7_75t_SL g15 ( .A1(n_14), .A2(n_1), .B1(n_3), .B2(n_12), .C1(n_5), .C2(n_6), .Y(n_15) );
endmodule