module fake_jpeg_31711_n_90 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_90);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_90;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_24),
.Y(n_40)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_13),
.B(n_19),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_30),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_15),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_31),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_17),
.B1(n_11),
.B2(n_21),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_17),
.B1(n_11),
.B2(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_10),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_50),
.B1(n_52),
.B2(n_46),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

AO221x1_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_71),
.B1(n_60),
.B2(n_56),
.C(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_74),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_57),
.C(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_76),
.B1(n_75),
.B2(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_79),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_36),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_82),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_6),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_6),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B(n_9),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_53),
.B(n_0),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);


endmodule