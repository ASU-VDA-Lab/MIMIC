module fake_aes_4591_n_30 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_3), .B(n_4), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
NAND3xp33_ASAP7_75t_SL g15 ( .A(n_10), .B(n_0), .C(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_5), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_11), .Y(n_17) );
AOI22xp33_ASAP7_75t_SL g18 ( .A1(n_16), .A2(n_12), .B1(n_13), .B2(n_8), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_19), .B(n_12), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_15), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx2_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_22), .B(n_12), .Y(n_25) );
AOI32xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_6), .A3(n_7), .B1(n_24), .B2(n_19), .Y(n_26) );
INVx4_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
endmodule