module real_jpeg_3361_n_16 (n_5, n_4, n_8, n_0, n_12, n_319, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_319;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_1),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_1),
.B(n_41),
.C(n_44),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_136),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_1),
.B(n_103),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_1),
.B(n_39),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_31),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_1),
.A2(n_31),
.B(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_87),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_1),
.A2(n_25),
.B(n_251),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_4),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_145),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_41),
.B1(n_45),
.B2(n_145),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_145),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_5),
.A2(n_25),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_36),
.B1(n_41),
.B2(n_45),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_5),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_116),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_6),
.A2(n_41),
.B1(n_45),
.B2(n_116),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_116),
.Y(n_236)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_66),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_11),
.A2(n_41),
.B1(n_45),
.B2(n_66),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_12),
.A2(n_41),
.B1(n_45),
.B2(n_53),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_12),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_13),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_13),
.A2(n_41),
.B1(n_45),
.B2(n_118),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_118),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_91),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_38),
.C(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_22)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_23),
.A2(n_35),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_23),
.A2(n_29),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_23),
.A2(n_29),
.B1(n_115),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_23),
.A2(n_117),
.B(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_23),
.A2(n_29),
.B1(n_144),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_23),
.A2(n_86),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_26),
.A2(n_30),
.B(n_135),
.C(n_137),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_27),
.B(n_136),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_27),
.B(n_28),
.C(n_31),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_29),
.A2(n_33),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_31),
.B1(n_61),
.B2(n_62),
.Y(n_69)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_31),
.A2(n_49),
.A3(n_62),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_71),
.C(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_38),
.A2(n_70),
.B1(n_76),
.B2(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_46),
.B(n_51),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_39),
.B(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_39),
.A2(n_46),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_39),
.A2(n_46),
.B1(n_179),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_40),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_40),
.A2(n_109),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_40),
.A2(n_129),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_40),
.B(n_52),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_41),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_41),
.B(n_192),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_46),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_46),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OA22x2_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_48),
.B(n_61),
.Y(n_215)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_49),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_52),
.A2(n_129),
.B(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_56),
.A2(n_68),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_60),
.B(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_68),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_59),
.A2(n_67),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_59),
.A2(n_67),
.B1(n_77),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_64),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_60),
.B(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_60),
.A2(n_68),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_60),
.A2(n_68),
.B1(n_142),
.B2(n_236),
.Y(n_252)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_71),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_71),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_75),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_76),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_87),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_299),
.B(n_313),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_279),
.B(n_298),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_167),
.B(n_278),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_146),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_95),
.B(n_146),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_120),
.C(n_131),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_96),
.B(n_120),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_112),
.B2(n_113),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_114),
.C(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_99),
.B(n_108),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_106),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_100),
.A2(n_102),
.B(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_100),
.A2(n_102),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_100),
.A2(n_106),
.B(n_124),
.Y(n_216)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_101),
.A2(n_123),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_101),
.A2(n_103),
.B1(n_136),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_101),
.A2(n_103),
.B1(n_194),
.B2(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_102),
.A2(n_126),
.B(n_140),
.Y(n_241)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_130),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_131),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.C(n_143),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_132),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_133),
.A2(n_134),
.B1(n_138),
.B2(n_258),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_138),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_141),
.B(n_143),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_166),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_150),
.B(n_156),
.C(n_166),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_151),
.A2(n_152),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_152),
.B(n_153),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_152),
.A2(n_287),
.B(n_290),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_159),
.B(n_162),
.C(n_165),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_163),
.Y(n_295)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI321xp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_260),
.A3(n_270),
.B1(n_276),
.B2(n_277),
.C(n_319),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_244),
.B(n_259),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_225),
.B(n_243),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_207),
.B(n_224),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_188),
.B(n_206),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_181),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_181),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_178),
.C(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_200),
.B(n_205),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_195),
.B(n_199),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_204),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_217),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_218),
.C(n_221),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_242),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_242),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_231),
.C(n_232),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_256),
.C(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_248),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.CI(n_253),
.CON(n_248),
.SN(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_263),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_269),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_297),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_297),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_285),
.C(n_291),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_294),
.B(n_296),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_305),
.C(n_309),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_305),
.CI(n_309),
.CON(n_312),
.SN(n_312)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_310),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_312),
.Y(n_317)
);


endmodule