module fake_ariane_2019_n_1084 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_255, n_122, n_257, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1084);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_257;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1084;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_398;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_611;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_851;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_106),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_46),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_112),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_31),
.Y(n_265)
);

BUFx8_ASAP7_75t_SL g266 ( 
.A(n_156),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_120),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_24),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_95),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_204),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_5),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_192),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_69),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_202),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_222),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_99),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_68),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_206),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_127),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_260),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_129),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_0),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_108),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_116),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_113),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_180),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_28),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_1),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_118),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_173),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_10),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_35),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_103),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_196),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_60),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_94),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_28),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_125),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_157),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_181),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_133),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_179),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_115),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_88),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_195),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_52),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_264),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_266),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_299),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_266),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_265),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_291),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_270),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_291),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_291),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_262),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_312),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_298),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_0),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_261),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_263),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_265),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_265),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_271),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_272),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_269),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_273),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_275),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_279),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g369 ( 
.A1(n_359),
.A2(n_315),
.B(n_301),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_320),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_326),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_331),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_364),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_322),
.C(n_289),
.Y(n_384)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_277),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_352),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_334),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_333),
.B(n_289),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_361),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_361),
.B(n_280),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_325),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_346),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_405),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_410),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_349),
.Y(n_419)
);

OR2x6_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_355),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_392),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_351),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_385),
.A2(n_343),
.B1(n_335),
.B2(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_274),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_405),
.B(n_394),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_297),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_386),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_307),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_405),
.B(n_324),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_411),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_410),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_321),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_411),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_281),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_283),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_385),
.A2(n_322),
.B1(n_320),
.B2(n_323),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_320),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_320),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_369),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_284),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_1),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_404),
.B(n_285),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_286),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_408),
.B(n_287),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_390),
.B(n_2),
.Y(n_470)
);

BUFx4f_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_292),
.Y(n_472)
);

BUFx8_ASAP7_75t_SL g473 ( 
.A(n_398),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_414),
.B(n_293),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_408),
.B(n_295),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_318),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_406),
.B(n_303),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_416),
.B(n_308),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_309),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_430),
.B(n_400),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_409),
.B1(n_407),
.B2(n_403),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_438),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_430),
.B(n_436),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_413),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_372),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_479),
.B(n_385),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_369),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_428),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_438),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_374),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_374),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_432),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_376),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_376),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_377),
.Y(n_504)
);

OAI221xp5_ASAP7_75t_L g505 ( 
.A1(n_453),
.A2(n_377),
.B1(n_370),
.B2(n_313),
.C(n_314),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_398),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_436),
.B(n_310),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_311),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_445),
.B(n_316),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_3),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_447),
.B(n_3),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_435),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_429),
.B(n_4),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_431),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_450),
.B(n_6),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

NAND2x1_ASAP7_75t_L g519 ( 
.A(n_417),
.B(n_454),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_7),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_419),
.B(n_7),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_476),
.B(n_8),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_471),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_427),
.B(n_9),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_473),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_457),
.B(n_11),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_418),
.B(n_11),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_447),
.B(n_12),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_423),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_423),
.B(n_12),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_424),
.B(n_13),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_424),
.B(n_13),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_14),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_449),
.B(n_14),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_472),
.B(n_15),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_459),
.B(n_15),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_453),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_474),
.B(n_16),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_445),
.B(n_17),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_420),
.B(n_18),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_19),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_449),
.B(n_482),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_19),
.C(n_20),
.Y(n_552)
);

BUFx2_ASAP7_75t_SL g553 ( 
.A(n_459),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

A2O1A1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_544),
.A2(n_471),
.B(n_467),
.C(n_481),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_496),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_491),
.A2(n_481),
.B1(n_477),
.B2(n_460),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_491),
.B(n_477),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_500),
.A2(n_429),
.B1(n_417),
.B2(n_441),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_493),
.A2(n_508),
.B(n_489),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_520),
.B(n_451),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_504),
.B(n_498),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_489),
.A2(n_462),
.B(n_452),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_544),
.A2(n_455),
.B(n_464),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_523),
.A2(n_480),
.B(n_439),
.C(n_458),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_502),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_503),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_506),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_534),
.A2(n_439),
.B(n_461),
.C(n_456),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_542),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_490),
.B(n_420),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_SL g578 ( 
.A1(n_510),
.A2(n_456),
.B(n_461),
.C(n_417),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_535),
.A2(n_439),
.B(n_426),
.C(n_460),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_488),
.A2(n_439),
.B(n_460),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_498),
.B(n_420),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_497),
.A2(n_41),
.B(n_40),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_540),
.B(n_426),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_492),
.B(n_473),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_519),
.A2(n_43),
.B(n_42),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_21),
.Y(n_586)
);

INVx6_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

O2A1O1Ixp5_ASAP7_75t_L g588 ( 
.A1(n_521),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_530),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_532),
.B(n_22),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_539),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_591)
);

INVx11_ASAP7_75t_L g592 ( 
.A(n_528),
.Y(n_592)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_526),
.A2(n_45),
.B(n_44),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_513),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_507),
.A2(n_48),
.B(n_47),
.Y(n_595)
);

OAI321xp33_ASAP7_75t_L g596 ( 
.A1(n_543),
.A2(n_26),
.A3(n_27),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_485),
.A2(n_50),
.B(n_49),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_521),
.B(n_484),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g599 ( 
.A(n_486),
.B(n_51),
.Y(n_599)
);

O2A1O1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_512),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_507),
.A2(n_54),
.B(n_53),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_483),
.A2(n_516),
.B(n_514),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_518),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_483),
.A2(n_56),
.B(n_55),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_522),
.A2(n_59),
.B(n_58),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_542),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_543),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_527),
.A2(n_62),
.B(n_61),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_485),
.A2(n_64),
.B(n_63),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_32),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_533),
.B(n_33),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_515),
.A2(n_66),
.B(n_65),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_517),
.A2(n_71),
.B(n_70),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_537),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_495),
.B(n_34),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_561),
.B(n_545),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_598),
.A2(n_552),
.B(n_505),
.C(n_538),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_566),
.B(n_547),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_567),
.A2(n_531),
.B(n_511),
.Y(n_621)
);

OAI22x1_ASAP7_75t_L g622 ( 
.A1(n_583),
.A2(n_550),
.B1(n_511),
.B2(n_531),
.Y(n_622)
);

INVx3_ASAP7_75t_SL g623 ( 
.A(n_573),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_563),
.A2(n_546),
.B(n_542),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_558),
.A2(n_552),
.B(n_541),
.C(n_524),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_577),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_554),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_564),
.A2(n_560),
.B(n_562),
.Y(n_628)
);

OAI21x1_ASAP7_75t_SL g629 ( 
.A1(n_602),
.A2(n_529),
.B(n_541),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_597),
.A2(n_546),
.B(n_542),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_557),
.A2(n_548),
.B(n_546),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_568),
.A2(n_512),
.B1(n_553),
.B2(n_546),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_576),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_587),
.B(n_548),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_581),
.B(n_548),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

AOI21x1_ASAP7_75t_SL g638 ( 
.A1(n_586),
.A2(n_548),
.B(n_35),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_571),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_580),
.A2(n_73),
.B(n_72),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_574),
.B(n_36),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_593),
.A2(n_75),
.B(n_74),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_578),
.A2(n_77),
.B(n_76),
.Y(n_643)
);

AO31x2_ASAP7_75t_L g644 ( 
.A1(n_575),
.A2(n_172),
.A3(n_258),
.B(n_257),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_SL g645 ( 
.A1(n_568),
.A2(n_36),
.B(n_37),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_605),
.A2(n_79),
.B(n_78),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_579),
.B(n_37),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_615),
.A2(n_611),
.B(n_610),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_587),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_589),
.B(n_38),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_589),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_565),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_559),
.B(n_584),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_612),
.B(n_38),
.C(n_39),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_606),
.A2(n_81),
.B(n_80),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_572),
.B(n_39),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_570),
.A2(n_82),
.B(n_83),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_596),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_616),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_594),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_584),
.B(n_259),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

AO21x2_ASAP7_75t_L g663 ( 
.A1(n_590),
.A2(n_87),
.B(n_89),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_585),
.A2(n_90),
.B(n_91),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_576),
.B(n_92),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_607),
.Y(n_666)
);

AO31x2_ASAP7_75t_L g667 ( 
.A1(n_603),
.A2(n_93),
.A3(n_97),
.B(n_98),
.Y(n_667)
);

AOI21xp33_ASAP7_75t_L g668 ( 
.A1(n_609),
.A2(n_100),
.B(n_101),
.Y(n_668)
);

NAND2x1p5_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_599),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_595),
.A2(n_601),
.B(n_614),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_102),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_592),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_596),
.B(n_600),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_604),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_613),
.A2(n_104),
.B(n_105),
.C(n_107),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_582),
.A2(n_109),
.B(n_110),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_608),
.B(n_111),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_625),
.A2(n_588),
.B(n_591),
.C(n_119),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_651),
.B(n_591),
.Y(n_679)
);

OR2x2_ASAP7_75t_SL g680 ( 
.A(n_654),
.B(n_114),
.Y(n_680)
);

OAI21xp33_ASAP7_75t_L g681 ( 
.A1(n_645),
.A2(n_117),
.B(n_121),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_635),
.B(n_256),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_628),
.A2(n_122),
.B(n_123),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_672),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_651),
.B(n_124),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g686 ( 
.A1(n_624),
.A2(n_126),
.B(n_128),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_620),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_623),
.B(n_134),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_633),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_635),
.B(n_255),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_649),
.B(n_135),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_626),
.B(n_627),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_633),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_SL g695 ( 
.A1(n_668),
.A2(n_643),
.B(n_641),
.C(n_657),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_635),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_619),
.A2(n_136),
.B(n_137),
.C(n_138),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_639),
.B(n_139),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_659),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_674),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_631),
.A2(n_140),
.B(n_141),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_645),
.A2(n_142),
.B(n_143),
.C(n_144),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_145),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_658),
.A2(n_146),
.B(n_147),
.C(n_148),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_618),
.B(n_149),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_632),
.A2(n_673),
.B1(n_654),
.B2(n_636),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_633),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_660),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_653),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_632),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_618),
.B(n_158),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_670),
.A2(n_159),
.B(n_160),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_622),
.B(n_161),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_647),
.A2(n_162),
.B(n_163),
.C(n_164),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_668),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_652),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_666),
.B(n_661),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_656),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_666),
.B(n_254),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_669),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_677),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_671),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_640),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_675),
.A2(n_168),
.B(n_169),
.C(n_170),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_629),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_621),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_665),
.B(n_253),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_718),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_690),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_703),
.A2(n_663),
.B1(n_676),
.B2(n_655),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_718),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_684),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_682),
.B(n_644),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_693),
.Y(n_737)
);

BUFx10_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_687),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_699),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_700),
.Y(n_741)
);

OA21x2_ASAP7_75t_L g742 ( 
.A1(n_728),
.A2(n_630),
.B(n_648),
.Y(n_742)
);

BUFx12f_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_707),
.A2(n_663),
.B1(n_664),
.B2(n_642),
.Y(n_744)
);

INVx8_ASAP7_75t_L g745 ( 
.A(n_682),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_679),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_720),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_705),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_681),
.A2(n_725),
.B1(n_724),
.B2(n_721),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_719),
.B(n_644),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_709),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_729),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_715),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_678),
.A2(n_646),
.B(n_638),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_696),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_726),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_712),
.A2(n_644),
.B1(n_667),
.B2(n_175),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_690),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_690),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_694),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_680),
.A2(n_702),
.B1(n_704),
.B2(n_692),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_694),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_691),
.A2(n_667),
.B1(n_174),
.B2(n_176),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_710),
.B(n_667),
.Y(n_765)
);

AO21x2_ASAP7_75t_L g766 ( 
.A1(n_695),
.A2(n_714),
.B(n_717),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_694),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_685),
.B(n_252),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_701),
.A2(n_171),
.B(n_178),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_708),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_683),
.A2(n_182),
.B(n_183),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_708),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_698),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_708),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_713),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_776)
);

BUFx2_ASAP7_75t_R g777 ( 
.A(n_706),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_723),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_697),
.A2(n_197),
.B(n_198),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_691),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_722),
.Y(n_781)
);

AO21x2_ASAP7_75t_L g782 ( 
.A1(n_716),
.A2(n_205),
.B(n_207),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_727),
.A2(n_208),
.B(n_209),
.Y(n_783)
);

AO21x2_ASAP7_75t_L g784 ( 
.A1(n_688),
.A2(n_210),
.B(n_211),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_689),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_726),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_710),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_693),
.B(n_212),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_693),
.B(n_251),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_746),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_737),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_736),
.B(n_213),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_740),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_741),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_734),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_790),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_752),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_790),
.Y(n_802)
);

BUFx2_ASAP7_75t_SL g803 ( 
.A(n_738),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_751),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_752),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_747),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_762),
.A2(n_215),
.B(n_216),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_786),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_758),
.A2(n_217),
.B(n_218),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_756),
.Y(n_810)
);

AO21x1_ASAP7_75t_SL g811 ( 
.A1(n_753),
.A2(n_219),
.B(n_220),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_750),
.B(n_221),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_747),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_748),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_786),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

AO21x1_ASAP7_75t_SL g817 ( 
.A1(n_744),
.A2(n_223),
.B(n_224),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_758),
.A2(n_765),
.B(n_754),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_745),
.B(n_225),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_748),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_743),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_786),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_755),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_773),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_756),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_742),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_742),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_735),
.B(n_230),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_781),
.B(n_233),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_773),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_779),
.A2(n_234),
.B(n_235),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_742),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_736),
.B(n_763),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_736),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_785),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_763),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_759),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_771),
.A2(n_783),
.B(n_757),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_749),
.A2(n_236),
.B(n_238),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_782),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_745),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_782),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_801),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_794),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_794),
.B(n_745),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_834),
.B(n_782),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_787),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_833),
.B(n_738),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_805),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_833),
.B(n_738),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_834),
.B(n_770),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_836),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_807),
.A2(n_745),
.B1(n_733),
.B2(n_764),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_808),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_818),
.B(n_808),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_805),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_816),
.B(n_787),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_792),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_793),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_839),
.A2(n_831),
.B1(n_743),
.B2(n_842),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_818),
.B(n_770),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_822),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_835),
.B(n_772),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_795),
.B(n_770),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_806),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_816),
.B(n_789),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_818),
.B(n_759),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_822),
.B(n_732),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_797),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_798),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_796),
.B(n_759),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_822),
.B(n_732),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_799),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_800),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_802),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_823),
.B(n_774),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_815),
.B(n_774),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_815),
.B(n_774),
.Y(n_879)
);

INVx5_ASAP7_75t_SL g880 ( 
.A(n_819),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_824),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_810),
.B(n_732),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_842),
.B(n_784),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_826),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_841),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_803),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_810),
.B(n_784),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_814),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_826),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_820),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_848),
.B(n_803),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_848),
.B(n_841),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_850),
.B(n_825),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_855),
.B(n_827),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_853),
.B(n_828),
.C(n_837),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_860),
.B(n_812),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_843),
.B(n_812),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_855),
.B(n_827),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_850),
.B(n_832),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_859),
.B(n_825),
.Y(n_901)
);

NAND3xp33_ASAP7_75t_L g902 ( 
.A(n_862),
.B(n_840),
.C(n_829),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_862),
.B(n_840),
.C(n_829),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_884),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_858),
.B(n_832),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_880),
.B(n_794),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_886),
.B(n_847),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_883),
.A2(n_788),
.B1(n_775),
.B2(n_780),
.C(n_831),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_858),
.B(n_813),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_878),
.B(n_817),
.Y(n_910)
);

OAI221xp5_ASAP7_75t_L g911 ( 
.A1(n_861),
.A2(n_821),
.B1(n_839),
.B2(n_768),
.C(n_819),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_878),
.B(n_817),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_847),
.B(n_831),
.Y(n_913)
);

NAND3xp33_ASAP7_75t_L g914 ( 
.A(n_868),
.B(n_839),
.C(n_776),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_867),
.B(n_760),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_867),
.B(n_760),
.Y(n_916)
);

OAI221xp5_ASAP7_75t_L g917 ( 
.A1(n_883),
.A2(n_819),
.B1(n_778),
.B2(n_769),
.C(n_767),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_844),
.B(n_735),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_SL g919 ( 
.A1(n_888),
.A2(n_777),
.B(n_811),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_849),
.B(n_767),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_L g921 ( 
.A1(n_888),
.A2(n_809),
.B1(n_784),
.B2(n_766),
.C(n_767),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_868),
.B(n_819),
.C(n_761),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_854),
.B(n_838),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_852),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_SL g925 ( 
.A(n_857),
.B(n_811),
.C(n_761),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_924),
.B(n_900),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_895),
.B(n_854),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_895),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_899),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_900),
.B(n_879),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_919),
.B(n_885),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_910),
.B(n_882),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_901),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_904),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_894),
.B(n_879),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_905),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_899),
.B(n_849),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_909),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_898),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_912),
.B(n_882),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_923),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_923),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_915),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_916),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_920),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_907),
.B(n_852),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_892),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_907),
.B(n_885),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_893),
.B(n_863),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_925),
.B(n_922),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_939),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_939),
.B(n_856),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_931),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_948),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_937),
.B(n_856),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_934),
.B(n_897),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_932),
.B(n_913),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_944),
.Y(n_959)
);

AND2x4_ASAP7_75t_SL g960 ( 
.A(n_947),
.B(n_845),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_946),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_940),
.B(n_857),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_926),
.B(n_913),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_931),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_937),
.B(n_896),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_944),
.B(n_864),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_961),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_955),
.B(n_932),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_965),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_954),
.B(n_943),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_964),
.B(n_933),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_961),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_953),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_953),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_963),
.B(n_933),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_962),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_965),
.B(n_945),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_958),
.B(n_943),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_959),
.B(n_945),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_977),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_969),
.A2(n_921),
.B(n_951),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_967),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_972),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_969),
.B(n_966),
.Y(n_984)
);

INVxp67_ASAP7_75t_SL g985 ( 
.A(n_968),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_979),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_976),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_980),
.B(n_976),
.Y(n_988)
);

NOR2x1_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_978),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_981),
.A2(n_974),
.B1(n_973),
.B2(n_978),
.C(n_957),
.Y(n_990)
);

OAI221xp5_ASAP7_75t_SL g991 ( 
.A1(n_984),
.A2(n_911),
.B1(n_908),
.B2(n_917),
.C(n_970),
.Y(n_991)
);

AOI322xp5_ASAP7_75t_L g992 ( 
.A1(n_987),
.A2(n_942),
.A3(n_970),
.B1(n_929),
.B2(n_930),
.C1(n_952),
.C2(n_971),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_988),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_989),
.B(n_986),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_991),
.B(n_982),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_975),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_990),
.B(n_985),
.Y(n_997)
);

NOR3x1_ASAP7_75t_L g998 ( 
.A(n_994),
.B(n_983),
.C(n_968),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_994),
.A2(n_956),
.B(n_947),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_997),
.A2(n_914),
.B1(n_942),
.B2(n_906),
.Y(n_1000)
);

AOI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_993),
.A2(n_902),
.B1(n_903),
.B2(n_956),
.C(n_946),
.Y(n_1001)
);

OAI32xp33_ASAP7_75t_L g1002 ( 
.A1(n_995),
.A2(n_948),
.A3(n_927),
.B1(n_926),
.B2(n_938),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_996),
.A2(n_933),
.B1(n_941),
.B2(n_960),
.Y(n_1003)
);

OAI211xp5_ASAP7_75t_SL g1004 ( 
.A1(n_994),
.A2(n_877),
.B(n_906),
.C(n_872),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_1003),
.Y(n_1006)
);

NOR3x1_ASAP7_75t_L g1007 ( 
.A(n_1002),
.B(n_863),
.C(n_865),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_1004),
.B(n_771),
.C(n_783),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_SL g1010 ( 
.A(n_1001),
.B(n_918),
.C(n_761),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1009),
.B(n_1006),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_1005),
.B(n_1000),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_935),
.C(n_928),
.Y(n_1013)
);

OAI211xp5_ASAP7_75t_SL g1014 ( 
.A1(n_1010),
.A2(n_935),
.B(n_928),
.C(n_918),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_SL g1015 ( 
.A(n_1007),
.B(n_870),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_SL g1016 ( 
.A(n_1005),
.B(n_949),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1009),
.Y(n_1017)
);

NOR2x1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_949),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1011),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1018),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1017),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_1012),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_1014),
.B(n_941),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1016),
.Y(n_1024)
);

NOR2x1_ASAP7_75t_L g1025 ( 
.A(n_1015),
.B(n_941),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1013),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1011),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1012),
.A2(n_880),
.B1(n_845),
.B2(n_809),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1018),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1012),
.A2(n_880),
.B1(n_845),
.B2(n_809),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1011),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1011),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1011),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1011),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1022),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1024),
.B(n_936),
.Y(n_1037)
);

OR3x1_ASAP7_75t_L g1038 ( 
.A(n_1019),
.B(n_880),
.C(n_950),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_838),
.C(n_887),
.Y(n_1039)
);

AO221x2_ASAP7_75t_L g1040 ( 
.A1(n_1027),
.A2(n_950),
.B1(n_936),
.B2(n_873),
.C(n_869),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_L g1041 ( 
.A(n_1031),
.B(n_887),
.C(n_884),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_1032),
.B(n_870),
.C(n_871),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1033),
.A2(n_882),
.B(n_769),
.Y(n_1043)
);

AND3x4_ASAP7_75t_L g1044 ( 
.A(n_1023),
.B(n_873),
.C(n_869),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_845),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1029),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1025),
.A2(n_844),
.B1(n_766),
.B2(n_846),
.Y(n_1047)
);

AND2x2_ASAP7_75t_SL g1048 ( 
.A(n_1021),
.B(n_769),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_1026),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_1028),
.B(n_869),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1030),
.A2(n_873),
.B1(n_844),
.B2(n_884),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1022),
.B(n_890),
.C(n_871),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1035),
.B(n_890),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_1046),
.B(n_844),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_1037),
.Y(n_1055)
);

XOR2x1_ASAP7_75t_L g1056 ( 
.A(n_1036),
.B(n_882),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1040),
.B(n_890),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1038),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1044),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_1049),
.Y(n_1060)
);

OAI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1045),
.A2(n_875),
.B1(n_874),
.B2(n_889),
.Y(n_1061)
);

NAND3x1_ASAP7_75t_L g1062 ( 
.A(n_1041),
.B(n_1043),
.C(n_1047),
.Y(n_1062)
);

AO22x2_ASAP7_75t_L g1063 ( 
.A1(n_1060),
.A2(n_1055),
.B1(n_1058),
.B2(n_1059),
.Y(n_1063)
);

AOI22x1_ASAP7_75t_L g1064 ( 
.A1(n_1057),
.A2(n_1050),
.B1(n_1040),
.B2(n_1042),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1062),
.A2(n_1048),
.B1(n_1039),
.B2(n_1051),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1053),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1056),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1061),
.Y(n_1068)
);

OAI321xp33_ASAP7_75t_L g1069 ( 
.A1(n_1067),
.A2(n_1054),
.A3(n_1052),
.B1(n_844),
.B2(n_874),
.C(n_875),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_766),
.B1(n_846),
.B2(n_889),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_1068),
.B(n_1066),
.C(n_1063),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1064),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1072),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1071),
.B(n_1070),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1073),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_1069),
.B(n_846),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1074),
.A2(n_846),
.B1(n_881),
.B2(n_876),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1075),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_SL g1079 ( 
.A1(n_1076),
.A2(n_239),
.B(n_240),
.Y(n_1079)
);

OA22x2_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_1079),
.B1(n_1077),
.B2(n_851),
.Y(n_1080)
);

AOI221xp5_ASAP7_75t_L g1081 ( 
.A1(n_1078),
.A2(n_881),
.B1(n_876),
.B2(n_891),
.C(n_851),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1080),
.A2(n_891),
.B(n_866),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_R g1083 ( 
.A1(n_1082),
.A2(n_1081),
.B1(n_242),
.B2(n_243),
.C(n_244),
.Y(n_1083)
);

AOI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_241),
.B(n_246),
.C(n_247),
.Y(n_1084)
);


endmodule