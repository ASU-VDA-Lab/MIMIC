module real_jpeg_5991_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_0),
.A2(n_159),
.B1(n_163),
.B2(n_166),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_0),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_0),
.B(n_179),
.C(n_183),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_0),
.B(n_73),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_0),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_0),
.B(n_125),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_0),
.B(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_1),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_1),
.Y(n_293)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_1),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_2),
.A2(n_62),
.B1(n_211),
.B2(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_2),
.A2(n_62),
.B1(n_81),
.B2(n_219),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_2),
.A2(n_62),
.B1(n_378),
.B2(n_455),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_98),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_98),
.B1(n_135),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_3),
.A2(n_98),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_4),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_4),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_4),
.Y(n_368)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_4),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_4),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g441 ( 
.A(n_4),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_5),
.A2(n_51),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_5),
.A2(n_51),
.B1(n_219),
.B2(n_403),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_5),
.A2(n_51),
.B1(n_295),
.B2(n_413),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_6),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_8),
.A2(n_190),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_8),
.A2(n_159),
.B1(n_195),
.B2(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_8),
.A2(n_195),
.B1(n_375),
.B2(n_377),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_8),
.A2(n_195),
.B1(n_416),
.B2(n_418),
.Y(n_415)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_9),
.Y(n_544)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_12),
.A2(n_170),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_12),
.A2(n_170),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_12),
.A2(n_170),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_86),
.B1(n_88),
.B2(n_92),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_15),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_15),
.A2(n_92),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_15),
.A2(n_92),
.B1(n_241),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_15),
.A2(n_92),
.B1(n_382),
.B2(n_423),
.Y(n_422)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_17),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_17),
.A2(n_221),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_17),
.A2(n_221),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_17),
.A2(n_221),
.B1(n_440),
.B2(n_442),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_18),
.A2(n_283),
.B1(n_287),
.B2(n_288),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_18),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_18),
.A2(n_105),
.B1(n_287),
.B2(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_18),
.A2(n_287),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_L g467 ( 
.A1(n_18),
.A2(n_287),
.B1(n_362),
.B2(n_468),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_542),
.B(n_545),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_148),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_146),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_139),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_23),
.B(n_139),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_130),
.C(n_136),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_24),
.A2(n_25),
.B1(n_538),
.B2(n_539),
.Y(n_537)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_63),
.C(n_99),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_26),
.B(n_530),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_27),
.A2(n_52),
.B1(n_131),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_27),
.A2(n_366),
.B(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_27),
.A2(n_40),
.B1(n_415),
.B2(n_439),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_28),
.A2(n_361),
.B(n_365),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_28),
.B(n_367),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_39),
.Y(n_343)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_40),
.B(n_166),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_40)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_41),
.Y(n_341)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_43),
.Y(n_278)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_44),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_45),
.Y(n_315)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_46),
.Y(n_376)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_46),
.Y(n_379)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_47),
.Y(n_277)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_52),
.A2(n_439),
.B(n_469),
.Y(n_479)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_53),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_53),
.B(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_57),
.Y(n_443)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_63),
.A2(n_99),
.B1(n_100),
.B2(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_63),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_64),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_64),
.A2(n_93),
.B1(n_313),
.B2(n_374),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_64),
.A2(n_93),
.B1(n_409),
.B2(n_412),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_64),
.A2(n_85),
.B1(n_93),
.B2(n_519),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_73),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_67),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_69),
.Y(n_410)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_70),
.Y(n_302)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

AOI22x1_ASAP7_75t_L g444 ( 
.A1(n_73),
.A2(n_137),
.B1(n_317),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_73),
.A2(n_137),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_79),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_80),
.Y(n_296)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_80),
.Y(n_405)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_93),
.B(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_93),
.A2(n_313),
.B(n_316),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_95),
.Y(n_411)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_99),
.A2(n_100),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_99),
.B(n_514),
.C(n_517),
.Y(n_525)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_124),
.B(n_126),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_158),
.B(n_167),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_101),
.A2(n_124),
.B1(n_218),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_101),
.A2(n_167),
.B(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_101),
.A2(n_124),
.B1(n_381),
.B2(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_102),
.B(n_168),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_102),
.A2(n_125),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_102),
.A2(n_125),
.B1(n_406),
.B2(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_102),
.A2(n_125),
.B1(n_422),
.B2(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_106),
.Y(n_223)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_113),
.A2(n_218),
.B(n_224),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_121),
.Y(n_242)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_121),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_121),
.Y(n_398)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_124),
.A2(n_224),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_126),
.Y(n_458)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_130),
.B(n_136),
.Y(n_539)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_137),
.A2(n_269),
.B(n_275),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_137),
.B(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_137),
.A2(n_275),
.B(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_143),
.B(n_166),
.Y(n_347)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_536),
.B(n_541),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_508),
.B(n_533),
.Y(n_149)
);

OAI311xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_386),
.A3(n_484),
.B1(n_502),
.C1(n_503),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_331),
.B(n_385),
.Y(n_151)
);

AO21x1_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_304),
.B(n_330),
.Y(n_152)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_257),
.B(n_303),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_227),
.B(n_256),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_187),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_156),
.B(n_187),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_173),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_157),
.A2(n_173),
.B1(n_174),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_165),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_166),
.A2(n_199),
.B(n_207),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g269 ( 
.A1(n_166),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_166),
.A2(n_347),
.B(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_186),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_215),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_188),
.B(n_216),
.C(n_226),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_199),
.B(n_207),
.Y(n_188)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_194),
.Y(n_395)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_198),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_199),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_199),
.A2(n_392),
.B1(n_396),
.B2(n_397),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_199),
.A2(n_397),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_210),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_208),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_200),
.A2(n_282),
.B1(n_321),
.B2(n_327),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_200),
.A2(n_353),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_203),
.Y(n_328)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_203),
.Y(n_436)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_225),
.B2(n_226),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_222),
.B(n_301),
.Y(n_300)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_249),
.B(n_255),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_237),
.B(n_248),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_233),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_247),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_247),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_245),
.B(n_246),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_281),
.B(n_291),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_259),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_279),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_267),
.B2(n_268),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_262),
.B(n_267),
.C(n_279),
.Y(n_305)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI32xp33_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_295),
.A3(n_296),
.B1(n_297),
.B2(n_300),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_294),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_294),
.Y(n_310)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_305),
.B(n_306),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_311),
.B2(n_329),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_310),
.C(n_329),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_319),
.C(n_320),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_315),
.A2(n_338),
.A3(n_340),
.B1(n_342),
.B2(n_347),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_332),
.B(n_333),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_358),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_348),
.B2(n_349),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_337),
.B(n_348),
.Y(n_480)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_355),
.B(n_356),
.C(n_358),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_372),
.B2(n_384),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_359),
.B(n_373),
.C(n_380),
.Y(n_493)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_470),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_387),
.A2(n_470),
.B(n_504),
.C(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_446),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_388),
.B(n_446),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_419),
.C(n_429),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g483 ( 
.A(n_389),
.B(n_419),
.CI(n_429),
.CON(n_483),
.SN(n_483)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_407),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_390),
.B(n_408),
.C(n_414),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_401),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_391),
.B(n_401),
.Y(n_476)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

INVx4_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_414),
.Y(n_407)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_425),
.B2(n_428),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_425),
.Y(n_462)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_425),
.A2(n_428),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_425),
.A2(n_462),
.B(n_465),
.Y(n_511)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_437),
.C(n_444),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_431),
.B(n_433),
.Y(n_492)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_437),
.A2(n_438),
.B1(n_444),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_444),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_450),
.C(n_460),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_460),
.B2(n_461),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_456),
.B(n_459),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_457),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_454),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_459),
.B(n_511),
.CI(n_512),
.CON(n_510),
.SN(n_510)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_459),
.B(n_511),
.C(n_512),
.Y(n_532)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_467),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_483),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_471),
.B(n_483),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_476),
.C(n_477),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_472),
.A2(n_473),
.B1(n_476),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_480),
.C(n_481),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_478),
.A2(n_479),
.B1(n_481),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_481),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_483),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_497),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_505),
.B(n_506),
.Y(n_504)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_494),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_494),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_491),
.C(n_493),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_500),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_492),
.B1(n_493),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_493),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_499),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_522),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_521),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_521),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g548 ( 
.A(n_510),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_516),
.B2(n_520),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_513),
.A2(n_514),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_524),
.C(n_528),
.Y(n_540)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_516),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_522),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_523),
.B(n_532),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_532),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_525),
.B1(n_526),
.B2(n_527),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_540),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_540),
.Y(n_541)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_543),
.Y(n_546)
);

INVx13_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_547),
.Y(n_545)
);


endmodule