module fake_jpeg_13338_n_454 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_48),
.Y(n_140)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_50),
.Y(n_127)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_78),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_6),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_79),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_8),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_95),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_38),
.B(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_34),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_96),
.B(n_135),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_18),
.B1(n_15),
.B2(n_39),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_109),
.B1(n_114),
.B2(n_122),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_36),
.B(n_33),
.C(n_43),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_106),
.B(n_120),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_18),
.B1(n_15),
.B2(n_30),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_110),
.A2(n_0),
.B(n_2),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_54),
.A2(n_18),
.B1(n_34),
.B2(n_68),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_36),
.B(n_43),
.C(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_56),
.A2(n_34),
.B1(n_32),
.B2(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_146),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_59),
.A2(n_40),
.B1(n_31),
.B2(n_21),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_139),
.B1(n_101),
.B2(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_28),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_62),
.A2(n_21),
.B1(n_40),
.B2(n_31),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_140),
.B1(n_125),
.B2(n_127),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_31),
.B1(n_40),
.B2(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_47),
.B(n_31),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_63),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_64),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_153),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_98),
.B(n_40),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_155),
.B(n_172),
.Y(n_223)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_94),
.B1(n_93),
.B2(n_88),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_111),
.B1(n_147),
.B2(n_105),
.Y(n_225)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_180),
.B1(n_109),
.B2(n_114),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_87),
.C(n_85),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_192),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_101),
.A2(n_116),
.B1(n_113),
.B2(n_40),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_163),
.Y(n_217)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_73),
.B1(n_70),
.B2(n_41),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_167),
.Y(n_222)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_41),
.C(n_8),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_8),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_188),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_184),
.Y(n_213)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_107),
.B(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_97),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_5),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_121),
.B(n_9),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_198),
.A2(n_153),
.B1(n_168),
.B2(n_151),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_190),
.B(n_161),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_152),
.B(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_112),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_214),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_130),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_130),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_228),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_133),
.B1(n_132),
.B2(n_136),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_171),
.B(n_121),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_157),
.B1(n_165),
.B2(n_164),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_231),
.A2(n_243),
.B1(n_252),
.B2(n_260),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_224),
.C(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_180),
.B1(n_147),
.B2(n_111),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_239),
.B1(n_242),
.B2(n_256),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_215),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_214),
.A2(n_170),
.B(n_127),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_193),
.B1(n_192),
.B2(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_249),
.B1(n_250),
.B2(n_212),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_102),
.B1(n_136),
.B2(n_132),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_203),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_169),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_174),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_119),
.B1(n_123),
.B2(n_145),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_202),
.A2(n_119),
.B1(n_123),
.B2(n_145),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_217),
.A2(n_154),
.B1(n_166),
.B2(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_202),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_179),
.B1(n_175),
.B2(n_177),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_158),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_212),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_225),
.B1(n_197),
.B2(n_216),
.Y(n_288)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_217),
.A2(n_178),
.B1(n_162),
.B2(n_143),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_265),
.C(n_232),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_224),
.C(n_223),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_256),
.B1(n_239),
.B2(n_260),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_278),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_273),
.B(n_279),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_280),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_197),
.B(n_215),
.C(n_206),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_206),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_246),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_281),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_257),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_282),
.Y(n_295)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_197),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_259),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_286),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_216),
.B1(n_203),
.B2(n_211),
.Y(n_311)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_290),
.B(n_208),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_258),
.B(n_234),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_292),
.A2(n_266),
.B(n_276),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_232),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_304),
.C(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_267),
.A2(n_231),
.B1(n_268),
.B2(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_296),
.A2(n_307),
.B1(n_313),
.B2(n_274),
.Y(n_340)
);

XOR2x1_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_237),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_211),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_258),
.B(n_235),
.Y(n_300)
);

AOI21x1_ASAP7_75t_SL g341 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_270),
.A2(n_247),
.B(n_242),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_233),
.B(n_253),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_241),
.B1(n_249),
.B2(n_250),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_303),
.A2(n_311),
.B1(n_218),
.B2(n_209),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_265),
.B(n_280),
.C(n_269),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_277),
.C(n_281),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_245),
.B(n_240),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_286),
.B(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_314),
.Y(n_323)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_263),
.A2(n_209),
.B1(n_218),
.B2(n_219),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_276),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_334),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_283),
.B1(n_275),
.B2(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_328),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_324),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_283),
.Y(n_322)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_295),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_329),
.Y(n_359)
);

XOR2x2_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_272),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_301),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_296),
.A2(n_289),
.B1(n_287),
.B2(n_284),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_333),
.B(n_292),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_226),
.C(n_219),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_336),
.C(n_308),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_304),
.B(n_243),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_332),
.B(n_306),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_315),
.A2(n_200),
.B(n_210),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_200),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_335),
.B(n_338),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_210),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_307),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_274),
.Y(n_339)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_340),
.A2(n_342),
.B1(n_303),
.B2(n_311),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_292),
.A2(n_274),
.B1(n_230),
.B2(n_208),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_201),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_201),
.Y(n_345)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_345),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_347),
.A2(n_368),
.B1(n_320),
.B2(n_313),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_348),
.A2(n_318),
.B(n_339),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_298),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_316),
.Y(n_353)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_334),
.B(n_317),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_369),
.C(n_338),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_306),
.B1(n_302),
.B2(n_298),
.Y(n_362)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_344),
.B1(n_293),
.B2(n_230),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_292),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_367),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_314),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_330),
.A2(n_313),
.B1(n_312),
.B2(n_310),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_383),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_326),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_371),
.B(n_384),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_336),
.C(n_331),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_375),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_335),
.C(n_328),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_363),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_353),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_321),
.C(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_380),
.C(n_357),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_350),
.B1(n_349),
.B2(n_346),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_341),
.C(n_333),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_323),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_352),
.A2(n_342),
.B1(n_344),
.B2(n_308),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_347),
.B1(n_368),
.B2(n_360),
.Y(n_404)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_388),
.Y(n_398)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_405),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_355),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_143),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_374),
.C(n_370),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_394),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_380),
.A2(n_350),
.B(n_387),
.Y(n_394)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_378),
.A2(n_358),
.B(n_348),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_399),
.A2(n_375),
.B(n_381),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_383),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_379),
.Y(n_409)
);

OAI221xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_354),
.B1(n_361),
.B2(n_355),
.C(n_293),
.Y(n_405)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_382),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_414),
.Y(n_423)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

BUFx4f_ASAP7_75t_SL g416 ( 
.A(n_404),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_418),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_382),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_419),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g418 ( 
.A(n_390),
.B(n_386),
.CI(n_10),
.CON(n_418),
.SN(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_392),
.C(n_400),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_422),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_401),
.C(n_393),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_401),
.C(n_389),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_428),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_395),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_426),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_394),
.C(n_399),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_430),
.B(n_431),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_143),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_420),
.B(n_415),
.Y(n_432)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_432),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_427),
.A2(n_406),
.B(n_408),
.C(n_418),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_436),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_429),
.B(n_416),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_416),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_424),
.B1(n_425),
.B2(n_421),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_9),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_9),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_442),
.A2(n_9),
.B(n_11),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_434),
.A2(n_440),
.B(n_432),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_445),
.C(n_439),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_447),
.C(n_448),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_433),
.C(n_422),
.Y(n_447)
);

AOI321xp33_ASAP7_75t_L g449 ( 
.A1(n_447),
.A2(n_441),
.A3(n_444),
.B1(n_3),
.B2(n_4),
.C(n_10),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_449),
.B(n_4),
.C(n_11),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_451),
.A2(n_450),
.B(n_4),
.Y(n_452)
);

OAI21x1_ASAP7_75t_SL g453 ( 
.A1(n_452),
.A2(n_13),
.B(n_0),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_13),
.B(n_2),
.Y(n_454)
);


endmodule