module fake_jpeg_6053_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_40),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_53),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_51),
.Y(n_68)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_64),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_63),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_40),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_33),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_27),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_91),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_37),
.B1(n_22),
.B2(n_30),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_92),
.B1(n_95),
.B2(n_100),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_86),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_98),
.B1(n_99),
.B2(n_50),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_50),
.B1(n_22),
.B2(n_29),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_87),
.A2(n_45),
.B1(n_44),
.B2(n_10),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_45),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_20),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_25),
.B1(n_20),
.B2(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_15),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_20),
.C(n_34),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_0),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_3),
.Y(n_134)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_34),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_91),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_45),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_132),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_94),
.B1(n_86),
.B2(n_67),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_13),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_2),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_125),
.B(n_116),
.C(n_120),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_70),
.B1(n_84),
.B2(n_81),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_3),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_101),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_97),
.B1(n_100),
.B2(n_58),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_143),
.B1(n_157),
.B2(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_61),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_144),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_68),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_142),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_70),
.B1(n_58),
.B2(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_59),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_77),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_77),
.Y(n_151)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_164),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_62),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_102),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_57),
.B(n_103),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.C(n_166),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_123),
.B(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_63),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_159),
.B1(n_169),
.B2(n_124),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_74),
.B(n_62),
.C(n_72),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_82),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_67),
.B1(n_62),
.B2(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_112),
.B(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_62),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_56),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_3),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_4),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_179),
.B1(n_186),
.B2(n_205),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_125),
.B1(n_113),
.B2(n_128),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_113),
.B(n_134),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_197),
.B(n_151),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_128),
.B1(n_106),
.B2(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_164),
.B(n_106),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_111),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_152),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_107),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_147),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_133),
.B1(n_130),
.B2(n_111),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_143),
.A2(n_130),
.B1(n_117),
.B2(n_119),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_117),
.B1(n_119),
.B2(n_56),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_140),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_139),
.A2(n_119),
.B1(n_7),
.B2(n_8),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_224),
.B1(n_234),
.B2(n_235),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_153),
.B1(n_159),
.B2(n_161),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_217),
.B(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_137),
.B(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_225),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_180),
.B1(n_199),
.B2(n_178),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_236),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_150),
.B(n_142),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_146),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_149),
.C(n_148),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_231),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_155),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_230),
.C(n_233),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_146),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_176),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_196),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_141),
.C(n_154),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_159),
.B1(n_169),
.B2(n_172),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_177),
.A2(n_207),
.B1(n_190),
.B2(n_193),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_145),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_163),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_194),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_244),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_248),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_216),
.A2(n_210),
.B1(n_199),
.B2(n_203),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_260),
.B1(n_185),
.B2(n_226),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_192),
.B(n_178),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_257),
.B(n_181),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_258),
.B1(n_197),
.B2(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_175),
.B1(n_179),
.B2(n_190),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_217),
.B1(n_214),
.B2(n_206),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_218),
.A2(n_203),
.B1(n_196),
.B2(n_206),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_251),
.B(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_237),
.C(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_233),
.C(n_228),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_222),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_277),
.C(n_248),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_205),
.B1(n_232),
.B2(n_224),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_214),
.C(n_201),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_231),
.C(n_197),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_186),
.C(n_226),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_241),
.B(n_189),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_184),
.C(n_185),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_272),
.B(n_277),
.C(n_255),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_284),
.B(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

INVxp33_ASAP7_75t_SL g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_289),
.C(n_276),
.Y(n_292)
);

OAI322xp33_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_251),
.A3(n_239),
.B1(n_259),
.B2(n_242),
.C1(n_244),
.C2(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_269),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_256),
.A3(n_239),
.B1(n_247),
.B2(n_254),
.C1(n_241),
.C2(n_195),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_224),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_302),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_306)
);

NAND4xp25_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_182),
.C(n_102),
.D(n_208),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_300),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_282),
.B(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_264),
.B1(n_263),
.B2(n_157),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_279),
.B1(n_281),
.B2(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_278),
.B(n_171),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_278),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_292),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_310),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_281),
.B(n_173),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_5),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_296),
.A2(n_279),
.B1(n_107),
.B2(n_83),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_145),
.A3(n_183),
.B1(n_162),
.B2(n_83),
.C1(n_56),
.C2(n_14),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_313),
.B(n_317),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_309),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_311),
.Y(n_319)
);

AOI31xp33_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_14),
.A3(n_5),
.B(n_8),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_310),
.B1(n_10),
.B2(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_14),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_315),
.B(n_318),
.C(n_313),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_322),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_321),
.Y(n_327)
);


endmodule