module fake_jpeg_20107_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_20),
.Y(n_45)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_15),
.B1(n_25),
.B2(n_23),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_14),
.B1(n_25),
.B2(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_43),
.B1(n_29),
.B2(n_36),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_22),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_38),
.B(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_16),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_61),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_60),
.B1(n_33),
.B2(n_30),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_33),
.B1(n_35),
.B2(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_35),
.B(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_42),
.B1(n_43),
.B2(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_79),
.B1(n_51),
.B2(n_49),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_75),
.B(n_53),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_24),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_21),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_39),
.B(n_35),
.C(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_76),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_86),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_83),
.B1(n_65),
.B2(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_24),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_90),
.B(n_93),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OA21x2_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_50),
.B(n_27),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_66),
.C(n_85),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_97),
.B(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_68),
.C(n_67),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_79),
.B1(n_73),
.B2(n_75),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_92),
.B1(n_82),
.B2(n_3),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

XNOR2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_74),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_112),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_80),
.B(n_83),
.C(n_89),
.D(n_91),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_97),
.C(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_118),
.C(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_95),
.C(n_98),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_109),
.B(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_17),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_82),
.C(n_109),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_8),
.B(n_11),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_7),
.B(n_12),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_27),
.C(n_6),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_115),
.C(n_27),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_10),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_11),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_10),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_133),
.B(n_1),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_135),
.B(n_4),
.Y(n_136)
);

AOI21x1_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_2),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_3),
.Y(n_138)
);


endmodule