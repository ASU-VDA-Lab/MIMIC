module fake_netlist_6_714_n_2424 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2424);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2424;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_107),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_66),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_17),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_69),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_133),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_75),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_22),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_34),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_40),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_98),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_129),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_103),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_69),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_106),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_102),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_78),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_8),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_138),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_122),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_88),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_9),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_229),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_10),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_179),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_79),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_14),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_102),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_113),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_192),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_108),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_152),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_16),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_71),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_123),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_199),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_0),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_209),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_91),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_99),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_115),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_57),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_92),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_158),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_134),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_80),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_234),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_114),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_140),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_35),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_159),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_71),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_93),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_55),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_2),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_223),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_8),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_92),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_108),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_202),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_6),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_126),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_0),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_67),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_70),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_68),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_172),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_225),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_169),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_168),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_31),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_76),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_56),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_58),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_33),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_28),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_22),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_63),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_34),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_143),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_25),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_125),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_176),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_215),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_77),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_43),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_42),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_110),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_89),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_35),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_191),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_146),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_38),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_212),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_15),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_77),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_21),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_17),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_2),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_84),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_100),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_203),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_165),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_13),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_147),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_26),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_38),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_52),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_211),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_149),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_144),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_148),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_52),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_120),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_93),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_100),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_44),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_59),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_67),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_81),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_132),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_73),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_214),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_85),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_15),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_182),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_150),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_128),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_195),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_70),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_119),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_40),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_208),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_205),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_224),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_90),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_20),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_157),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_19),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_4),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_164),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_57),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_37),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_36),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_84),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_130),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_49),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_96),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_155),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_154),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_112),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_27),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_31),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_207),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_78),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_142),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_189),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_55),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_63),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_39),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_99),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_101),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_74),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_151),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_36),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_97),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_194),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_1),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_30),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_47),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_124),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_41),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_97),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_190),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_5),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_117),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_85),
.Y(n_448)
);

BUFx2_ASAP7_75t_SL g449 ( 
.A(n_106),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_25),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_173),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_41),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_193),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_217),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_153),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_66),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_183),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_6),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_135),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_42),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_30),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_188),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_252),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_311),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_248),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_272),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_284),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_392),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_251),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_237),
.B(n_1),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_262),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_237),
.B(n_3),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_277),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_266),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_459),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_268),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_311),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_311),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_311),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_279),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_311),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_277),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_364),
.B(n_405),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_319),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_330),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_447),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_405),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_330),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_304),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_330),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_303),
.B(n_3),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_287),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_289),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_330),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_447),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_294),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_305),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_238),
.B(n_4),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_306),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_330),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_272),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_330),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_284),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_239),
.B(n_5),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_308),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_303),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_309),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_337),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_312),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_337),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_238),
.B(n_7),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_313),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_314),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_337),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_337),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_337),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_284),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_337),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_325),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_326),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_333),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_334),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_335),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_376),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_239),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_336),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_349),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_351),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_376),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_353),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_304),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_331),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_449),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_376),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_357),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_376),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_331),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_361),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_376),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_376),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_363),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_371),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_365),
.B(n_7),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_276),
.B(n_417),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_276),
.B(n_10),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_417),
.B(n_11),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_242),
.B(n_11),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_372),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_374),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_378),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_458),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_242),
.B(n_12),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_380),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_394),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_397),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_400),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_404),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_256),
.B(n_265),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_420),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_421),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_422),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_435),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_244),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_244),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_350),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_438),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_260),
.B(n_12),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_444),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_350),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_368),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_444),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_442),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_368),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_389),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_256),
.B(n_16),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_451),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_446),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_446),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_449),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_246),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_453),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_517),
.B(n_454),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_528),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_519),
.B(n_324),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_465),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_470),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_472),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_463),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_475),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_468),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_477),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_521),
.B(n_445),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

BUFx8_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_478),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_481),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_478),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_479),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_537),
.B(n_457),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_479),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_566),
.B(n_365),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_469),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_423),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_480),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_482),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_493),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_467),
.A2(n_302),
.B(n_286),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_482),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_494),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_484),
.B(n_434),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_511),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_514),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_502),
.B(n_505),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_492),
.B(n_296),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_522),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_497),
.B(n_235),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_534),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_523),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_466),
.B(n_286),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_487),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_476),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_489),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_489),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_525),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_488),
.B(n_265),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_491),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_526),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_533),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_491),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_495),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_550),
.B(n_423),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_501),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_501),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_503),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_503),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_541),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_510),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_510),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_512),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_512),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_544),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_504),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_518),
.B(n_302),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_527),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_527),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_532),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_532),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_246),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_539),
.B(n_316),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_520),
.A2(n_341),
.B(n_316),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_553),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_498),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_539),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_341),
.Y(n_676)
);

AND2x2_ASAP7_75t_SL g677 ( 
.A(n_551),
.B(n_296),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_554),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_542),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_535),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_543),
.B(n_425),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_496),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_543),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_548),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_548),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_549),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_555),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_466),
.B(n_425),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_666),
.B(n_558),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_609),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_669),
.B(n_466),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_591),
.B(n_560),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_602),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_666),
.B(n_561),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_602),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_609),
.Y(n_696)
);

BUFx4f_ASAP7_75t_L g697 ( 
.A(n_677),
.Y(n_697)
);

INVx6_ASAP7_75t_L g698 ( 
.A(n_635),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_635),
.B(n_267),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_627),
.B(n_574),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_666),
.B(n_580),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_677),
.B(n_267),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_629),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_635),
.B(n_269),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_609),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_688),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_669),
.B(n_579),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_680),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_635),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_677),
.B(n_269),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_595),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_591),
.B(n_590),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_594),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_594),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_599),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_598),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_598),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_601),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_SL g720 ( 
.A1(n_680),
.A2(n_575),
.B1(n_298),
.B2(n_342),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_627),
.B(n_531),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_631),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_618),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_618),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_620),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_674),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_602),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_614),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_593),
.B(n_531),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_601),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_593),
.B(n_531),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_605),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_688),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_618),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_688),
.B(n_536),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_605),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_620),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_637),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_649),
.B(n_296),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_602),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_649),
.B(n_296),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_607),
.Y(n_743)
);

BUFx2_ASAP7_75t_SL g744 ( 
.A(n_629),
.Y(n_744)
);

OR2x2_ASAP7_75t_SL g745 ( 
.A(n_613),
.B(n_490),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_672),
.B(n_271),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_613),
.B(n_588),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_623),
.B(n_507),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_596),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_597),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_621),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_666),
.B(n_490),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_672),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_604),
.B(n_549),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_607),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_632),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_687),
.B(n_535),
.Y(n_758)
);

AND2x6_ASAP7_75t_L g759 ( 
.A(n_641),
.B(n_296),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_634),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_636),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_621),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_610),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_615),
.B(n_557),
.C(n_552),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_604),
.B(n_540),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_612),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_606),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_636),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_629),
.A2(n_583),
.B1(n_485),
.B2(n_509),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_612),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_600),
.B(n_500),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_672),
.Y(n_773)
);

XNOR2xp5_ASAP7_75t_L g774 ( 
.A(n_682),
.B(n_575),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_617),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_603),
.B(n_506),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_617),
.Y(n_778)
);

BUFx4f_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_611),
.B(n_556),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_611),
.B(n_629),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_629),
.B(n_556),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_634),
.B(n_296),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_592),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_632),
.A2(n_508),
.B1(n_524),
.B2(n_516),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_629),
.B(n_271),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_616),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_592),
.B(n_559),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_592),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_625),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_617),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_616),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_592),
.B(n_559),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_592),
.B(n_564),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_564),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_617),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_625),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_638),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_663),
.B(n_293),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_608),
.B(n_529),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_639),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_639),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_634),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_639),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_615),
.A2(n_483),
.B1(n_515),
.B2(n_474),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_606),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_682),
.B(n_434),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_638),
.B(n_565),
.Y(n_808)
);

INVx4_ASAP7_75t_SL g809 ( 
.A(n_617),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_634),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_650),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_643),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_650),
.Y(n_813)
);

OA22x2_ASAP7_75t_L g814 ( 
.A1(n_663),
.A2(n_247),
.B1(n_258),
.B2(n_257),
.Y(n_814)
);

NAND3x1_ASAP7_75t_L g815 ( 
.A(n_670),
.B(n_257),
.C(n_247),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_619),
.B(n_530),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_643),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_650),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_646),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_622),
.B(n_538),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_642),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_624),
.B(n_562),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_646),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_647),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_647),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_648),
.B(n_565),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_648),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_652),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_642),
.B(n_293),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_651),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_606),
.A2(n_473),
.B1(n_546),
.B2(n_471),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_670),
.B(n_300),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_626),
.A2(n_259),
.B1(n_318),
.B2(n_243),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_651),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_652),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_630),
.B(n_563),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_652),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_653),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_653),
.B(n_528),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_676),
.B(n_499),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_676),
.B(n_499),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_655),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_633),
.B(n_567),
.Y(n_843)
);

INVx5_ASAP7_75t_L g844 ( 
.A(n_642),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_655),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_640),
.B(n_568),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_617),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_659),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_644),
.B(n_645),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_714),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_753),
.B(n_300),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_708),
.Y(n_854)
);

NAND2x1_ASAP7_75t_L g855 ( 
.A(n_725),
.B(n_642),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_700),
.B(n_606),
.Y(n_856)
);

AO22x1_ASAP7_75t_L g857 ( 
.A1(n_786),
.A2(n_310),
.B1(n_328),
.B2(n_301),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_715),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_707),
.B(n_654),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_706),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_715),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_702),
.A2(n_301),
.B1(n_328),
.B2(n_310),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_721),
.B(n_660),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_729),
.B(n_673),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_678),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_692),
.B(n_661),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_712),
.B(n_661),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_754),
.B(n_661),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_717),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_717),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_765),
.A2(n_473),
.B1(n_546),
.B2(n_471),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_697),
.A2(n_360),
.B(n_379),
.C(n_352),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_780),
.B(n_661),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_718),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_748),
.B(n_569),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_766),
.B(n_570),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_702),
.B(n_662),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_SL g878 ( 
.A(n_833),
.B(n_240),
.C(n_236),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_702),
.B(n_662),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_707),
.B(n_585),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_710),
.A2(n_360),
.B1(n_379),
.B2(n_352),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_747),
.B(n_528),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_710),
.A2(n_765),
.B1(n_697),
.B2(n_746),
.Y(n_883)
);

NAND2x1_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_734),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_718),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_706),
.B(n_381),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_753),
.B(n_381),
.Y(n_887)
);

AND2x6_ASAP7_75t_SL g888 ( 
.A(n_772),
.B(n_258),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_766),
.B(n_528),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_821),
.B(n_662),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_747),
.B(n_320),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_830),
.B(n_671),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_830),
.B(n_671),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_708),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_725),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_834),
.B(n_671),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_719),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_831),
.B(n_320),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_698),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_719),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_697),
.B(n_320),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_691),
.B(n_589),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_746),
.A2(n_384),
.B1(n_398),
.B2(n_382),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_834),
.B(n_671),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_691),
.B(n_656),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_730),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_722),
.B(n_841),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_781),
.B(n_656),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_698),
.A2(n_382),
.B1(n_398),
.B2(n_384),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_814),
.A2(n_815),
.B1(n_840),
.B2(n_699),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_746),
.A2(n_402),
.B1(n_406),
.B2(n_399),
.Y(n_911)
);

AND2x6_ASAP7_75t_SL g912 ( 
.A(n_800),
.B(n_261),
.Y(n_912)
);

AOI22x1_ASAP7_75t_SL g913 ( 
.A1(n_739),
.A2(n_343),
.B1(n_377),
.B2(n_283),
.Y(n_913)
);

OAI22xp33_ASAP7_75t_L g914 ( 
.A1(n_840),
.A2(n_399),
.B1(n_406),
.B2(n_402),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_730),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_814),
.A2(n_387),
.B1(n_403),
.B2(n_396),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_841),
.B(n_320),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_732),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_725),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_749),
.B(n_413),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_732),
.B(n_657),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_737),
.B(n_657),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_698),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_737),
.B(n_658),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_743),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_698),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_755),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_755),
.B(n_763),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_770),
.B(n_736),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_763),
.B(n_658),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_736),
.B(n_320),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_725),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_734),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_764),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_806),
.B(n_513),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_764),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_805),
.B(n_245),
.C(n_241),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_746),
.A2(n_832),
.B1(n_799),
.B2(n_840),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_709),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_767),
.B(n_665),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_749),
.B(n_431),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_750),
.B(n_250),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_767),
.B(n_771),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_774),
.A2(n_410),
.B1(n_441),
.B2(n_366),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_757),
.B(n_758),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_771),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_779),
.B(n_409),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_787),
.B(n_665),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_787),
.B(n_667),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_734),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_689),
.B(n_461),
.Y(n_951)
);

AND2x2_ASAP7_75t_SL g952 ( 
.A(n_779),
.B(n_320),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_694),
.B(n_253),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_699),
.A2(n_427),
.B(n_428),
.C(n_409),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_792),
.B(n_667),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_792),
.B(n_812),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_812),
.B(n_668),
.Y(n_957)
);

AND2x2_ASAP7_75t_SL g958 ( 
.A(n_779),
.B(n_412),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_817),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_701),
.B(n_254),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_788),
.A2(n_681),
.B(n_675),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_840),
.B(n_589),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_799),
.A2(n_427),
.B1(n_455),
.B2(n_428),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_817),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_819),
.B(n_823),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_840),
.B(n_668),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_SL g967 ( 
.A1(n_720),
.A2(n_373),
.B1(n_278),
.B2(n_274),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_709),
.B(n_455),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_819),
.Y(n_969)
);

INVxp33_ASAP7_75t_L g970 ( 
.A(n_774),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_823),
.B(n_824),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_824),
.Y(n_972)
);

AND2x2_ASAP7_75t_SL g973 ( 
.A(n_786),
.B(n_412),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_825),
.B(n_675),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_799),
.A2(n_462),
.B1(n_412),
.B2(n_385),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_825),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_745),
.B(n_255),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_827),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_713),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_827),
.B(n_679),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_799),
.A2(n_462),
.B1(n_412),
.B2(n_385),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_806),
.B(n_412),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_681),
.B(n_679),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_832),
.A2(n_412),
.B1(n_385),
.B2(n_284),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_734),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_745),
.B(n_264),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_838),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_838),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_842),
.B(n_684),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_842),
.B(n_684),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_807),
.B(n_270),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_832),
.B(n_686),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_734),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_713),
.A2(n_513),
.B1(n_686),
.B2(n_460),
.Y(n_994)
);

NAND2x1_ASAP7_75t_L g995 ( 
.A(n_738),
.B(n_659),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_845),
.B(n_685),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_807),
.B(n_273),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_845),
.B(n_685),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_284),
.B1(n_385),
.B2(n_664),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_794),
.A2(n_683),
.B(n_664),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_703),
.B(n_664),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_733),
.B(n_685),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_733),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_690),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_690),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_696),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_786),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_699),
.B(n_571),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_696),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_699),
.B(n_685),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_693),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_839),
.B(n_282),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_703),
.B(n_285),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_704),
.B(n_685),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_703),
.B(n_288),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_705),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_703),
.B(n_290),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_704),
.B(n_685),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_705),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_704),
.B(n_693),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_704),
.A2(n_520),
.B(n_281),
.C(n_261),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_693),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_785),
.B(n_292),
.C(n_291),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_894),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_902),
.B(n_814),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_895),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_894),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_863),
.B(n_789),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_851),
.B(n_789),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_895),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_852),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_852),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_902),
.B(n_962),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_858),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_880),
.B(n_761),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_858),
.Y(n_1036)
);

BUFx12f_ASAP7_75t_L g1037 ( 
.A(n_854),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_929),
.A2(n_938),
.B1(n_883),
.B2(n_856),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_851),
.B(n_861),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_854),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_869),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_869),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_695),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_992),
.A2(n_962),
.B1(n_898),
.B2(n_881),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_854),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_920),
.B(n_750),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_875),
.B(n_864),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_895),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_935),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_860),
.B(n_768),
.Y(n_1050)
);

INVx3_ASAP7_75t_SL g1051 ( 
.A(n_859),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_874),
.B(n_695),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_941),
.B(n_716),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_870),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_870),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_874),
.B(n_695),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_900),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_885),
.B(n_727),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_860),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_900),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_915),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_885),
.B(n_727),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_915),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_918),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_918),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_992),
.A2(n_786),
.B1(n_759),
.B2(n_742),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_925),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_SL g1068 ( 
.A1(n_914),
.A2(n_280),
.B1(n_275),
.B2(n_263),
.C(n_281),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_925),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_897),
.B(n_727),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_966),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_865),
.B(n_816),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_934),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_895),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_966),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_934),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_886),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_897),
.B(n_768),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_976),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_935),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1003),
.A2(n_843),
.B1(n_847),
.B2(n_822),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_976),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_988),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_895),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_886),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_988),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1011),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1004),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1003),
.A2(n_777),
.B1(n_836),
.B2(n_820),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1007),
.B(n_850),
.Y(n_1090)
);

OR2x4_ASAP7_75t_L g1091 ( 
.A(n_977),
.B(n_263),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1007),
.B(n_744),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_906),
.B(n_711),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_939),
.B(n_979),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_876),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_919),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_919),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_935),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_886),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_906),
.B(n_741),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_936),
.B(n_946),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_936),
.B(n_946),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1004),
.Y(n_1103)
);

OR2x2_ASAP7_75t_SL g1104 ( 
.A(n_937),
.B(n_720),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1005),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_853),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1005),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_945),
.B(n_739),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_952),
.B(n_711),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_942),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1011),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_907),
.B(n_769),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_951),
.B(n_752),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_935),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_R g1116 ( 
.A(n_882),
.B(n_297),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_952),
.B(n_711),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1006),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_913),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_R g1120 ( 
.A(n_889),
.B(n_711),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_919),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_959),
.B(n_741),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_959),
.B(n_741),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1009),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_952),
.B(n_703),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_958),
.B(n_703),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_964),
.B(n_760),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_939),
.A2(n_759),
.B1(n_784),
.B2(n_744),
.Y(n_1128)
);

AO21x2_ASAP7_75t_L g1129 ( 
.A1(n_901),
.A2(n_782),
.B(n_798),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1009),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1016),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_884),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_862),
.A2(n_738),
.B1(n_773),
.B2(n_829),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_932),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1016),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_979),
.B(n_728),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_913),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_932),
.B(n_950),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1019),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_964),
.B(n_760),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_969),
.B(n_972),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_888),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1008),
.B(n_760),
.Y(n_1143)
);

BUFx4f_ASAP7_75t_L g1144 ( 
.A(n_853),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1019),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_969),
.B(n_803),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_917),
.A2(n_803),
.B(n_808),
.C(n_795),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_978),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_978),
.B(n_803),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_987),
.Y(n_1150)
);

BUFx4f_ASAP7_75t_L g1151 ( 
.A(n_853),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_903),
.A2(n_759),
.B1(n_740),
.B2(n_742),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_932),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_987),
.B(n_759),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_910),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1008),
.B(n_738),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_905),
.B(n_759),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_958),
.B(n_726),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_SL g1159 ( 
.A(n_967),
.B(n_307),
.C(n_299),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_927),
.B(n_928),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1022),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1022),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_968),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_950),
.B(n_815),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_SL g1165 ( 
.A(n_967),
.B(n_317),
.C(n_315),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_970),
.B(n_738),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_916),
.B(n_738),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_991),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_933),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_968),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1020),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_996),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_933),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_933),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_993),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_910),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_866),
.A2(n_759),
.B1(n_740),
.B2(n_742),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_958),
.B(n_773),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_968),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_853),
.Y(n_1180)
);

AOI211xp5_ASAP7_75t_L g1181 ( 
.A1(n_997),
.A2(n_338),
.B(n_321),
.C(n_322),
.Y(n_1181)
);

NOR2xp67_ASAP7_75t_L g1182 ( 
.A(n_953),
.B(n_826),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_943),
.B(n_759),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_956),
.B(n_773),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_871),
.B(n_773),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_853),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_891),
.A2(n_829),
.B(n_846),
.C(n_837),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_998),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_965),
.B(n_971),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_871),
.B(n_773),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_892),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_986),
.B(n_329),
.C(n_327),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_960),
.B(n_1012),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_923),
.B(n_809),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_877),
.A2(n_796),
.B(n_776),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_893),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_896),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_867),
.B(n_911),
.Y(n_1198)
);

AO22x1_ASAP7_75t_L g1199 ( 
.A1(n_853),
.A2(n_740),
.B1(n_742),
.B2(n_280),
.Y(n_1199)
);

AND2x2_ASAP7_75t_SL g1200 ( 
.A(n_950),
.B(n_275),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_973),
.B(n_829),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_904),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_985),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1010),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_887),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_985),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_916),
.B(n_332),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_923),
.B(n_809),
.Y(n_1208)
);

CKINVDCx8_ASAP7_75t_R g1209 ( 
.A(n_912),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_993),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1014),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_985),
.B(n_778),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_899),
.B(n_926),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_921),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_973),
.B(n_899),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_993),
.B(n_740),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_R g1217 ( 
.A(n_899),
.B(n_740),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_995),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1047),
.B(n_1023),
.C(n_878),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1072),
.B(n_908),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1096),
.A2(n_884),
.B(n_879),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1053),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1195),
.A2(n_995),
.B(n_855),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1185),
.A2(n_973),
.B(n_961),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1033),
.B(n_944),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1187),
.A2(n_947),
.B(n_1002),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1038),
.A2(n_947),
.B1(n_926),
.B2(n_963),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1190),
.A2(n_983),
.B(n_947),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_872),
.A3(n_954),
.B(n_909),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1218),
.A2(n_1018),
.B(n_1000),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1096),
.A2(n_1001),
.B(n_890),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1212),
.A2(n_1141),
.B(n_1039),
.Y(n_1232)
);

AO21x1_ASAP7_75t_L g1233 ( 
.A1(n_1193),
.A2(n_982),
.B(n_924),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1218),
.A2(n_930),
.B(n_922),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1216),
.A2(n_948),
.B(n_940),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1150),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1155),
.A2(n_1021),
.A3(n_955),
.B(n_957),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1097),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1147),
.A2(n_974),
.B(n_949),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1096),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1150),
.A2(n_989),
.B(n_980),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1160),
.A2(n_926),
.B1(n_981),
.B2(n_975),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1189),
.A2(n_868),
.B1(n_873),
.B2(n_990),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1033),
.B(n_994),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1138),
.A2(n_931),
.B(n_999),
.Y(n_1245)
);

INVx6_ASAP7_75t_L g1246 ( 
.A(n_1037),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1184),
.A2(n_887),
.B(n_1013),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1029),
.A2(n_1017),
.B(n_1015),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1138),
.A2(n_984),
.B(n_1001),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1138),
.A2(n_724),
.B(n_723),
.Y(n_1250)
);

INVx3_ASAP7_75t_SL g1251 ( 
.A(n_1111),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1096),
.A2(n_796),
.B(n_776),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1161),
.A2(n_724),
.B(n_723),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1214),
.B(n_1168),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1153),
.B(n_1203),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1166),
.B(n_887),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1025),
.B(n_887),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1184),
.A2(n_887),
.B(n_742),
.Y(n_1258)
);

OA22x2_ASAP7_75t_L g1259 ( 
.A1(n_1089),
.A2(n_295),
.B1(n_356),
.B2(n_362),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1178),
.A2(n_751),
.B(n_735),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1035),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1075),
.B(n_887),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1035),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1093),
.B(n_249),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1162),
.A2(n_762),
.B(n_756),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1166),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1097),
.A2(n_356),
.B(n_295),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1043),
.A2(n_790),
.B(n_775),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1046),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1167),
.A2(n_796),
.B1(n_848),
.B2(n_776),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_1207),
.A2(n_340),
.B(n_339),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1153),
.B(n_778),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1157),
.A2(n_790),
.B(n_775),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1075),
.B(n_809),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1042),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1093),
.B(n_249),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1153),
.A2(n_848),
.B(n_791),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1171),
.B(n_857),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_1108),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1052),
.A2(n_801),
.B(n_797),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1056),
.A2(n_801),
.B(n_797),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1148),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1027),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1148),
.Y(n_1284)
);

AO22x2_ASAP7_75t_L g1285 ( 
.A1(n_1167),
.A2(n_1117),
.B1(n_1109),
.B2(n_1158),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_L g1286 ( 
.A1(n_1028),
.A2(n_857),
.B(n_848),
.C(n_849),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1058),
.A2(n_804),
.B(n_802),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

O2A1O1Ixp5_ASAP7_75t_L g1289 ( 
.A1(n_1198),
.A2(n_1125),
.B(n_1126),
.C(n_1183),
.Y(n_1289)
);

NOR2xp67_ASAP7_75t_L g1290 ( 
.A(n_1111),
.B(n_111),
.Y(n_1290)
);

OA22x2_ASAP7_75t_L g1291 ( 
.A1(n_1081),
.A2(n_448),
.B1(n_436),
.B2(n_390),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1177),
.A2(n_804),
.B(n_802),
.Y(n_1292)
);

AOI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1031),
.A2(n_813),
.B(n_811),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1156),
.A2(n_742),
.B(n_740),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1156),
.A2(n_742),
.B(n_740),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1031),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1153),
.A2(n_1203),
.B(n_1084),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1155),
.A2(n_828),
.A3(n_846),
.B(n_837),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1042),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1026),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1153),
.A2(n_791),
.B(n_778),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1062),
.A2(n_813),
.B(n_811),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1171),
.B(n_818),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1101),
.B(n_1102),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1101),
.B(n_818),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1070),
.A2(n_835),
.B(n_828),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1026),
.Y(n_1307)
);

AO32x2_ASAP7_75t_L g1308 ( 
.A1(n_1071),
.A2(n_408),
.A3(n_407),
.B1(n_395),
.B2(n_436),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1203),
.A2(n_791),
.B(n_778),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1120),
.A2(n_249),
.B1(n_323),
.B2(n_393),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1054),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1025),
.A2(n_418),
.B(n_362),
.C(n_369),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1100),
.A2(n_849),
.B(n_835),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1097),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1054),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1122),
.A2(n_683),
.B(n_572),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1102),
.A2(n_418),
.B(n_369),
.C(n_370),
.Y(n_1317)
);

AOI211x1_ASAP7_75t_L g1318 ( 
.A1(n_1215),
.A2(n_395),
.B(n_390),
.C(n_386),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1176),
.A2(n_430),
.A3(n_433),
.B(n_429),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1203),
.A2(n_791),
.B(n_778),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1095),
.B(n_1136),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1181),
.B(n_345),
.C(n_344),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1206),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1176),
.B(n_346),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1123),
.A2(n_683),
.B(n_572),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1172),
.B(n_1188),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1172),
.B(n_791),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1154),
.A2(n_573),
.B(n_571),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1203),
.A2(n_844),
.B(n_810),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_SL g1330 ( 
.A1(n_1090),
.A2(n_783),
.B(n_809),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1114),
.A2(n_783),
.B1(n_383),
.B2(n_416),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1188),
.B(n_347),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1084),
.B(n_1200),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1204),
.B(n_1211),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_L g1335 ( 
.A(n_1113),
.B(n_354),
.C(n_348),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1204),
.B(n_355),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1211),
.B(n_358),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1200),
.A2(n_429),
.B(n_386),
.C(n_370),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1034),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1206),
.A2(n_407),
.B(n_419),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1034),
.A2(n_577),
.B(n_573),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_SL g1342 ( 
.A1(n_1206),
.A2(n_408),
.B(n_430),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1059),
.B(n_419),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1156),
.A2(n_1196),
.B(n_1191),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1106),
.A2(n_1144),
.B(n_1151),
.C(n_1044),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1090),
.A2(n_783),
.B(n_284),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_SL g1347 ( 
.A(n_1037),
.B(n_249),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_L g1348 ( 
.A(n_1090),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1191),
.B(n_359),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1196),
.B(n_367),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1127),
.A2(n_1146),
.B(n_1140),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1149),
.A2(n_581),
.B(n_577),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1169),
.A2(n_582),
.B(n_578),
.Y(n_1353)
);

AO21x1_ASAP7_75t_L g1354 ( 
.A1(n_1197),
.A2(n_448),
.B(n_433),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1036),
.A2(n_582),
.A3(n_587),
.B(n_578),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1027),
.B(n_581),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1026),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1036),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1084),
.A2(n_844),
.B(n_810),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1169),
.A2(n_587),
.B(n_586),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1197),
.A2(n_783),
.B(n_844),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1084),
.A2(n_432),
.B1(n_411),
.B2(n_375),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1095),
.B(n_323),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1106),
.A2(n_439),
.B(n_388),
.C(n_401),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1202),
.A2(n_783),
.B(n_844),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1071),
.A2(n_783),
.B1(n_391),
.B2(n_440),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1173),
.A2(n_1175),
.B(n_1174),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1173),
.A2(n_586),
.B(n_584),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1202),
.A2(n_783),
.B(n_844),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_SL g1370 ( 
.A1(n_1077),
.A2(n_584),
.B(n_174),
.Y(n_1370)
);

AND2x6_ASAP7_75t_L g1371 ( 
.A(n_1121),
.B(n_284),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1094),
.B(n_414),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1084),
.A2(n_844),
.B(n_810),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1121),
.A2(n_810),
.B(n_184),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1121),
.A2(n_810),
.B(n_181),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1094),
.B(n_415),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1136),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1128),
.A2(n_810),
.B(n_456),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1024),
.B(n_1136),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1134),
.A2(n_178),
.B(n_118),
.Y(n_1380)
);

NOR2x1_ASAP7_75t_L g1381 ( 
.A(n_1040),
.B(n_1099),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1134),
.A2(n_180),
.B(n_121),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1106),
.A2(n_452),
.B(n_450),
.C(n_443),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1240),
.B(n_1134),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1253),
.A2(n_1065),
.B(n_1060),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1236),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1345),
.A2(n_1077),
.B(n_1085),
.C(n_1055),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1266),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1228),
.A2(n_1182),
.B(n_1057),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1288),
.Y(n_1390)
);

AO32x2_ASAP7_75t_L g1391 ( 
.A1(n_1227),
.A2(n_1085),
.A3(n_1068),
.B1(n_1091),
.B2(n_1104),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1220),
.A2(n_1179),
.B1(n_1099),
.B2(n_1170),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1300),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1233),
.A2(n_1057),
.B(n_1055),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1265),
.A2(n_1065),
.B(n_1060),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1354),
.A2(n_1338),
.A3(n_1312),
.B(n_1243),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1223),
.A2(n_1069),
.B(n_1067),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1300),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1283),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1254),
.B(n_1078),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1240),
.B(n_1026),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1257),
.B(n_1143),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1269),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1377),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1240),
.B(n_1026),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1223),
.A2(n_1280),
.B(n_1268),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1324),
.B(n_1095),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1271),
.A2(n_1163),
.B1(n_1170),
.B2(n_1179),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1262),
.B(n_1213),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1324),
.B(n_1051),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1325),
.B(n_1316),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1282),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1268),
.A2(n_1069),
.B(n_1067),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1316),
.A2(n_1063),
.B(n_1061),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1284),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1304),
.B(n_1115),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1275),
.Y(n_1417)
);

CKINVDCx14_ASAP7_75t_R g1418 ( 
.A(n_1222),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1280),
.A2(n_1086),
.B(n_1082),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1275),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1257),
.B(n_1143),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1289),
.A2(n_1201),
.B(n_1143),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1288),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1300),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1299),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1299),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1311),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1281),
.A2(n_1086),
.B(n_1082),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1281),
.A2(n_1063),
.B(n_1061),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1225),
.A2(n_1115),
.B1(n_1080),
.B2(n_1049),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1261),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1255),
.B(n_1030),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1269),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1287),
.A2(n_1073),
.B(n_1064),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1287),
.A2(n_1073),
.B(n_1064),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1325),
.A2(n_1079),
.B(n_1076),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1311),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1345),
.B(n_1164),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1315),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1326),
.B(n_1076),
.Y(n_1440)
);

AOI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1219),
.A2(n_1376),
.B(n_1372),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1302),
.A2(n_1079),
.B(n_1174),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1255),
.A2(n_1151),
.B(n_1144),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1344),
.A2(n_1278),
.B(n_1242),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1238),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1302),
.A2(n_1041),
.B(n_1032),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1296),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1339),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1306),
.A2(n_1083),
.B(n_1129),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1307),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1306),
.A2(n_1199),
.B(n_1105),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1358),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1305),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1313),
.A2(n_1129),
.B(n_1217),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1238),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1338),
.A2(n_1159),
.B1(n_1165),
.B2(n_1142),
.C(n_1051),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1313),
.A2(n_1112),
.B(n_1087),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1286),
.A2(n_1201),
.B(n_1066),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1234),
.A2(n_1175),
.B(n_1210),
.Y(n_1459)
);

INVx4_ASAP7_75t_SL g1460 ( 
.A(n_1371),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1234),
.A2(n_1210),
.B(n_1088),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1235),
.A2(n_1144),
.B(n_1151),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1353),
.Y(n_1463)
);

INVx3_ASAP7_75t_SL g1464 ( 
.A(n_1251),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1334),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1263),
.B(n_1104),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1321),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1222),
.A2(n_1078),
.B1(n_1050),
.B2(n_1142),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1279),
.B(n_1349),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1379),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1352),
.A2(n_1124),
.B(n_1105),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1352),
.A2(n_1103),
.B(n_1124),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1367),
.A2(n_1118),
.B(n_1088),
.Y(n_1473)
);

AO31x2_ASAP7_75t_L g1474 ( 
.A1(n_1312),
.A2(n_1205),
.A3(n_1131),
.B(n_1130),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1367),
.A2(n_1145),
.B(n_1139),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1370),
.A2(n_1145),
.B(n_1110),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1235),
.A2(n_1247),
.B(n_1256),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_SL g1478 ( 
.A1(n_1364),
.A2(n_1098),
.B(n_1103),
.C(n_1131),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1244),
.B(n_1094),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1238),
.B(n_1030),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1356),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1347),
.A2(n_1209),
.B1(n_1119),
.B2(n_1137),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1348),
.A2(n_1205),
.B1(n_1074),
.B2(n_1186),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1348),
.A2(n_1180),
.B1(n_1186),
.B2(n_1092),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1293),
.A2(n_1250),
.B(n_1226),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1332),
.B(n_1164),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1348),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1226),
.A2(n_1239),
.B(n_1258),
.Y(n_1488)
);

O2A1O1Ixp5_ASAP7_75t_L g1489 ( 
.A1(n_1333),
.A2(n_1132),
.B(n_1199),
.C(n_1050),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1490)
);

INVx4_ASAP7_75t_SL g1491 ( 
.A(n_1371),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1250),
.A2(n_1230),
.B(n_1353),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1230),
.A2(n_1118),
.B(n_1107),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1267),
.A2(n_1342),
.B(n_1340),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1360),
.A2(n_1135),
.B(n_1107),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1360),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1303),
.Y(n_1497)
);

BUFx12f_ASAP7_75t_L g1498 ( 
.A(n_1246),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1259),
.B(n_1110),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1355),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1239),
.A2(n_1130),
.B(n_1139),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1350),
.B(n_1264),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1256),
.A2(n_1180),
.B1(n_1092),
.B2(n_1030),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1314),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1368),
.A2(n_1135),
.B(n_1152),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1355),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1276),
.A2(n_1091),
.B1(n_1050),
.B2(n_1119),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1333),
.B(n_1164),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1317),
.B(n_1091),
.Y(n_1509)
);

CKINVDCx9p33_ASAP7_75t_R g1510 ( 
.A(n_1251),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1314),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1361),
.A2(n_1129),
.B(n_1192),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1259),
.B(n_1164),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1241),
.A2(n_1030),
.B(n_1048),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1246),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1355),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1355),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1298),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1298),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1262),
.B(n_1030),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1241),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1307),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1351),
.A2(n_1346),
.B(n_1221),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1291),
.B(n_1213),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1291),
.B(n_1213),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1317),
.B(n_1116),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1246),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1262),
.B(n_1319),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1298),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1298),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_SL g1532 ( 
.A1(n_1232),
.A2(n_1048),
.B(n_1092),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1341),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1363),
.B(n_1048),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1327),
.Y(n_1535)
);

AOI221x1_ASAP7_75t_L g1536 ( 
.A1(n_1285),
.A2(n_1048),
.B1(n_1194),
.B2(n_1208),
.C(n_1092),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1237),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_SL g1538 ( 
.A(n_1290),
.B(n_1209),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1237),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1297),
.A2(n_1048),
.B(n_1194),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1260),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1322),
.A2(n_1343),
.B1(n_1335),
.B2(n_1310),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1237),
.B(n_1045),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1237),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1319),
.B(n_1045),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1362),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1319),
.B(n_1285),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1307),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1274),
.B(n_1194),
.Y(n_1549)
);

BUFx12f_ASAP7_75t_L g1550 ( 
.A(n_1307),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1365),
.A2(n_1369),
.B(n_1292),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1274),
.B(n_1208),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1260),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1274),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1318),
.B(n_1208),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1351),
.A2(n_284),
.B(n_385),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1381),
.B(n_1040),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1378),
.A2(n_426),
.B(n_424),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1273),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1249),
.A2(n_385),
.B(n_284),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1285),
.A2(n_1137),
.B1(n_393),
.B2(n_323),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1357),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1390),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1554),
.B(n_1300),
.Y(n_1564)
);

OAI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1466),
.A2(n_1546),
.B1(n_1507),
.B2(n_1490),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1558),
.A2(n_323),
.B1(n_393),
.B2(n_1380),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1412),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_L g1568 ( 
.A(n_1465),
.B(n_1314),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1502),
.B(n_1364),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1465),
.B(n_1383),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1400),
.B(n_1383),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1431),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1407),
.B(n_1319),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1410),
.A2(n_1331),
.B1(n_1357),
.B2(n_1366),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1416),
.B(n_1481),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1441),
.B(n_1382),
.C(n_1375),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1474),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1412),
.Y(n_1578)
);

INVx8_ASAP7_75t_L g1579 ( 
.A(n_1550),
.Y(n_1579)
);

AOI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1561),
.A2(n_1374),
.B1(n_1270),
.B2(n_1294),
.C(n_1295),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1456),
.B(n_1248),
.C(n_1272),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1416),
.B(n_1371),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1466),
.A2(n_1509),
.B1(n_1527),
.B2(n_1546),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_SL g1584 ( 
.A(n_1542),
.B(n_1231),
.C(n_1272),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1390),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1415),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_SL g1587 ( 
.A1(n_1555),
.A2(n_1323),
.B(n_1320),
.C(n_1309),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1479),
.B(n_1371),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1486),
.A2(n_393),
.B1(n_1292),
.B2(n_385),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1467),
.B(n_1308),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1486),
.A2(n_1323),
.B1(n_1357),
.B2(n_1301),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1498),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1468),
.A2(n_1323),
.B1(n_1277),
.B2(n_1252),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1469),
.A2(n_1371),
.B1(n_1245),
.B2(n_1249),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1399),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1507),
.B(n_1538),
.C(n_1408),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1430),
.A2(n_1273),
.B1(n_1329),
.B2(n_1359),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1467),
.B(n_1308),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1444),
.A2(n_1273),
.B(n_1373),
.Y(n_1599)
);

NAND2x1_ASAP7_75t_L g1600 ( 
.A(n_1393),
.B(n_1330),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1399),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1415),
.Y(n_1602)
);

AOI222xp33_ASAP7_75t_L g1603 ( 
.A1(n_1514),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_23),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1438),
.A2(n_385),
.B1(n_1328),
.B2(n_1308),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1447),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1386),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1470),
.A2(n_1229),
.B1(n_1328),
.B2(n_1308),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_L g1608 ( 
.A(n_1550),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1545),
.A2(n_1229),
.B1(n_385),
.B2(n_24),
.C(n_27),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_L g1610 ( 
.A(n_1482),
.B(n_1229),
.C(n_23),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1447),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1388),
.A2(n_1229),
.B1(n_24),
.B2(n_28),
.C(n_29),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1534),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1448),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1452),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1450),
.B(n_116),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1438),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_R g1618 ( 
.A(n_1403),
.B(n_231),
.Y(n_1618)
);

AND2x2_ASAP7_75t_SL g1619 ( 
.A(n_1547),
.B(n_45),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1514),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1453),
.B(n_46),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1545),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.C(n_51),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1417),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1492),
.A2(n_221),
.B(n_219),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1392),
.A2(n_48),
.B(n_50),
.C(n_51),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1403),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1402),
.B(n_53),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1453),
.B(n_53),
.Y(n_1628)
);

INVx5_ASAP7_75t_L g1629 ( 
.A(n_1424),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1402),
.B(n_54),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1420),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1528),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1497),
.B(n_54),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1498),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1440),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1510),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1549),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1425),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1421),
.B(n_60),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1421),
.B(n_1525),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1438),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1474),
.Y(n_1642)
);

AO31x2_ASAP7_75t_L g1643 ( 
.A1(n_1536),
.A2(n_62),
.A3(n_64),
.B(n_65),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1422),
.B(n_1440),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1424),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1528),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1549),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1424),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1497),
.B(n_65),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1409),
.B(n_216),
.Y(n_1650)
);

AO221x1_ASAP7_75t_L g1651 ( 
.A1(n_1494),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.C(n_74),
.Y(n_1651)
);

AND2x2_ASAP7_75t_SL g1652 ( 
.A(n_1547),
.B(n_72),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1438),
.A2(n_75),
.B1(n_81),
.B2(n_83),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1389),
.A2(n_206),
.B(n_137),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1409),
.B(n_131),
.Y(n_1655)
);

O2A1O1Ixp5_ASAP7_75t_L g1656 ( 
.A1(n_1477),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1409),
.B(n_139),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1425),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1464),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1508),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1393),
.Y(n_1661)
);

INVxp67_ASAP7_75t_SL g1662 ( 
.A(n_1404),
.Y(n_1662)
);

INVx4_ASAP7_75t_L g1663 ( 
.A(n_1393),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_L g1664 ( 
.A(n_1424),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1665)
);

OAI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1543),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.C(n_96),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1525),
.B(n_1526),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1543),
.B(n_94),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1526),
.B(n_95),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1557),
.B(n_161),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1389),
.A2(n_163),
.B(n_201),
.Y(n_1671)
);

NAND2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1424),
.B(n_98),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1433),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1393),
.Y(n_1674)
);

NAND2x1_ASAP7_75t_L g1675 ( 
.A(n_1398),
.B(n_160),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1433),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1389),
.A2(n_1462),
.B(n_1443),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1499),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1418),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1499),
.A2(n_105),
.B1(n_109),
.B2(n_127),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1529),
.A2(n_204),
.B1(n_156),
.B2(n_166),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1458),
.A2(n_141),
.B(n_167),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1529),
.B(n_170),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1535),
.A2(n_198),
.B1(n_171),
.B2(n_196),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1489),
.A2(n_1540),
.B(n_1387),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1536),
.A2(n_1508),
.B1(n_1464),
.B2(n_1557),
.Y(n_1686)
);

A2O1A1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1537),
.A2(n_1539),
.B(n_1544),
.C(n_1484),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1537),
.A2(n_1544),
.B1(n_1539),
.B2(n_1557),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1423),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1549),
.B(n_1552),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1464),
.A2(n_1557),
.B1(n_1478),
.B2(n_1503),
.C(n_1483),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1554),
.B(n_1549),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1398),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1521),
.A2(n_1504),
.B1(n_1552),
.B2(n_1516),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1521),
.A2(n_1552),
.B1(n_1398),
.B2(n_1432),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1521),
.A2(n_1552),
.B1(n_1398),
.B2(n_1432),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1562),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_R g1698 ( 
.A(n_1521),
.B(n_1445),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1513),
.A2(n_1476),
.B(n_1494),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1513),
.A2(n_1409),
.B1(n_1518),
.B2(n_1517),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1532),
.A2(n_1394),
.B(n_1406),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1548),
.B(n_1426),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1548),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1450),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1427),
.B(n_1437),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1427),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1513),
.A2(n_1518),
.B1(n_1517),
.B2(n_1506),
.Y(n_1707)
);

AOI221xp5_ASAP7_75t_L g1708 ( 
.A1(n_1476),
.A2(n_1500),
.B1(n_1506),
.B2(n_1531),
.C(n_1530),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1439),
.B(n_1396),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1500),
.A2(n_1531),
.B1(n_1530),
.B2(n_1519),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1445),
.A2(n_1511),
.B1(n_1455),
.B2(n_1523),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1533),
.A2(n_1519),
.B(n_1520),
.C(n_1560),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1520),
.A2(n_1533),
.B1(n_1522),
.B2(n_1551),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1450),
.Y(n_1715)
);

NAND2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1445),
.B(n_1511),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1450),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1391),
.A2(n_1396),
.B1(n_1522),
.B2(n_1511),
.C(n_1455),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1450),
.A2(n_1455),
.B1(n_1384),
.B2(n_1432),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1473),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1450),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1401),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1551),
.A2(n_1384),
.B(n_1532),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1394),
.A2(n_1406),
.B(n_1485),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1473),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1480),
.A2(n_1384),
.B1(n_1405),
.B2(n_1401),
.Y(n_1728)
);

CKINVDCx8_ASAP7_75t_R g1729 ( 
.A(n_1460),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1474),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1474),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1460),
.A2(n_1491),
.B1(n_1551),
.B2(n_1480),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1391),
.B(n_1474),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1480),
.B(n_1405),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1460),
.A2(n_1491),
.B1(n_1454),
.B2(n_1488),
.Y(n_1735)
);

AO21x2_ASAP7_75t_L g1736 ( 
.A1(n_1485),
.A2(n_1524),
.B(n_1556),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1401),
.A2(n_1405),
.B1(n_1463),
.B2(n_1512),
.C(n_1496),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1460),
.B(n_1491),
.Y(n_1738)
);

BUFx4f_ASAP7_75t_SL g1739 ( 
.A(n_1541),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1475),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1488),
.A2(n_1411),
.B(n_1515),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1449),
.A2(n_1457),
.B1(n_1541),
.B2(n_1553),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1515),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1391),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1491),
.B(n_1459),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1553),
.B(n_1559),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1475),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1457),
.B(n_1449),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1459),
.B(n_1461),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1559),
.A2(n_1457),
.B1(n_1512),
.B2(n_1463),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1429),
.B(n_1434),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1457),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_L g1753 ( 
.A(n_1596),
.B(n_1524),
.C(n_1556),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1622),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1619),
.A2(n_1449),
.B1(n_1436),
.B2(n_1414),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1666),
.A2(n_1496),
.B1(n_1488),
.B2(n_1436),
.C(n_1414),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1667),
.B(n_1435),
.Y(n_1757)
);

BUFx4f_ASAP7_75t_SL g1758 ( 
.A(n_1697),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1640),
.B(n_1435),
.Y(n_1759)
);

CKINVDCx6p67_ASAP7_75t_R g1760 ( 
.A(n_1592),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1741),
.A2(n_1713),
.B(n_1699),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1617),
.A2(n_1436),
.B1(n_1471),
.B2(n_1472),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1575),
.B(n_1501),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1629),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1653),
.A2(n_1411),
.B1(n_1446),
.B2(n_1454),
.C(n_1434),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1583),
.A2(n_1472),
.B1(n_1471),
.B2(n_1451),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1583),
.A2(n_1472),
.B1(n_1471),
.B2(n_1501),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_1626),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1617),
.A2(n_1472),
.B1(n_1471),
.B2(n_1501),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1641),
.A2(n_1501),
.B(n_1429),
.C(n_1461),
.Y(n_1770)
);

NAND2xp33_ASAP7_75t_R g1771 ( 
.A(n_1738),
.B(n_1397),
.Y(n_1771)
);

AO21x1_ASAP7_75t_L g1772 ( 
.A1(n_1653),
.A2(n_1442),
.B(n_1397),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1563),
.B(n_1385),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1627),
.B(n_1505),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1665),
.B(n_1569),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1641),
.A2(n_1446),
.B1(n_1428),
.B2(n_1413),
.C(n_1419),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1630),
.B(n_1505),
.Y(n_1777)
);

NAND2xp33_ASAP7_75t_R g1778 ( 
.A(n_1738),
.B(n_1493),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1577),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1565),
.A2(n_1446),
.B1(n_1442),
.B2(n_1413),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1679),
.A2(n_1493),
.B1(n_1419),
.B2(n_1395),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1565),
.A2(n_1385),
.B1(n_1395),
.B2(n_1495),
.Y(n_1782)
);

AOI222xp33_ASAP7_75t_L g1783 ( 
.A1(n_1678),
.A2(n_1495),
.B1(n_1680),
.B2(n_1612),
.C1(n_1635),
.C2(n_1660),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1668),
.B(n_1573),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1568),
.A2(n_1576),
.B(n_1682),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1563),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1673),
.A2(n_1676),
.B(n_1569),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1566),
.A2(n_1636),
.B1(n_1681),
.B2(n_1680),
.Y(n_1788)
);

OAI21xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1681),
.A2(n_1684),
.B(n_1678),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1567),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1609),
.A2(n_1613),
.B1(n_1625),
.B2(n_1566),
.C(n_1610),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1572),
.B(n_1621),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1578),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1651),
.A2(n_1574),
.B1(n_1691),
.B2(n_1618),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1659),
.A2(n_1697),
.B1(n_1689),
.B2(n_1620),
.Y(n_1796)
);

AOI222xp33_ASAP7_75t_L g1797 ( 
.A1(n_1672),
.A2(n_1684),
.B1(n_1644),
.B2(n_1628),
.C1(n_1669),
.C2(n_1649),
.Y(n_1797)
);

AOI222xp33_ASAP7_75t_L g1798 ( 
.A1(n_1672),
.A2(n_1644),
.B1(n_1633),
.B2(n_1570),
.C1(n_1639),
.C2(n_1662),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1592),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1581),
.A2(n_1584),
.B1(n_1618),
.B2(n_1580),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1601),
.B(n_1690),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1721),
.A2(n_1688),
.B1(n_1686),
.B2(n_1729),
.Y(n_1802)
);

BUFx4f_ASAP7_75t_SL g1803 ( 
.A(n_1634),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1637),
.B(n_1647),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1694),
.A2(n_1683),
.B1(n_1650),
.B2(n_1655),
.Y(n_1805)
);

AOI222xp33_ASAP7_75t_L g1806 ( 
.A1(n_1744),
.A2(n_1655),
.B1(n_1650),
.B2(n_1657),
.C1(n_1686),
.C2(n_1582),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1650),
.A2(n_1657),
.B1(n_1655),
.B2(n_1670),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1637),
.B(n_1647),
.Y(n_1808)
);

AO21x2_ASAP7_75t_L g1809 ( 
.A1(n_1599),
.A2(n_1677),
.B(n_1713),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1664),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1586),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1656),
.A2(n_1607),
.B1(n_1718),
.B2(n_1604),
.C(n_1589),
.Y(n_1812)
);

OAI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1589),
.A2(n_1688),
.B(n_1700),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1657),
.A2(n_1604),
.B1(n_1692),
.B2(n_1615),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1585),
.B(n_1692),
.Y(n_1815)
);

CKINVDCx6p67_ASAP7_75t_R g1816 ( 
.A(n_1634),
.Y(n_1816)
);

NAND2x1_ASAP7_75t_L g1817 ( 
.A(n_1722),
.B(n_1738),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1721),
.A2(n_1585),
.B1(n_1739),
.B2(n_1588),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1593),
.A2(n_1675),
.B1(n_1695),
.B2(n_1696),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1602),
.A2(n_1605),
.B1(n_1611),
.B2(n_1614),
.Y(n_1820)
);

AOI21xp33_ASAP7_75t_L g1821 ( 
.A1(n_1591),
.A2(n_1597),
.B(n_1594),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1654),
.A2(n_1671),
.B1(n_1632),
.B2(n_1616),
.C(n_1646),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1724),
.A2(n_1727),
.B1(n_1598),
.B2(n_1590),
.C1(n_1733),
.C2(n_1568),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1646),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1698),
.A2(n_1739),
.B1(n_1616),
.B2(n_1732),
.Y(n_1825)
);

INVxp33_ASAP7_75t_L g1826 ( 
.A(n_1608),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1703),
.B(n_1606),
.Y(n_1827)
);

AOI222xp33_ASAP7_75t_L g1828 ( 
.A1(n_1638),
.A2(n_1658),
.B1(n_1706),
.B2(n_1687),
.C1(n_1710),
.C2(n_1730),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1752),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1608),
.A2(n_1693),
.B1(n_1661),
.B2(n_1663),
.Y(n_1830)
);

AOI222xp33_ASAP7_75t_L g1831 ( 
.A1(n_1687),
.A2(n_1731),
.B1(n_1705),
.B2(n_1709),
.C1(n_1700),
.C2(n_1642),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_R g1832 ( 
.A(n_1745),
.B(n_1734),
.Y(n_1832)
);

OAI21xp33_ASAP7_75t_L g1833 ( 
.A1(n_1707),
.A2(n_1714),
.B(n_1642),
.Y(n_1833)
);

AOI33xp33_ASAP7_75t_L g1834 ( 
.A1(n_1707),
.A2(n_1711),
.A3(n_1714),
.B1(n_1708),
.B2(n_1742),
.B3(n_1719),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1712),
.A2(n_1693),
.B1(n_1674),
.B2(n_1661),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1674),
.B(n_1564),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1629),
.A2(n_1645),
.B1(n_1648),
.B2(n_1579),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1629),
.A2(n_1645),
.B1(n_1648),
.B2(n_1579),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1698),
.A2(n_1645),
.B1(n_1648),
.B2(n_1629),
.Y(n_1839)
);

OAI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1735),
.A2(n_1587),
.B1(n_1723),
.B2(n_1600),
.C(n_1715),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1645),
.B(n_1648),
.Y(n_1841)
);

BUFx4f_ASAP7_75t_SL g1842 ( 
.A(n_1608),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_SL g1843 ( 
.A1(n_1737),
.A2(n_1722),
.B1(n_1728),
.B2(n_1748),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1608),
.A2(n_1579),
.B1(n_1711),
.B2(n_1564),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_SL g1845 ( 
.A1(n_1624),
.A2(n_1664),
.B1(n_1745),
.B2(n_1704),
.Y(n_1845)
);

OAI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1742),
.A2(n_1623),
.B(n_1631),
.C(n_1643),
.Y(n_1846)
);

BUFx5_ASAP7_75t_L g1847 ( 
.A(n_1740),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1623),
.B(n_1664),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1643),
.B(n_1704),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1717),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1587),
.A2(n_1719),
.B(n_1716),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_1745),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1746),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1716),
.B(n_1701),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1720),
.A2(n_1726),
.B1(n_1747),
.B2(n_1701),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1726),
.A2(n_1747),
.B1(n_1750),
.B2(n_1749),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1743),
.A2(n_1751),
.B1(n_1749),
.B2(n_1643),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1743),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1643),
.A2(n_1751),
.B1(n_1725),
.B2(n_1736),
.Y(n_1859)
);

A2O1A1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1751),
.A2(n_1047),
.B(n_697),
.C(n_1193),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1736),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1725),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1626),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1729),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1869)
);

INVx8_ASAP7_75t_L g1870 ( 
.A(n_1579),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1871)
);

AO21x2_ASAP7_75t_L g1872 ( 
.A1(n_1599),
.A2(n_1699),
.B(n_1685),
.Y(n_1872)
);

BUFx12f_ASAP7_75t_L g1873 ( 
.A(n_1626),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1622),
.A2(n_748),
.B1(n_1271),
.B2(n_1047),
.C(n_1207),
.Y(n_1876)
);

OAI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1566),
.A2(n_875),
.B1(n_1047),
.B2(n_1072),
.C(n_748),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1622),
.A2(n_748),
.B1(n_1271),
.B2(n_1047),
.C(n_1207),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1567),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1575),
.B(n_1668),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1563),
.B(n_1585),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1622),
.A2(n_1666),
.B1(n_1653),
.B2(n_1609),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1601),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1885)
);

AOI222xp33_ASAP7_75t_L g1886 ( 
.A1(n_1619),
.A2(n_967),
.B1(n_1207),
.B2(n_1652),
.C1(n_623),
.C2(n_720),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1565),
.B(n_1410),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1563),
.Y(n_1888)
);

AOI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1565),
.A2(n_875),
.B(n_1047),
.C(n_748),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1892)
);

NOR2x1_ASAP7_75t_SL g1893 ( 
.A(n_1584),
.B(n_1438),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1595),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_SL g1896 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_875),
.B2(n_1047),
.Y(n_1896)
);

BUFx4f_ASAP7_75t_SL g1897 ( 
.A(n_1697),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1898)
);

AOI221xp5_ASAP7_75t_L g1899 ( 
.A1(n_1622),
.A2(n_748),
.B1(n_1271),
.B2(n_1047),
.C(n_1207),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1596),
.A2(n_875),
.B1(n_1047),
.B2(n_1072),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1697),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1567),
.Y(n_1903)
);

BUFx12f_ASAP7_75t_L g1904 ( 
.A(n_1626),
.Y(n_1904)
);

OAI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1566),
.A2(n_875),
.B1(n_1047),
.B2(n_1072),
.C(n_748),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1575),
.B(n_1465),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1702),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_SL g1909 ( 
.A(n_1584),
.B(n_1438),
.Y(n_1909)
);

OAI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1666),
.A2(n_1622),
.B1(n_1609),
.B2(n_1561),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1617),
.A2(n_1047),
.B(n_697),
.C(n_1193),
.Y(n_1912)
);

OAI222xp33_ASAP7_75t_L g1913 ( 
.A1(n_1617),
.A2(n_1641),
.B1(n_1620),
.B2(n_1622),
.C1(n_1666),
.C2(n_1678),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1567),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1622),
.A2(n_1666),
.B1(n_1653),
.B2(n_1609),
.Y(n_1916)
);

OAI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1583),
.A2(n_1047),
.B1(n_1546),
.B2(n_875),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1619),
.A2(n_1652),
.B1(n_1603),
.B2(n_1047),
.Y(n_1918)
);

AOI222xp33_ASAP7_75t_L g1919 ( 
.A1(n_1619),
.A2(n_967),
.B1(n_1207),
.B2(n_1652),
.C1(n_623),
.C2(n_720),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1857),
.B(n_1779),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1775),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1790),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1877),
.A2(n_1905),
.B1(n_1899),
.B2(n_1876),
.C(n_1878),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1829),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1794),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1811),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1858),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1879),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1903),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1779),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1847),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1757),
.B(n_1849),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1852),
.B(n_1773),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1852),
.B(n_1773),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1809),
.B(n_1759),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1809),
.B(n_1823),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1915),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1862),
.B(n_1859),
.Y(n_1938)
);

INVx4_ASAP7_75t_L g1939 ( 
.A(n_1841),
.Y(n_1939)
);

AND2x4_ASAP7_75t_SL g1940 ( 
.A(n_1819),
.B(n_1764),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1763),
.B(n_1853),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1859),
.B(n_1784),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1896),
.A2(n_1908),
.B1(n_1898),
.B2(n_1883),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1872),
.B(n_1861),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1856),
.B(n_1872),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1856),
.B(n_1855),
.Y(n_1946)
);

NOR2x1_ASAP7_75t_L g1947 ( 
.A(n_1839),
.B(n_1822),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1855),
.B(n_1755),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1755),
.B(n_1761),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1851),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1761),
.B(n_1854),
.Y(n_1951)
);

INVxp67_ASAP7_75t_SL g1952 ( 
.A(n_1772),
.Y(n_1952)
);

CKINVDCx14_ASAP7_75t_R g1953 ( 
.A(n_1768),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1761),
.B(n_1767),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1828),
.B(n_1831),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1854),
.B(n_1774),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1777),
.B(n_1833),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1780),
.B(n_1765),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1834),
.B(n_1860),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1865),
.A2(n_1874),
.B1(n_1917),
.B2(n_1871),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1834),
.B(n_1860),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1839),
.B(n_1825),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1906),
.B(n_1820),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1766),
.B(n_1769),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1762),
.B(n_1782),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1762),
.B(n_1782),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1832),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1786),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1832),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1786),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1756),
.B(n_1866),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1820),
.B(n_1792),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1869),
.B(n_1875),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1885),
.B(n_1894),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1776),
.B(n_1893),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1846),
.Y(n_1976)
);

AND2x4_ASAP7_75t_SL g1977 ( 
.A(n_1764),
.B(n_1807),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1907),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1909),
.B(n_1753),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1825),
.B(n_1840),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1848),
.B(n_1821),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1813),
.B(n_1806),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1881),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1827),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1801),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1778),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1887),
.B(n_1800),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1887),
.B(n_1800),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1880),
.B(n_1770),
.Y(n_1989)
);

NOR2x1_ASAP7_75t_SL g1990 ( 
.A(n_1802),
.B(n_1844),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1812),
.B(n_1781),
.Y(n_1991)
);

OA21x2_ASAP7_75t_L g1992 ( 
.A1(n_1785),
.A2(n_1781),
.B(n_1912),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1778),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1886),
.A2(n_1919),
.B1(n_1918),
.B2(n_1914),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1845),
.B(n_1814),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1804),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_SL g1997 ( 
.A(n_1888),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1808),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1817),
.Y(n_1999)
);

NAND2x1_ASAP7_75t_L g2000 ( 
.A(n_1807),
.B(n_1835),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_SL g2001 ( 
.A(n_1818),
.B(n_1810),
.Y(n_2001)
);

OAI321xp33_ASAP7_75t_L g2002 ( 
.A1(n_1889),
.A2(n_1918),
.A3(n_1914),
.B1(n_1911),
.B2(n_1863),
.C(n_1900),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1843),
.Y(n_2003)
);

INVxp67_ASAP7_75t_L g2004 ( 
.A(n_1771),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1771),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1850),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1863),
.A2(n_1867),
.B1(n_1911),
.B2(n_1890),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1912),
.B(n_1884),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1798),
.B(n_1901),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1932),
.B(n_1902),
.Y(n_2010)
);

INVxp33_ASAP7_75t_SL g2011 ( 
.A(n_1967),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_1968),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1956),
.B(n_1895),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1924),
.Y(n_2014)
);

INVxp67_ASAP7_75t_SL g2015 ( 
.A(n_1967),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1923),
.A2(n_1867),
.B1(n_1890),
.B2(n_1900),
.C(n_1891),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1923),
.A2(n_1789),
.B(n_1892),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1932),
.B(n_1815),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_R g2019 ( 
.A(n_1953),
.B(n_1864),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1932),
.B(n_1805),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1922),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1921),
.B(n_1793),
.Y(n_2022)
);

O2A1O1Ixp33_ASAP7_75t_L g2023 ( 
.A1(n_2002),
.A2(n_1910),
.B(n_1913),
.C(n_1916),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1956),
.B(n_1795),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1922),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_1921),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1960),
.B(n_1892),
.C(n_1891),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1994),
.A2(n_1754),
.B1(n_1788),
.B2(n_1916),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_1994),
.A2(n_1754),
.B1(n_1791),
.B2(n_1796),
.C(n_1797),
.Y(n_2029)
);

OAI322xp33_ASAP7_75t_L g2030 ( 
.A1(n_1955),
.A2(n_1882),
.A3(n_1787),
.B1(n_1824),
.B2(n_1830),
.C1(n_1868),
.C2(n_1799),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1933),
.B(n_1836),
.Y(n_2031)
);

INVx3_ASAP7_75t_SL g2032 ( 
.A(n_1970),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1968),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1985),
.B(n_1882),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2002),
.A2(n_1826),
.B1(n_1868),
.B2(n_1870),
.C(n_1836),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1985),
.B(n_1783),
.Y(n_2036)
);

AOI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_2009),
.A2(n_1870),
.B1(n_1838),
.B2(n_1837),
.C(n_1758),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1956),
.B(n_1760),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1987),
.B(n_1758),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1942),
.B(n_1816),
.Y(n_2040)
);

INVx3_ASAP7_75t_SL g2041 ( 
.A(n_1970),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1925),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2007),
.A2(n_1943),
.B1(n_1987),
.B2(n_1988),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_L g2044 ( 
.A(n_2009),
.B(n_1897),
.C(n_1803),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1942),
.B(n_1870),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1925),
.Y(n_2046)
);

AOI221x1_ASAP7_75t_SL g2047 ( 
.A1(n_1955),
.A2(n_1897),
.B1(n_1803),
.B2(n_1842),
.C(n_1873),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1935),
.B(n_1904),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1933),
.B(n_1842),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1926),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1930),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1935),
.B(n_1936),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1978),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_1988),
.B(n_2003),
.C(n_1958),
.Y(n_2054)
);

AOI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_1936),
.A2(n_1982),
.B1(n_1958),
.B2(n_1959),
.C(n_1961),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1930),
.Y(n_2056)
);

OAI33xp33_ASAP7_75t_L g2057 ( 
.A1(n_2003),
.A2(n_1972),
.A3(n_1989),
.B1(n_1963),
.B2(n_1937),
.B3(n_1941),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1982),
.A2(n_1991),
.B1(n_1959),
.B2(n_1961),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1982),
.A2(n_1980),
.B1(n_1991),
.B2(n_1959),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1927),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1927),
.Y(n_2061)
);

NAND4xp25_ASAP7_75t_L g2062 ( 
.A(n_1972),
.B(n_1936),
.C(n_1989),
.D(n_1991),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1969),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1928),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1978),
.Y(n_2065)
);

NAND4xp25_ASAP7_75t_L g2066 ( 
.A(n_1989),
.B(n_1958),
.C(n_1961),
.D(n_1980),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_L g2067 ( 
.A(n_1963),
.B(n_1950),
.C(n_2008),
.D(n_1947),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1928),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1929),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1999),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1929),
.Y(n_2071)
);

NAND4xp25_ASAP7_75t_L g2072 ( 
.A(n_1950),
.B(n_2008),
.C(n_1947),
.D(n_1971),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1933),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1962),
.A2(n_2000),
.B1(n_1969),
.B2(n_2006),
.Y(n_2074)
);

OAI211xp5_ASAP7_75t_L g2075 ( 
.A1(n_1976),
.A2(n_1952),
.B(n_2000),
.C(n_1992),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1935),
.B(n_1986),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1962),
.A2(n_2006),
.B1(n_1976),
.B2(n_1940),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1983),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1986),
.B(n_1993),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1970),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1940),
.A2(n_1995),
.B1(n_1977),
.B2(n_2004),
.Y(n_2081)
);

OAI31xp33_ASAP7_75t_L g2082 ( 
.A1(n_1995),
.A2(n_1940),
.A3(n_1965),
.B(n_1966),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2008),
.A2(n_1995),
.B1(n_1971),
.B2(n_1966),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1993),
.B(n_2005),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1978),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1942),
.B(n_2005),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1971),
.A2(n_1966),
.B1(n_1965),
.B2(n_1975),
.Y(n_2087)
);

AOI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1992),
.A2(n_1952),
.B(n_1990),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_SL g2089 ( 
.A1(n_1990),
.A2(n_1965),
.B1(n_2001),
.B2(n_1992),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2004),
.B(n_1957),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2052),
.B(n_1937),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2032),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2063),
.Y(n_2093)
);

NAND2x1_ASAP7_75t_L g2094 ( 
.A(n_2070),
.B(n_1931),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2052),
.B(n_2087),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2014),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2076),
.B(n_1951),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2051),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2039),
.B(n_1973),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2032),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2090),
.B(n_1951),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2026),
.B(n_1941),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2090),
.B(n_1951),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2079),
.B(n_1949),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2079),
.B(n_1938),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2084),
.B(n_1984),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_2056),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2086),
.B(n_1954),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2084),
.B(n_1938),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2015),
.B(n_1984),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2073),
.B(n_2049),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2073),
.B(n_1949),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_2074),
.B(n_1999),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2028),
.A2(n_1992),
.B1(n_1975),
.B2(n_1964),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2086),
.B(n_1949),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_2041),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2053),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2053),
.Y(n_2118)
);

INVx1_ASAP7_75t_SL g2119 ( 
.A(n_2041),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2083),
.B(n_1996),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2065),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2010),
.B(n_1975),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2010),
.B(n_1979),
.Y(n_2123)
);

OR2x2_ASAP7_75t_L g2124 ( 
.A(n_2085),
.B(n_1954),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2013),
.B(n_2062),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2021),
.B(n_1954),
.Y(n_2126)
);

OR2x6_ASAP7_75t_L g2127 ( 
.A(n_2088),
.B(n_1979),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2025),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_2042),
.B(n_1920),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2018),
.B(n_1979),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_2039),
.B(n_1974),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_2046),
.B(n_1920),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2018),
.B(n_2060),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2050),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2020),
.B(n_1945),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2020),
.B(n_1945),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2060),
.B(n_1964),
.Y(n_2137)
);

INVx4_ASAP7_75t_L g2138 ( 
.A(n_2070),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2061),
.B(n_1964),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2061),
.B(n_1934),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2064),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2048),
.B(n_1934),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2068),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2069),
.B(n_1998),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_2092),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2128),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2120),
.B(n_2054),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2128),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2120),
.B(n_2022),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2128),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2108),
.B(n_2126),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2102),
.B(n_2055),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2104),
.B(n_2048),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2104),
.B(n_2038),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2104),
.B(n_2038),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2141),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2102),
.B(n_2072),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2141),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2141),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_L g2160 ( 
.A(n_2113),
.B(n_2029),
.C(n_2023),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2099),
.B(n_2059),
.Y(n_2161)
);

NAND2x1p5_ASAP7_75t_L g2162 ( 
.A(n_2094),
.B(n_1992),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2111),
.B(n_2070),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2135),
.B(n_2070),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2129),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_2100),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2129),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2132),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2135),
.B(n_2078),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2135),
.B(n_2011),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2136),
.B(n_2089),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2134),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2136),
.B(n_2031),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_2111),
.B(n_2031),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2136),
.B(n_2031),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2134),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2143),
.Y(n_2177)
);

NOR2x1_ASAP7_75t_SL g2178 ( 
.A(n_2127),
.B(n_2075),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2132),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2096),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2101),
.B(n_2012),
.Y(n_2181)
);

AOI32xp33_ASAP7_75t_L g2182 ( 
.A1(n_2095),
.A2(n_2058),
.A3(n_2043),
.B1(n_2016),
.B2(n_2024),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2143),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2117),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2108),
.B(n_1920),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2101),
.B(n_2012),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2125),
.B(n_2122),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2117),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2118),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_2138),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2101),
.B(n_2033),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2096),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2125),
.B(n_2011),
.Y(n_2193)
);

NOR2x1p5_ASAP7_75t_SL g2194 ( 
.A(n_2126),
.B(n_1944),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2111),
.B(n_2080),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2122),
.B(n_2067),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2118),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2121),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2103),
.B(n_2033),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2091),
.B(n_2071),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2121),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2152),
.B(n_2095),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2157),
.B(n_2123),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2185),
.B(n_2091),
.Y(n_2204)
);

NOR2x1_ASAP7_75t_L g2205 ( 
.A(n_2145),
.B(n_2066),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2183),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2183),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2180),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2147),
.A2(n_2017),
.B(n_2057),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2149),
.B(n_2166),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2180),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2192),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2178),
.B(n_2171),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2178),
.B(n_2115),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2160),
.A2(n_2027),
.B1(n_2114),
.B2(n_2036),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2185),
.B(n_2093),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2171),
.B(n_2115),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2161),
.B(n_2123),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2174),
.B(n_2115),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2165),
.B(n_2093),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2192),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2182),
.B(n_2024),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2193),
.B(n_2058),
.C(n_2114),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_2145),
.Y(n_2224)
);

BUFx3_ASAP7_75t_L g2225 ( 
.A(n_2190),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2196),
.B(n_2105),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2172),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2174),
.B(n_2195),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2154),
.B(n_2105),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_2170),
.B(n_2131),
.Y(n_2230)
);

NAND4xp25_ASAP7_75t_L g2231 ( 
.A(n_2187),
.B(n_2047),
.C(n_2034),
.D(n_2044),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2174),
.B(n_2130),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2174),
.B(n_2130),
.Y(n_2233)
);

AND2x4_ASAP7_75t_L g2234 ( 
.A(n_2190),
.B(n_2127),
.Y(n_2234)
);

NAND2xp33_ASAP7_75t_R g2235 ( 
.A(n_2190),
.B(n_2019),
.Y(n_2235)
);

NOR2x1_ASAP7_75t_L g2236 ( 
.A(n_2163),
.B(n_2138),
.Y(n_2236)
);

INVxp67_ASAP7_75t_L g2237 ( 
.A(n_2164),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2176),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2177),
.Y(n_2239)
);

NOR3xp33_ASAP7_75t_SL g2240 ( 
.A(n_2165),
.B(n_2030),
.C(n_2077),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2184),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_2195),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2167),
.B(n_2124),
.Y(n_2243)
);

NAND4xp25_ASAP7_75t_L g2244 ( 
.A(n_2167),
.B(n_2037),
.C(n_2082),
.D(n_2035),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2146),
.Y(n_2245)
);

NOR2xp67_ASAP7_75t_SL g2246 ( 
.A(n_2164),
.B(n_2040),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2184),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2195),
.B(n_2111),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2188),
.Y(n_2249)
);

INVx3_ASAP7_75t_L g2250 ( 
.A(n_2195),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2163),
.B(n_2092),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2168),
.B(n_2179),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2163),
.B(n_2103),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2153),
.B(n_2100),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2188),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2189),
.Y(n_2256)
);

AOI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_2209),
.A2(n_2127),
.B(n_2110),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2215),
.B(n_2153),
.Y(n_2258)
);

AOI21xp33_ASAP7_75t_SL g2259 ( 
.A1(n_2222),
.A2(n_2127),
.B(n_2162),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2253),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_2224),
.Y(n_2261)
);

INVx1_ASAP7_75t_SL g2262 ( 
.A(n_2205),
.Y(n_2262)
);

XNOR2x1_ASAP7_75t_L g2263 ( 
.A(n_2205),
.B(n_2154),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_L g2264 ( 
.A1(n_2223),
.A2(n_1948),
.B1(n_1945),
.B2(n_1946),
.Y(n_2264)
);

AO21x1_ASAP7_75t_L g2265 ( 
.A1(n_2235),
.A2(n_2163),
.B(n_2138),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2228),
.B(n_2173),
.Y(n_2266)
);

INVxp33_ASAP7_75t_L g2267 ( 
.A(n_2246),
.Y(n_2267)
);

NOR3xp33_ASAP7_75t_L g2268 ( 
.A(n_2223),
.B(n_2138),
.C(n_2081),
.Y(n_2268)
);

OAI21xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2213),
.A2(n_2175),
.B(n_2173),
.Y(n_2269)
);

AOI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2213),
.A2(n_2127),
.B1(n_2168),
.B2(n_2179),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2244),
.A2(n_1948),
.B1(n_1946),
.B2(n_2127),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2254),
.A2(n_2246),
.B1(n_2237),
.B2(n_2202),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2253),
.Y(n_2273)
);

AOI311xp33_ASAP7_75t_L g2274 ( 
.A1(n_2206),
.A2(n_2158),
.A3(n_2148),
.B(n_2150),
.C(n_2156),
.Y(n_2274)
);

OAI221xp5_ASAP7_75t_SL g2275 ( 
.A1(n_2244),
.A2(n_2119),
.B1(n_2116),
.B2(n_2151),
.C(n_2045),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2240),
.B(n_2155),
.Y(n_2276)
);

NAND2xp33_ASAP7_75t_L g2277 ( 
.A(n_2236),
.B(n_2019),
.Y(n_2277)
);

OAI21xp5_ASAP7_75t_L g2278 ( 
.A1(n_2236),
.A2(n_2162),
.B(n_2119),
.Y(n_2278)
);

OA22x2_ASAP7_75t_L g2279 ( 
.A1(n_2224),
.A2(n_2116),
.B1(n_2169),
.B2(n_2107),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2206),
.Y(n_2280)
);

OAI21xp33_ASAP7_75t_L g2281 ( 
.A1(n_2231),
.A2(n_2194),
.B(n_2200),
.Y(n_2281)
);

AND2x4_ASAP7_75t_SL g2282 ( 
.A(n_2224),
.B(n_2251),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2210),
.B(n_2155),
.Y(n_2283)
);

AOI21xp33_ASAP7_75t_L g2284 ( 
.A1(n_2251),
.A2(n_2045),
.B(n_2200),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2225),
.B(n_2175),
.Y(n_2285)
);

OAI21xp33_ASAP7_75t_SL g2286 ( 
.A1(n_2214),
.A2(n_2169),
.B(n_2151),
.Y(n_2286)
);

NAND2x1p5_ASAP7_75t_L g2287 ( 
.A(n_2225),
.B(n_2094),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2219),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2207),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2203),
.A2(n_2162),
.B(n_2110),
.Y(n_2290)
);

AO22x1_ASAP7_75t_L g2291 ( 
.A1(n_2214),
.A2(n_2107),
.B1(n_2098),
.B2(n_2137),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2226),
.B(n_2106),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2207),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2227),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2228),
.B(n_2181),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2242),
.A2(n_2158),
.B(n_2146),
.Y(n_2296)
);

NAND2xp33_ASAP7_75t_SL g2297 ( 
.A(n_2242),
.B(n_2098),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2219),
.Y(n_2298)
);

OAI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2262),
.A2(n_2218),
.B1(n_2250),
.B2(n_2216),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2275),
.B(n_2252),
.C(n_2238),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2267),
.B(n_2230),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2280),
.Y(n_2302)
);

OAI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_2271),
.A2(n_2217),
.B(n_2252),
.Y(n_2303)
);

NAND4xp25_ASAP7_75t_L g2304 ( 
.A(n_2271),
.B(n_2217),
.C(n_2250),
.D(n_2234),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2276),
.B(n_2229),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2282),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2277),
.A2(n_2250),
.B1(n_2248),
.B2(n_2234),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2261),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2289),
.Y(n_2309)
);

O2A1O1Ixp33_ASAP7_75t_L g2310 ( 
.A1(n_2277),
.A2(n_2281),
.B(n_2257),
.C(n_2268),
.Y(n_2310)
);

OAI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2267),
.A2(n_2216),
.B1(n_2204),
.B2(n_2220),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2261),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_2282),
.B(n_2248),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_SL g2314 ( 
.A1(n_2263),
.A2(n_2001),
.B1(n_2234),
.B2(n_1948),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2265),
.B(n_2234),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2258),
.B(n_2232),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2293),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2294),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2264),
.B(n_2232),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_2261),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2260),
.Y(n_2321)
);

NOR3xp33_ASAP7_75t_L g2322 ( 
.A(n_2297),
.B(n_2238),
.C(n_2239),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2272),
.B(n_2204),
.Y(n_2323)
);

NAND3xp33_ASAP7_75t_L g2324 ( 
.A(n_2264),
.B(n_2239),
.C(n_2227),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2263),
.A2(n_2233),
.B1(n_2220),
.B2(n_2243),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2279),
.A2(n_2211),
.B(n_2212),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2260),
.B(n_2233),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2297),
.A2(n_2256),
.B1(n_2255),
.B2(n_2249),
.C(n_2247),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2273),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2320),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2320),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2314),
.B(n_2279),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2312),
.Y(n_2333)
);

OAI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2310),
.A2(n_2300),
.B(n_2322),
.Y(n_2334)
);

INVxp67_ASAP7_75t_SL g2335 ( 
.A(n_2322),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2321),
.Y(n_2336)
);

NOR3xp33_ASAP7_75t_SL g2337 ( 
.A(n_2304),
.B(n_2278),
.C(n_2286),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2313),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2301),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2306),
.B(n_2273),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2329),
.Y(n_2341)
);

INVx2_ASAP7_75t_SL g2342 ( 
.A(n_2313),
.Y(n_2342)
);

AOI322xp5_ASAP7_75t_L g2343 ( 
.A1(n_2323),
.A2(n_2269),
.A3(n_2284),
.B1(n_2298),
.B2(n_2288),
.C1(n_2270),
.C2(n_2283),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2316),
.B(n_2288),
.Y(n_2344)
);

XOR2xp5_ASAP7_75t_L g2345 ( 
.A(n_2307),
.B(n_2285),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_R g2346 ( 
.A(n_2326),
.B(n_2259),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2314),
.B(n_2266),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2315),
.A2(n_2287),
.B(n_2296),
.Y(n_2348)
);

INVx1_ASAP7_75t_SL g2349 ( 
.A(n_2325),
.Y(n_2349)
);

NOR3xp33_ASAP7_75t_SL g2350 ( 
.A(n_2299),
.B(n_2290),
.C(n_2247),
.Y(n_2350)
);

CKINVDCx20_ASAP7_75t_R g2351 ( 
.A(n_2305),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2303),
.B(n_2285),
.Y(n_2352)
);

INVx2_ASAP7_75t_SL g2353 ( 
.A(n_2342),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2342),
.B(n_2311),
.Y(n_2354)
);

NOR3xp33_ASAP7_75t_L g2355 ( 
.A(n_2334),
.B(n_2319),
.C(n_2308),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2339),
.B(n_2324),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2351),
.B(n_2327),
.Y(n_2357)
);

OAI21xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2332),
.A2(n_2328),
.B(n_2308),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2338),
.B(n_2318),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2338),
.B(n_2302),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2335),
.B(n_2349),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_L g2362 ( 
.A(n_2340),
.B(n_2317),
.C(n_2309),
.Y(n_2362)
);

AOI21xp33_ASAP7_75t_SL g2363 ( 
.A1(n_2345),
.A2(n_2348),
.B(n_2352),
.Y(n_2363)
);

OAI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2350),
.A2(n_2298),
.B1(n_2285),
.B2(n_2287),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2351),
.B(n_2295),
.Y(n_2365)
);

NOR3xp33_ASAP7_75t_L g2366 ( 
.A(n_2344),
.B(n_2291),
.C(n_2292),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2348),
.A2(n_2241),
.B(n_2256),
.Y(n_2367)
);

AO21x1_ASAP7_75t_L g2368 ( 
.A1(n_2363),
.A2(n_2331),
.B(n_2330),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2353),
.B(n_2333),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2355),
.A2(n_2347),
.B1(n_2345),
.B2(n_2337),
.Y(n_2370)
);

NAND4xp25_ASAP7_75t_L g2371 ( 
.A(n_2357),
.B(n_2361),
.C(n_2356),
.D(n_2354),
.Y(n_2371)
);

NAND4xp25_ASAP7_75t_SL g2372 ( 
.A(n_2358),
.B(n_2343),
.C(n_2366),
.D(n_2365),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2362),
.B(n_2333),
.Y(n_2373)
);

AOI21xp33_ASAP7_75t_L g2374 ( 
.A1(n_2364),
.A2(n_2346),
.B(n_2331),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2359),
.B(n_2360),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2367),
.A2(n_2347),
.B1(n_2330),
.B2(n_2336),
.Y(n_2376)
);

O2A1O1Ixp33_ASAP7_75t_L g2377 ( 
.A1(n_2363),
.A2(n_2341),
.B(n_2336),
.C(n_2274),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2353),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_2365),
.B(n_2341),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2358),
.A2(n_2255),
.B(n_2249),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_L g2381 ( 
.A(n_2365),
.B(n_2243),
.Y(n_2381)
);

XNOR2xp5_ASAP7_75t_L g2382 ( 
.A(n_2365),
.B(n_1977),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_R g2383 ( 
.A(n_2378),
.B(n_1997),
.Y(n_2383)
);

OAI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_2370),
.A2(n_2241),
.B(n_2212),
.Y(n_2384)
);

AOI221xp5_ASAP7_75t_L g2385 ( 
.A1(n_2372),
.A2(n_2221),
.B1(n_2211),
.B2(n_2208),
.C(n_2245),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2369),
.Y(n_2386)
);

XNOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2376),
.B(n_2194),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2368),
.A2(n_2221),
.B(n_2208),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2373),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2374),
.A2(n_2245),
.B(n_2148),
.Y(n_2390)
);

AOI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2377),
.A2(n_2201),
.B1(n_2189),
.B2(n_2198),
.C(n_2197),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_R g2392 ( 
.A(n_2375),
.B(n_2137),
.Y(n_2392)
);

NOR3xp33_ASAP7_75t_L g2393 ( 
.A(n_2389),
.B(n_2371),
.C(n_2379),
.Y(n_2393)
);

NOR2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2386),
.B(n_2381),
.Y(n_2394)
);

NOR4xp75_ASAP7_75t_L g2395 ( 
.A(n_2384),
.B(n_2380),
.C(n_2382),
.D(n_2106),
.Y(n_2395)
);

NAND4xp25_ASAP7_75t_L g2396 ( 
.A(n_2391),
.B(n_2139),
.C(n_1999),
.D(n_2109),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2387),
.Y(n_2397)
);

NOR2x1_ASAP7_75t_L g2398 ( 
.A(n_2388),
.B(n_2150),
.Y(n_2398)
);

NAND4xp75_ASAP7_75t_L g2399 ( 
.A(n_2390),
.B(n_2139),
.C(n_2199),
.D(n_2186),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2383),
.Y(n_2400)
);

NAND3xp33_ASAP7_75t_SL g2401 ( 
.A(n_2393),
.B(n_2385),
.C(n_2392),
.Y(n_2401)
);

XOR2xp5_ASAP7_75t_L g2402 ( 
.A(n_2400),
.B(n_2142),
.Y(n_2402)
);

AOI211xp5_ASAP7_75t_L g2403 ( 
.A1(n_2397),
.A2(n_2109),
.B(n_2199),
.C(n_2181),
.Y(n_2403)
);

NOR3xp33_ASAP7_75t_L g2404 ( 
.A(n_2396),
.B(n_1939),
.C(n_2142),
.Y(n_2404)
);

OAI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2399),
.A2(n_2156),
.B1(n_2159),
.B2(n_2197),
.Y(n_2405)
);

AOI22xp33_ASAP7_75t_L g2406 ( 
.A1(n_2394),
.A2(n_1997),
.B1(n_1939),
.B2(n_1946),
.Y(n_2406)
);

NAND3xp33_ASAP7_75t_SL g2407 ( 
.A(n_2395),
.B(n_2186),
.C(n_2191),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2402),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2401),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2407),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2405),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2406),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2409),
.A2(n_2398),
.B(n_2404),
.Y(n_2413)
);

CKINVDCx20_ASAP7_75t_R g2414 ( 
.A(n_2408),
.Y(n_2414)
);

AND2x2_ASAP7_75t_SL g2415 ( 
.A(n_2414),
.B(n_2410),
.Y(n_2415)
);

INVxp67_ASAP7_75t_L g2416 ( 
.A(n_2415),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2415),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2416),
.A2(n_2412),
.B1(n_2411),
.B2(n_2413),
.Y(n_2418)
);

AOI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2417),
.A2(n_2411),
.B1(n_2412),
.B2(n_2403),
.C(n_2159),
.Y(n_2419)
);

NAND5xp2_ASAP7_75t_L g2420 ( 
.A(n_2419),
.B(n_1981),
.C(n_1957),
.D(n_2103),
.E(n_2191),
.Y(n_2420)
);

OR2x6_ASAP7_75t_L g2421 ( 
.A(n_2418),
.B(n_2133),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_L g2422 ( 
.A(n_2421),
.B(n_2201),
.C(n_2198),
.Y(n_2422)
);

AOI221xp5_ASAP7_75t_L g2423 ( 
.A1(n_2422),
.A2(n_2420),
.B1(n_1997),
.B2(n_2097),
.C(n_2133),
.Y(n_2423)
);

AOI211xp5_ASAP7_75t_L g2424 ( 
.A1(n_2423),
.A2(n_2112),
.B(n_2140),
.C(n_2144),
.Y(n_2424)
);


endmodule